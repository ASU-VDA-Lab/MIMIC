module fake_jpeg_29693_n_516 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_516);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_516;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_51),
.B(n_65),
.Y(n_129)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_75),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_81),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_14),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_14),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_34),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_91),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_41),
.B(n_22),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_99),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_13),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_93),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_13),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_81),
.CON(n_102),
.SN(n_102)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_102),
.B(n_105),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_47),
.B(n_42),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_32),
.C(n_49),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_125),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_47),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_117),
.B(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_47),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_50),
.B(n_32),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_126),
.B(n_132),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_56),
.A2(n_32),
.B1(n_29),
.B2(n_39),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_150),
.B1(n_27),
.B2(n_25),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_144),
.B(n_152),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_53),
.A2(n_32),
.B1(n_29),
.B2(n_40),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_40),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_63),
.A2(n_18),
.B1(n_45),
.B2(n_43),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_22),
.B1(n_25),
.B2(n_35),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_39),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_159),
.Y(n_208)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_158),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_39),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_105),
.A2(n_52),
.B1(n_88),
.B2(n_16),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_168),
.B1(n_177),
.B2(n_180),
.Y(n_207)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_27),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_173),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_29),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_169),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_112),
.A2(n_55),
.B1(n_57),
.B2(n_78),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_22),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_187),
.B1(n_197),
.B2(n_45),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_27),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_112),
.A2(n_67),
.B1(n_72),
.B2(n_77),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_76),
.B1(n_73),
.B2(n_74),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_185),
.B1(n_127),
.B2(n_16),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_111),
.A2(n_35),
.B1(n_18),
.B2(n_49),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_25),
.B1(n_43),
.B2(n_35),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_191),
.Y(n_239)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_194),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_21),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_200),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_21),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_101),
.A2(n_59),
.B1(n_87),
.B2(n_79),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_119),
.A2(n_62),
.B1(n_98),
.B2(n_99),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_102),
.B(n_88),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_123),
.B(n_124),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_135),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_101),
.B(n_46),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_46),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_134),
.A2(n_43),
.B1(n_18),
.B2(n_49),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_135),
.C(n_150),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_16),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_107),
.B1(n_100),
.B2(n_120),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_211),
.A2(n_212),
.B1(n_184),
.B2(n_164),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_107),
.B1(n_100),
.B2(n_120),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_221),
.B1(n_175),
.B2(n_207),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_207),
.B1(n_243),
.B2(n_197),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_133),
.B(n_115),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_175),
.B(n_162),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_103),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_244),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_226),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_227),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_148),
.B1(n_121),
.B2(n_103),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_235),
.B1(n_238),
.B2(n_198),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_183),
.A2(n_121),
.B1(n_108),
.B2(n_148),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_116),
.C(n_108),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_188),
.C(n_162),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_162),
.A2(n_180),
.B1(n_173),
.B2(n_170),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_159),
.B(n_193),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_245),
.A2(n_271),
.B1(n_274),
.B2(n_277),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_166),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_269),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_247),
.B(n_135),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_263),
.B1(n_266),
.B2(n_268),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_237),
.B(n_206),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_256),
.B(n_237),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_175),
.C(n_200),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_258),
.C(n_220),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_219),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_194),
.B(n_164),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_178),
.C(n_195),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_192),
.B1(n_179),
.B2(n_171),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_209),
.B(n_181),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_241),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_210),
.A2(n_161),
.B1(n_189),
.B2(n_119),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_267),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_212),
.B1(n_225),
.B2(n_208),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_224),
.B(n_204),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_209),
.A2(n_244),
.B1(n_211),
.B2(n_223),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_278),
.B1(n_279),
.B2(n_242),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_273),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_214),
.A2(n_186),
.B1(n_155),
.B2(n_158),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_191),
.B1(n_165),
.B2(n_190),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_227),
.A2(n_96),
.B1(n_163),
.B2(n_176),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_293),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_239),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_289),
.B(n_296),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_241),
.B1(n_232),
.B2(n_228),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_312),
.B1(n_263),
.B2(n_279),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_311),
.B(n_298),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_295),
.A2(n_301),
.B(n_247),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_216),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_270),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_300),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_231),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_249),
.A2(n_250),
.B(n_256),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_240),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_308),
.C(n_258),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_215),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_306),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_215),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_272),
.B1(n_266),
.B2(n_248),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_250),
.B1(n_271),
.B2(n_274),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_19),
.B(n_45),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_245),
.A2(n_232),
.B1(n_228),
.B2(n_240),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_220),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_313),
.B(n_260),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_220),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_282),
.B(n_246),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_317),
.B(n_343),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_318),
.A2(n_340),
.B1(n_304),
.B2(n_297),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_339),
.B(n_322),
.C(n_335),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_344),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_323),
.A2(n_326),
.B1(n_328),
.B2(n_336),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_330),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_311),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_307),
.A2(n_290),
.B1(n_293),
.B2(n_306),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_290),
.A2(n_278),
.B1(n_247),
.B2(n_255),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_276),
.B1(n_260),
.B2(n_252),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_331),
.A2(n_348),
.B1(n_281),
.B2(n_303),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_287),
.Y(n_334)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_253),
.B(n_257),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_335),
.A2(n_311),
.B(n_304),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_300),
.A2(n_276),
.B1(n_277),
.B2(n_252),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_259),
.B1(n_280),
.B2(n_267),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_349),
.B1(n_304),
.B2(n_310),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_338),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_282),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_339),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_294),
.A2(n_267),
.B1(n_273),
.B2(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_343),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_283),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_288),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_346),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_350),
.C(n_315),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_284),
.A2(n_232),
.B1(n_262),
.B2(n_229),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_294),
.A2(n_229),
.B1(n_174),
.B2(n_19),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_222),
.C(n_31),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_361),
.C(n_363),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_296),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_328),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_356),
.A2(n_358),
.B1(n_336),
.B2(n_319),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_323),
.A2(n_284),
.B1(n_305),
.B2(n_312),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_360),
.A2(n_378),
.B1(n_340),
.B2(n_322),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_315),
.C(n_289),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_289),
.C(n_313),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_368),
.C(n_369),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_302),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_363),
.Y(n_391)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_302),
.C(n_299),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_299),
.C(n_281),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_314),
.C(n_310),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_370),
.B(n_374),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_372),
.A2(n_318),
.B1(n_348),
.B2(n_331),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_381),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_285),
.C(n_304),
.Y(n_374)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_375),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_377),
.A2(n_349),
.B1(n_346),
.B2(n_345),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_326),
.A2(n_285),
.B1(n_222),
.B2(n_31),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_317),
.A2(n_31),
.B1(n_21),
.B2(n_19),
.Y(n_379)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_379),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_381),
.B(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_386),
.A2(n_387),
.B1(n_395),
.B2(n_411),
.Y(n_414)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_382),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_394),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_391),
.B(n_409),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_352),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_365),
.B(n_344),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_371),
.A2(n_319),
.B1(n_327),
.B2(n_337),
.Y(n_395)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_396),
.Y(n_433)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_397),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_327),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_401),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_399),
.A2(n_407),
.B1(n_412),
.B2(n_370),
.Y(n_415)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_353),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_376),
.B1(n_357),
.B2(n_61),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_341),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_405),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_368),
.B(n_321),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_0),
.C(n_1),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_334),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_316),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_408),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_356),
.A2(n_377),
.B1(n_371),
.B2(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_362),
.B(n_342),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_366),
.B(n_338),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_372),
.A2(n_338),
.B1(n_222),
.B2(n_44),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_377),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_384),
.A2(n_374),
.B(n_373),
.Y(n_413)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_413),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_418),
.B1(n_408),
.B2(n_2),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_398),
.A2(n_352),
.B(n_359),
.C(n_367),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_429),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_364),
.C(n_355),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_420),
.C(n_410),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_399),
.A2(n_378),
.B1(n_369),
.B2(n_362),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_380),
.C(n_359),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_422),
.B(n_423),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_383),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_431),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_46),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_46),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_2),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_46),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_46),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_389),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_435),
.A2(n_411),
.B1(n_395),
.B2(n_412),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_436),
.A2(n_401),
.B1(n_388),
.B2(n_403),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_392),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_440),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_438),
.A2(n_452),
.B1(n_424),
.B2(n_418),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_414),
.A2(n_407),
.B1(n_412),
.B2(n_385),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_433),
.Y(n_441)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_441),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_443),
.B(n_446),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g444 ( 
.A(n_425),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_444),
.B(n_445),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_SL g445 ( 
.A(n_434),
.B(n_409),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_405),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_455),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_451),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_414),
.A2(n_436),
.B1(n_421),
.B2(n_415),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_1),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_453),
.A2(n_456),
.B(n_416),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_5),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_3),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_3),
.C(n_5),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_468),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_460),
.B(n_465),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_439),
.A2(n_427),
.B(n_426),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_461),
.A2(n_469),
.B(n_449),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_427),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_466),
.Y(n_488)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_442),
.A2(n_426),
.B(n_434),
.C(n_423),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_429),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_456),
.A2(n_432),
.B(n_430),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_471),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_447),
.A2(n_455),
.B1(n_451),
.B2(n_454),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_13),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_6),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_473),
.B(n_463),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_5),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_477),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_458),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_481),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_465),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_11),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_7),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_484),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_7),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_13),
.C(n_10),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_487),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_488),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_7),
.C(n_10),
.Y(n_487)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_471),
.C(n_459),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_499),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_488),
.A2(n_464),
.B(n_463),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_12),
.B(n_494),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_495),
.B(n_497),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_475),
.A2(n_470),
.B(n_11),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_485),
.B(n_487),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_486),
.A2(n_10),
.B(n_11),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_498),
.A2(n_483),
.B(n_480),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_503),
.B(n_505),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_498),
.B(n_483),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_504),
.A2(n_501),
.B(n_500),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_11),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_499),
.C(n_492),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_491),
.B(n_12),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_505),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_509),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_511),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_513),
.A2(n_512),
.B(n_510),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_12),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_12),
.Y(n_516)
);


endmodule