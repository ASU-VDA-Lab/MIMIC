module fake_jpeg_27050_n_266 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_266);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_16),
.B(n_28),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_28),
.B(n_27),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_20),
.B1(n_26),
.B2(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_26),
.B1(n_25),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_34),
.B1(n_40),
.B2(n_30),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_25),
.B1(n_32),
.B2(n_23),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_37),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_18),
.B1(n_27),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_58),
.B1(n_43),
.B2(n_34),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_19),
.B1(n_24),
.B2(n_30),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_33),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_50),
.C(n_35),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_68),
.B1(n_80),
.B2(n_30),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_51),
.B1(n_34),
.B2(n_57),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_44),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_52),
.B1(n_48),
.B2(n_56),
.Y(n_100)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_52),
.B1(n_45),
.B2(n_31),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_34),
.B1(n_40),
.B2(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_21),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_108),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_50),
.C(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_98),
.C(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_48),
.C(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_52),
.B1(n_58),
.B2(n_49),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_85),
.B1(n_81),
.B2(n_84),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_67),
.C(n_63),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_73),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_64),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_106),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_61),
.B(n_24),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_35),
.C(n_30),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_75),
.B1(n_78),
.B2(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_65),
.B(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_29),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_68),
.B(n_63),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_125),
.B(n_127),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_118),
.B(n_125),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_135),
.B1(n_140),
.B2(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_130),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_84),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_12),
.B(n_15),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_99),
.B1(n_8),
.B2(n_10),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_29),
.B(n_31),
.C(n_7),
.D(n_11),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_108),
.A3(n_102),
.B1(n_97),
.B2(n_8),
.C1(n_5),
.C2(n_6),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_78),
.C(n_82),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_137),
.C(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_82),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_74),
.B1(n_31),
.B2(n_29),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_144),
.B(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_150),
.C(n_128),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_94),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_114),
.C(n_101),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_103),
.B(n_93),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_158),
.B(n_10),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_12),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_161),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_113),
.A3(n_108),
.B1(n_89),
.B2(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_162),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_106),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_102),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_106),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_128),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_90),
.B1(n_31),
.B2(n_29),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_164),
.B1(n_160),
.B2(n_169),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_190),
.B1(n_154),
.B2(n_31),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_128),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_177),
.C(n_188),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_129),
.B1(n_141),
.B2(n_142),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_187),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_179),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_122),
.B1(n_119),
.B2(n_109),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_119),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_90),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_166),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_31),
.C(n_29),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_152),
.C(n_145),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_144),
.B1(n_170),
.B2(n_159),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_198),
.B1(n_200),
.B2(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_203),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_157),
.B1(n_167),
.B2(n_163),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_148),
.B(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_207),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_180),
.B1(n_185),
.B2(n_174),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_205),
.C(n_208),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_148),
.C(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_29),
.C(n_7),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_7),
.C(n_13),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_211),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_14),
.C(n_6),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_182),
.B1(n_184),
.B2(n_14),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_198),
.B1(n_195),
.B2(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_204),
.B(n_183),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_215),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_227),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_201),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_201),
.B(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_223),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_208),
.C(n_194),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_240),
.C(n_223),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_175),
.C(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_246),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

OAI321xp33_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_221),
.A3(n_224),
.B1(n_227),
.B2(n_219),
.C(n_11),
.Y(n_248)
);

OAI21x1_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_1),
.B(n_2),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_249),
.A2(n_239),
.B1(n_236),
.B2(n_230),
.Y(n_256)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_250),
.A2(n_249),
.B1(n_233),
.B2(n_247),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_3),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_3),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_259),
.B(n_260),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_4),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_4),
.A3(n_252),
.B1(n_246),
.B2(n_235),
.C1(n_196),
.C2(n_232),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_262),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_264),
.Y(n_265)
);

XNOR2x2_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_261),
.Y(n_266)
);


endmodule