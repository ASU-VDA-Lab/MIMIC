module fake_jpeg_15561_n_267 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_37),
.Y(n_64)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_41),
.B(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_34),
.B1(n_18),
.B2(n_19),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_63),
.B1(n_39),
.B2(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_30),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_59),
.Y(n_76)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_60),
.B(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_70),
.B1(n_76),
.B2(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_39),
.B(n_37),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_77),
.C(n_97),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_37),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_24),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_39),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_40),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_82),
.B1(n_40),
.B2(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_66),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_92),
.Y(n_121)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_42),
.A3(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_96),
.B(n_99),
.C(n_24),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_19),
.B(n_34),
.C(n_23),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_42),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_22),
.C(n_43),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_40),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_30),
.B(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_29),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_97),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_74),
.B(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_118),
.B(n_67),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_78),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_20),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_120),
.B1(n_72),
.B2(n_93),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_79),
.B1(n_83),
.B2(n_57),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_22),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_22),
.C(n_20),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_40),
.B1(n_57),
.B2(n_26),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_125),
.B1(n_67),
.B2(n_92),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_0),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_77),
.B1(n_73),
.B2(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_81),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_57),
.B1(n_66),
.B2(n_33),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_131),
.B(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_156),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_108),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_140),
.C(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_69),
.C(n_95),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_145),
.B(n_118),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_144),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_155),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_84),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_69),
.C(n_89),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_69),
.C(n_89),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_121),
.B1(n_112),
.B2(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_109),
.B(n_22),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_86),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_173),
.CI(n_156),
.CON(n_188),
.SN(n_188)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_R g173 ( 
.A1(n_148),
.A2(n_117),
.B(n_104),
.C(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_131),
.A2(n_122),
.B(n_121),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_182),
.B(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_140),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_106),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_170),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_180),
.A2(n_175),
.B1(n_179),
.B2(n_174),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_190),
.B1(n_198),
.B2(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_138),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_162),
.C(n_178),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_172),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_139),
.B1(n_142),
.B2(n_151),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_197),
.B(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_136),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_204),
.B(n_167),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_163),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

AO221x1_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_0),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_206),
.C(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_178),
.C(n_166),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_172),
.A3(n_182),
.B1(n_160),
.B2(n_173),
.C1(n_177),
.C2(n_176),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_16),
.C(n_15),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_215),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_161),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_161),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_167),
.C(n_11),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_203),
.B1(n_200),
.B2(n_194),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_228),
.B1(n_211),
.B2(n_212),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_200),
.B1(n_203),
.B2(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

AOI31xp67_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_188),
.A3(n_196),
.B(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_191),
.B1(n_186),
.B2(n_198),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_188),
.B1(n_10),
.B2(n_13),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_3),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_219),
.B1(n_14),
.B2(n_211),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_206),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_205),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_219),
.B(n_214),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_231),
.B(n_225),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_229),
.B(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_226),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_234),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_242),
.A3(n_240),
.B1(n_239),
.B2(n_223),
.C1(n_233),
.C2(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_5),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_236),
.B1(n_4),
.B2(n_5),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_3),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_238),
.C(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_251),
.A2(n_249),
.B1(n_248),
.B2(n_8),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_252),
.C(n_6),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_6),
.C(n_261),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_262),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);


endmodule