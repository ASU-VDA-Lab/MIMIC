module fake_jpeg_27054_n_312 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_312);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_23),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_49),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_34),
.B1(n_19),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_16),
.C(n_15),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_27),
.Y(n_58)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_60),
.B1(n_69),
.B2(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_61),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_68),
.Y(n_87)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_59),
.Y(n_85)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_41),
.B1(n_44),
.B2(n_49),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_41),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_19),
.B1(n_24),
.B2(n_22),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_33),
.B1(n_29),
.B2(n_36),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_38),
.B1(n_48),
.B2(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_43),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_67),
.B1(n_66),
.B2(n_58),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_50),
.B1(n_48),
.B2(n_47),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_57),
.B1(n_40),
.B2(n_70),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_20),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_57),
.B1(n_68),
.B2(n_40),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_38),
.B1(n_24),
.B2(n_14),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_38),
.B1(n_60),
.B2(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_12),
.B1(n_45),
.B2(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_68),
.C(n_58),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_97),
.C(n_100),
.Y(n_119)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_15),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_72),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_101),
.B(n_85),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_68),
.C(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_76),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_57),
.B1(n_62),
.B2(n_40),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_70),
.B1(n_59),
.B2(n_52),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_32),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_110),
.C(n_28),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_55),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_78),
.B(n_82),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_123),
.B(n_127),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_129),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_76),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_105),
.Y(n_125)
);

AOI22x1_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_73),
.B1(n_76),
.B2(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_76),
.B1(n_78),
.B2(n_82),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_133),
.B1(n_54),
.B2(n_84),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_86),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_135),
.B(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_88),
.B1(n_85),
.B2(n_86),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_85),
.B1(n_61),
.B2(n_90),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_140),
.B1(n_54),
.B2(n_20),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_71),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_85),
.B1(n_90),
.B2(n_74),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_28),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_27),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_143),
.B(n_53),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_21),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_84),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_21),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_92),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_155),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_116),
.B1(n_118),
.B2(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_164),
.B1(n_176),
.B2(n_177),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_65),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_157),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_80),
.B(n_9),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_65),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_170),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_143),
.B(n_131),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_71),
.B(n_80),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_161),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_20),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_9),
.B(n_11),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_13),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_16),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

OR2x6_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_129),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_16),
.C(n_15),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_159),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_157),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_172),
.B(n_161),
.Y(n_229)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_198),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_141),
.B1(n_142),
.B2(n_132),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_146),
.B1(n_160),
.B2(n_165),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_115),
.B1(n_142),
.B2(n_134),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_153),
.B(n_132),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_168),
.Y(n_223)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_158),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_115),
.B1(n_126),
.B2(n_15),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_13),
.B1(n_1),
.B2(n_0),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_196),
.B1(n_191),
.B2(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx4_ASAP7_75t_SL g212 ( 
.A(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_155),
.B1(n_166),
.B2(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_220),
.B1(n_222),
.B2(n_224),
.Y(n_238)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_225),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_176),
.B1(n_150),
.B2(n_147),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_190),
.B1(n_184),
.B2(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_147),
.B(n_161),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_196),
.B1(n_183),
.B2(n_181),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_178),
.C(n_168),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_228),
.C(n_193),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_173),
.C(n_170),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_225),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_246),
.B1(n_171),
.B2(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_226),
.B1(n_209),
.B2(n_218),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_219),
.C(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_244),
.C(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_188),
.C(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_188),
.C(n_195),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_185),
.B1(n_174),
.B2(n_148),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_223),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_247),
.C(n_6),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_263),
.B1(n_264),
.B2(n_242),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_220),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_214),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_260),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_207),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_256),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_217),
.B1(n_154),
.B2(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_13),
.C(n_1),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_245),
.C(n_231),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_5),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI321xp33_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_238),
.A3(n_241),
.B1(n_246),
.B2(n_233),
.C(n_234),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_254),
.B1(n_249),
.B2(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_271),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_244),
.C(n_241),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_273),
.C(n_5),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_247),
.B1(n_6),
.B2(n_2),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_7),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_0),
.C(n_1),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_253),
.B1(n_250),
.B2(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_286),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_283),
.B1(n_2),
.B2(n_3),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_285),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_7),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_7),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_2),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_270),
.C(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_11),
.B(n_4),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_276),
.C(n_275),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_284),
.C(n_4),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_296),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_302),
.B(n_303),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_4),
.B(n_9),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_4),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_294),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_300),
.C(n_301),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_293),
.C(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_10),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_10),
.B(n_1),
.Y(n_312)
);


endmodule