module fake_jpeg_15862_n_375 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_42),
.B(n_46),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_56),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_31),
.Y(n_60)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_40),
.Y(n_82)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_0),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_17),
.Y(n_77)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_27),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_75),
.B(n_10),
.CON(n_129),
.SN(n_129)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_20),
.B1(n_41),
.B2(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_76),
.A2(n_79),
.B1(n_83),
.B2(n_91),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_77),
.B(n_115),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_41),
.B1(n_36),
.B2(n_33),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_36),
.B1(n_17),
.B2(n_35),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_81),
.A2(n_129),
.B1(n_4),
.B2(n_5),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_82),
.B(n_94),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_35),
.B1(n_38),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_29),
.B1(n_25),
.B2(n_39),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_84),
.A2(n_122),
.B1(n_127),
.B2(n_87),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_35),
.B1(n_62),
.B2(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_98),
.B(n_112),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_17),
.B1(n_24),
.B2(n_34),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_118),
.B1(n_121),
.B2(n_74),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_24),
.B1(n_38),
.B2(n_34),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_103),
.B1(n_107),
.B2(n_128),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_23),
.B1(n_32),
.B2(n_30),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_0),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_124),
.B(n_1),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_39),
.B1(n_32),
.B2(n_30),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_49),
.B(n_26),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_26),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_114),
.B(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_37),
.C(n_50),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_22),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_21),
.B1(n_37),
.B2(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_73),
.B(n_37),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_43),
.B(n_37),
.C(n_21),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_12),
.B1(n_1),
.B2(n_3),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_56),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_137),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_134),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_56),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_140),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_139),
.A2(n_171),
.B1(n_149),
.B2(n_135),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_80),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_141),
.B(n_145),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_100),
.B(n_4),
.CI(n_5),
.CON(n_142),
.SN(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_142),
.A2(n_166),
.B(n_144),
.C(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_146),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_6),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_150),
.Y(n_184)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_77),
.B(n_6),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_90),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_153),
.A2(n_167),
.B1(n_148),
.B2(n_158),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_7),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_156),
.Y(n_192)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_7),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_163),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_110),
.A2(n_8),
.B1(n_10),
.B2(n_88),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_170),
.B1(n_172),
.B2(n_175),
.Y(n_194)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_10),
.B1(n_81),
.B2(n_78),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_156),
.B(n_154),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_176),
.B1(n_181),
.B2(n_131),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_90),
.A2(n_97),
.B1(n_78),
.B2(n_93),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_81),
.A2(n_113),
.B1(n_126),
.B2(n_121),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_169),
.A2(n_176),
.B(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_93),
.B1(n_110),
.B2(n_116),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_102),
.A2(n_85),
.B1(n_124),
.B2(n_81),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_115),
.A2(n_86),
.B1(n_108),
.B2(n_97),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_86),
.A2(n_108),
.B1(n_92),
.B2(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_77),
.B(n_105),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_77),
.B(n_105),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_147),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_77),
.A2(n_122),
.B1(n_47),
.B2(n_51),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_76),
.A2(n_57),
.B1(n_62),
.B2(n_47),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_181),
.B1(n_165),
.B2(n_180),
.Y(n_205)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_191),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_201),
.B1(n_207),
.B2(n_222),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_193),
.A2(n_190),
.B1(n_201),
.B2(n_200),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_143),
.B1(n_172),
.B2(n_142),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_199),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_192),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_209),
.B1(n_146),
.B2(n_168),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_161),
.B(n_179),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_206),
.B(n_217),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_134),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_139),
.A2(n_169),
.B1(n_182),
.B2(n_155),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_142),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_143),
.A2(n_158),
.B1(n_169),
.B2(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_143),
.B(n_158),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_133),
.B(n_160),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_191),
.B1(n_214),
.B2(n_222),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_170),
.B(n_164),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_168),
.C(n_159),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_232),
.Y(n_277)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_211),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_174),
.C(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_207),
.Y(n_234)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_218),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_240),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_239),
.A2(n_185),
.B1(n_186),
.B2(n_204),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_243),
.B(n_217),
.Y(n_273)
);

NAND2x1p5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_188),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_242),
.B(n_262),
.Y(n_289)
);

AOI22x1_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_194),
.B1(n_209),
.B2(n_193),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_251),
.B1(n_188),
.B2(n_194),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_258),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_195),
.B(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_262),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_187),
.A2(n_183),
.B1(n_207),
.B2(n_208),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_254),
.A2(n_185),
.B1(n_219),
.B2(n_225),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_257),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_184),
.B(n_192),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_202),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_184),
.B(n_205),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_255),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_183),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_281),
.B1(n_242),
.B2(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_223),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_275),
.B(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_243),
.B(n_206),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_283),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_219),
.B(n_225),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_246),
.A2(n_189),
.B(n_215),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_196),
.B1(n_203),
.B2(n_215),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_196),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_245),
.B(n_203),
.Y(n_283)
);

OAI22x1_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_234),
.B1(n_257),
.B2(n_263),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_234),
.B1(n_249),
.B2(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_229),
.B(n_186),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_235),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_229),
.C(n_250),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_261),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_302),
.B1(n_306),
.B2(n_314),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_247),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_294),
.B(n_305),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_298),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_299),
.C(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_241),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_252),
.C(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_232),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_278),
.A2(n_239),
.B1(n_267),
.B2(n_281),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_304),
.A2(n_265),
.B1(n_268),
.B2(n_284),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_230),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_227),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_228),
.C(n_244),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_310),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_233),
.Y(n_310)
);

XOR2x2_ASAP7_75t_SL g313 ( 
.A(n_269),
.B(n_279),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_275),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_288),
.B1(n_272),
.B2(n_283),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_326),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_306),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_293),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_282),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_304),
.B1(n_302),
.B2(n_292),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_328),
.B1(n_330),
.B2(n_332),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_277),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_270),
.B1(n_266),
.B2(n_287),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_274),
.B1(n_270),
.B2(n_290),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_274),
.B1(n_265),
.B2(n_290),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_329),
.B(n_320),
.Y(n_338)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_342),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_300),
.B(n_311),
.C(n_298),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_327),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_344),
.B(n_345),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_332),
.B(n_266),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_303),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_347),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_310),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_326),
.C(n_323),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_356),
.C(n_353),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_341),
.B(n_330),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_354),
.B(n_355),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_323),
.C(n_299),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_349),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_344),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_359),
.B(n_361),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_334),
.Y(n_361)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_351),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_362),
.A2(n_363),
.B(n_357),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_333),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_365),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_360),
.A2(n_336),
.B1(n_348),
.B2(n_319),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g369 ( 
.A1(n_366),
.A2(n_343),
.B(n_339),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_369),
.B(n_355),
.Y(n_370)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_371),
.A3(n_367),
.B1(n_348),
.B2(n_318),
.C1(n_365),
.C2(n_335),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_368),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_372),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_373),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_364),
.Y(n_375)
);


endmodule