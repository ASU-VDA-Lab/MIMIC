module fake_jpeg_13380_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_0),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_19),
.B(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_56),
.B(n_51),
.C(n_60),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_56),
.B(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_48),
.B1(n_69),
.B2(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_61),
.B1(n_64),
.B2(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_91),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_54),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_49),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_85),
.B1(n_83),
.B2(n_82),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_109),
.B(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_108),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_25),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_104),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_100),
.Y(n_123)
);

OAI22x1_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_55),
.B1(n_74),
.B2(n_61),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_6),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_61),
.C(n_20),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_8),
.C(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_17),
.B1(n_45),
.B2(n_44),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_0),
.B(n_1),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_22),
.B1(n_43),
.B2(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_93),
.B(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_16),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_5),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_3),
.B(n_5),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_11),
.B(n_14),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_26),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_112),
.C(n_13),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_131),
.B1(n_107),
.B2(n_12),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_7),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_7),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_8),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_28),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_105),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_138),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_125),
.B1(n_133),
.B2(n_117),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_144),
.B1(n_129),
.B2(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_14),
.B1(n_15),
.B2(n_27),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_148),
.B1(n_126),
.B2(n_122),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_147),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_138),
.B(n_140),
.C(n_135),
.D(n_145),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_120),
.B(n_116),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_158),
.B(n_152),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_146),
.B(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.C(n_151),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_156),
.C(n_144),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_142),
.A3(n_115),
.B1(n_143),
.B2(n_40),
.C1(n_37),
.C2(n_47),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_123),
.Y(n_164)
);


endmodule