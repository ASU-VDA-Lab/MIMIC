module fake_jpeg_1033_n_709 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_709);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_709;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx11_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_60),
.B(n_62),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_61),
.B(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_63),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_64),
.Y(n_205)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_67),
.Y(n_169)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_69),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_84),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_80),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_27),
.B(n_9),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_92),
.Y(n_204)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_94),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_98),
.Y(n_224)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_103),
.B(n_107),
.Y(n_170)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_105),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_32),
.B(n_10),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_28),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_31),
.B(n_10),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_36),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_31),
.B(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_116),
.Y(n_176)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_42),
.B(n_7),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_122),
.Y(n_182)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_43),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_21),
.Y(n_127)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_26),
.Y(n_128)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_44),
.Y(n_130)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_46),
.Y(n_132)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_42),
.B(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_133),
.B(n_38),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_134),
.B(n_141),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_84),
.B(n_32),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_66),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_148),
.B(n_151),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_104),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_78),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_152),
.B(n_179),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_61),
.A2(n_29),
.B(n_56),
.Y(n_154)
);

OR2x2_ASAP7_75t_SL g241 ( 
.A(n_154),
.B(n_57),
.Y(n_241)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_163),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_189),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_86),
.A2(n_54),
.B1(n_46),
.B2(n_49),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_174),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_75),
.B(n_46),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_175),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_88),
.Y(n_179)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_193),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_64),
.B(n_38),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_214),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

BUFx4f_ASAP7_75t_SL g247 ( 
.A(n_200),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_69),
.B(n_28),
.Y(n_201)
);

INVx2_ASAP7_75t_R g270 ( 
.A(n_201),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_208),
.Y(n_248)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_65),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_92),
.B(n_40),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_132),
.B(n_37),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_228),
.Y(n_282)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_91),
.Y(n_219)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_81),
.B(n_49),
.C(n_54),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_220),
.B(n_54),
.C(n_52),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_80),
.B(n_49),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_98),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_231),
.Y(n_253)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_102),
.Y(n_225)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_94),
.B(n_40),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_87),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_109),
.Y(n_232)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_51),
.B1(n_30),
.B2(n_29),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_139),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_234),
.B(n_241),
.Y(n_331)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_238),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_136),
.A2(n_37),
.B(n_26),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_239),
.A2(n_242),
.B(n_212),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_51),
.B1(n_30),
.B2(n_29),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_240),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_136),
.A2(n_37),
.B(n_51),
.Y(n_242)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_244),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_245),
.B(n_304),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_139),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_246),
.B(n_252),
.Y(n_336)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_145),
.Y(n_250)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_177),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_256),
.Y(n_333)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

BUFx8_ASAP7_75t_L g375 ( 
.A(n_259),
.Y(n_375)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_146),
.A2(n_40),
.B1(n_129),
.B2(n_125),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_264),
.A2(n_278),
.B1(n_312),
.B2(n_143),
.Y(n_351)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_266),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_30),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_267),
.B(n_269),
.Y(n_337)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_221),
.A2(n_95),
.B1(n_126),
.B2(n_118),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_268),
.A2(n_293),
.B1(n_297),
.B2(n_299),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_26),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_176),
.B(n_33),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_272),
.B(n_273),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_170),
.B(n_33),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_170),
.B(n_33),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_274),
.B(n_277),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_195),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_279),
.Y(n_318)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_158),
.Y(n_276)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_178),
.B(n_184),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_146),
.A2(n_130),
.B1(n_111),
.B2(n_34),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_182),
.B(n_56),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_155),
.Y(n_280)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

CKINVDCx12_ASAP7_75t_R g281 ( 
.A(n_181),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_281),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_317),
.B1(n_219),
.B2(n_160),
.Y(n_330)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_172),
.Y(n_285)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_285),
.Y(n_347)
);

BUFx12_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

BUFx4f_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_182),
.B(n_57),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_294),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_191),
.Y(n_289)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_289),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_144),
.B(n_55),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_311),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_169),
.A2(n_55),
.B1(n_53),
.B2(n_34),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_180),
.B(n_53),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_190),
.Y(n_295)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_169),
.A2(n_53),
.B1(n_34),
.B2(n_49),
.Y(n_297)
);

CKINVDCx12_ASAP7_75t_R g298 ( 
.A(n_205),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_298),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_175),
.A2(n_54),
.B1(n_45),
.B2(n_52),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_185),
.B(n_0),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_305),
.Y(n_339)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_137),
.Y(n_301)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_194),
.Y(n_303)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_187),
.B(n_0),
.Y(n_305)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_198),
.Y(n_308)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_209),
.B(n_0),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_316),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_160),
.Y(n_310)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_223),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_167),
.A2(n_52),
.B1(n_13),
.B2(n_14),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_218),
.Y(n_313)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_150),
.B(n_13),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_315),
.Y(n_352)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_210),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_140),
.B(n_1),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_153),
.A2(n_52),
.B1(n_2),
.B2(n_3),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_323),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_163),
.B1(n_183),
.B2(n_147),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_327),
.A2(n_330),
.B1(n_361),
.B2(n_317),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_270),
.A2(n_165),
.B(n_213),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_329),
.A2(n_345),
.B(n_360),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_157),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_335),
.C(n_380),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_224),
.C(n_204),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_245),
.A2(n_138),
.B1(n_215),
.B2(n_166),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_340),
.A2(n_348),
.B1(n_360),
.B2(n_366),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_270),
.A2(n_199),
.B1(n_164),
.B2(n_171),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_344),
.A2(n_356),
.B1(n_364),
.B2(n_296),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_239),
.A2(n_135),
.B(n_156),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_245),
.A2(n_230),
.B1(n_229),
.B2(n_227),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_351),
.B(n_373),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_307),
.A2(n_192),
.B1(n_161),
.B2(n_203),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_197),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_374),
.Y(n_383)
);

OAI22x1_ASAP7_75t_L g360 ( 
.A1(n_251),
.A2(n_211),
.B1(n_194),
.B2(n_216),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_251),
.A2(n_143),
.B1(n_147),
.B2(n_202),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_294),
.A2(n_192),
.B1(n_203),
.B2(n_202),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_248),
.A2(n_216),
.B1(n_159),
.B2(n_186),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_288),
.A2(n_142),
.B1(n_223),
.B2(n_199),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_252),
.B(n_291),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_300),
.B(n_305),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_309),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_237),
.B(n_171),
.C(n_164),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_381),
.A2(n_395),
.B1(n_419),
.B2(n_427),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_370),
.B(n_242),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_382),
.B(n_392),
.Y(n_458)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_337),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_241),
.C(n_304),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_413),
.C(n_325),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_388),
.B(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_390),
.A2(n_393),
.B1(n_400),
.B2(n_402),
.Y(n_447)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_257),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_346),
.A2(n_316),
.B1(n_268),
.B2(n_161),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_292),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_399),
.Y(n_431)
);

BUFx24_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_336),
.Y(n_396)
);

INVx3_ASAP7_75t_SL g397 ( 
.A(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_318),
.B(n_253),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g399 ( 
.A1(n_319),
.A2(n_268),
.A3(n_255),
.B1(n_250),
.B2(n_236),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_346),
.A2(n_254),
.B1(n_260),
.B2(n_244),
.Y(n_400)
);

AOI221xp5_ASAP7_75t_L g401 ( 
.A1(n_331),
.A2(n_235),
.B1(n_247),
.B2(n_295),
.C(n_313),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_401),
.B(n_410),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_L g402 ( 
.A1(n_334),
.A2(n_243),
.B1(n_262),
.B2(n_280),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_367),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_420),
.Y(n_462)
);

INVx8_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_404),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_249),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_422),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_377),
.Y(n_408)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_327),
.A2(n_249),
.B1(n_258),
.B2(n_254),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_409),
.A2(n_426),
.B1(n_344),
.B2(n_356),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_319),
.B(n_332),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_355),
.A2(n_243),
.B1(n_260),
.B2(n_310),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_428),
.B1(n_247),
.B2(n_375),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_335),
.B(n_276),
.C(n_285),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_358),
.B(n_378),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_415),
.B(n_364),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_416),
.Y(n_453)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_341),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_417),
.B(n_423),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_424),
.B(n_373),
.Y(n_441)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_367),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_330),
.A2(n_258),
.B1(n_308),
.B2(n_315),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_421),
.A2(n_326),
.B1(n_347),
.B2(n_379),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_358),
.B(n_323),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_322),
.B(n_306),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_329),
.A2(n_265),
.B(n_256),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_271),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_429),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_355),
.A2(n_238),
.B1(n_263),
.B2(n_271),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_363),
.A2(n_289),
.B1(n_302),
.B2(n_263),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_363),
.A2(n_284),
.B1(n_306),
.B2(n_259),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_432),
.A2(n_446),
.B1(n_454),
.B2(n_464),
.Y(n_477)
);

OAI32xp33_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_345),
.A3(n_324),
.B1(n_325),
.B2(n_354),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_435),
.B(n_440),
.C(n_450),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_414),
.A2(n_390),
.B1(n_430),
.B2(n_418),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_438),
.A2(n_471),
.B1(n_441),
.B2(n_432),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_380),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_441),
.A2(n_397),
.B(n_371),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_388),
.B(n_361),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_443),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_354),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_425),
.Y(n_444)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_444),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_324),
.C(n_369),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_394),
.B(n_369),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_459),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_455),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_430),
.A2(n_343),
.B1(n_368),
.B2(n_320),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_333),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_368),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_383),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_460),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_399),
.B(n_362),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_472),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_396),
.A2(n_430),
.B1(n_429),
.B2(n_389),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_466),
.A2(n_386),
.B1(n_391),
.B2(n_419),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_385),
.B(n_379),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_400),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_393),
.A2(n_343),
.B1(n_320),
.B2(n_338),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_385),
.B(n_338),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_447),
.A2(n_405),
.B1(n_409),
.B2(n_424),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_474),
.A2(n_489),
.B1(n_512),
.B2(n_441),
.Y(n_516)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_475),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_450),
.C(n_506),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_372),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_484),
.B(n_365),
.Y(n_549)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_436),
.Y(n_485)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_449),
.Y(n_486)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_487),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_445),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_488),
.B(n_503),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_447),
.A2(n_402),
.B1(n_381),
.B2(n_417),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_490),
.A2(n_493),
.B1(n_495),
.B2(n_509),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_465),
.A2(n_426),
.B(n_420),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_491),
.A2(n_496),
.B(n_468),
.Y(n_536)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_492),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_431),
.A2(n_408),
.B1(n_404),
.B2(n_403),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_497),
.Y(n_524)
);

AOI32xp33_ASAP7_75t_L g498 ( 
.A1(n_431),
.A2(n_451),
.A3(n_472),
.B1(n_434),
.B2(n_437),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_498),
.B(n_452),
.Y(n_533)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_499),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_439),
.B(n_372),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_500),
.B(n_247),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_445),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_469),
.Y(n_504)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_505),
.Y(n_538)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_461),
.Y(n_507)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_507),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_463),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_433),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_434),
.A2(n_448),
.B1(n_442),
.B2(n_444),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_421),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_457),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_459),
.B(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_511),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_456),
.A2(n_416),
.B1(n_411),
.B2(n_376),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_376),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_513),
.A2(n_458),
.B1(n_454),
.B2(n_455),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_513),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_515),
.B(n_531),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_516),
.A2(n_525),
.B1(n_549),
.B2(n_476),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_478),
.B(n_491),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_519),
.A2(n_536),
.B(n_542),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_435),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_522),
.B(n_534),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_478),
.A2(n_495),
.B1(n_501),
.B2(n_489),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_527),
.B(n_552),
.Y(n_553)
);

AOI21xp33_ASAP7_75t_L g572 ( 
.A1(n_533),
.A2(n_475),
.B(n_504),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_479),
.B(n_440),
.Y(n_534)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_535),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_537),
.B(n_548),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_511),
.Y(n_539)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_488),
.B(n_438),
.Y(n_540)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_540),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_461),
.Y(n_541)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_541),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_471),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_467),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_543),
.B(n_353),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_474),
.B(n_457),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_546),
.A2(n_476),
.B1(n_477),
.B2(n_499),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_483),
.B(n_453),
.Y(n_547)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_547),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_502),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_483),
.B(n_453),
.Y(n_550)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_550),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_326),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_347),
.Y(n_584)
);

XNOR2x1_ASAP7_75t_L g605 ( 
.A(n_554),
.B(n_546),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_522),
.B(n_510),
.C(n_482),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_555),
.B(n_566),
.C(n_575),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_556),
.A2(n_546),
.B1(n_526),
.B2(n_536),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_525),
.A2(n_516),
.B1(n_519),
.B2(n_535),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_557),
.A2(n_565),
.B1(n_583),
.B2(n_546),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_529),
.A2(n_494),
.B1(n_497),
.B2(n_480),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_558),
.A2(n_554),
.B1(n_564),
.B2(n_563),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_492),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_559),
.B(n_579),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_528),
.A2(n_480),
.B1(n_486),
.B2(n_485),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_512),
.C(n_507),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_570),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_534),
.B(n_487),
.Y(n_571)
);

MAJx2_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_580),
.C(n_585),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_530),
.Y(n_574)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_574),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_551),
.B(n_505),
.C(n_357),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_523),
.B(n_357),
.C(n_321),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_521),
.C(n_532),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_547),
.B(n_481),
.Y(n_577)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_577),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_545),
.B(n_321),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_SL g580 ( 
.A(n_540),
.B(n_266),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_582),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_545),
.A2(n_473),
.B1(n_416),
.B2(n_365),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_584),
.B(n_587),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_524),
.B(n_473),
.Y(n_585)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_524),
.B(n_375),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_604),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_541),
.C(n_539),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_593),
.B(n_594),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_578),
.B(n_550),
.C(n_523),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_559),
.B(n_520),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_596),
.B(n_598),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_518),
.Y(n_597)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_597),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_553),
.B(n_555),
.C(n_571),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_599),
.A2(n_609),
.B1(n_365),
.B2(n_395),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_566),
.B(n_517),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_600),
.B(n_560),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_553),
.B(n_542),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_602),
.B(n_606),
.Y(n_618)
);

FAx1_ASAP7_75t_L g604 ( 
.A(n_569),
.B(n_557),
.CI(n_580),
.CON(n_604),
.SN(n_604)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_605),
.B(n_604),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_SL g606 ( 
.A(n_568),
.B(n_542),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_526),
.C(n_521),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_610),
.C(n_612),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_544),
.C(n_538),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_585),
.B(n_562),
.C(n_587),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_615),
.A2(n_581),
.B1(n_579),
.B2(n_583),
.Y(n_620)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_616),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_604),
.A2(n_569),
.B(n_558),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_617),
.B(n_625),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_593),
.B(n_561),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_637),
.Y(n_651)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_620),
.Y(n_645)
);

MAJx2_ASAP7_75t_L g659 ( 
.A(n_621),
.B(n_636),
.C(n_12),
.Y(n_659)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_613),
.Y(n_624)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_624),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_588),
.B(n_581),
.C(n_576),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_588),
.B(n_544),
.C(n_538),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_626),
.Y(n_652)
);

BUFx24_ASAP7_75t_SL g627 ( 
.A(n_611),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_627),
.B(n_614),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_532),
.C(n_353),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_629),
.B(n_634),
.C(n_52),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_630),
.B(n_605),
.Y(n_640)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_589),
.Y(n_632)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_632),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_598),
.B(n_591),
.C(n_594),
.Y(n_634)
);

AOI322xp5_ASAP7_75t_L g635 ( 
.A1(n_595),
.A2(n_395),
.A3(n_284),
.B1(n_407),
.B2(n_287),
.C1(n_259),
.C2(n_194),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_635),
.B(n_639),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_SL g636 ( 
.A(n_590),
.B(n_395),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_612),
.B(n_287),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_602),
.B(n_303),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_638),
.B(n_52),
.Y(n_657)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_592),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_640),
.A2(n_648),
.B1(n_649),
.B2(n_638),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_642),
.B(n_650),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_603),
.Y(n_644)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_644),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_621),
.A2(n_607),
.B(n_606),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_646),
.A2(n_5),
.B(n_17),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_631),
.A2(n_590),
.B1(n_610),
.B2(n_601),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_631),
.A2(n_628),
.B1(n_623),
.B2(n_619),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_633),
.B(n_301),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_622),
.A2(n_261),
.B1(n_211),
.B2(n_14),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_654),
.A2(n_656),
.B1(n_3),
.B2(n_4),
.Y(n_675)
);

AOI31xp33_ASAP7_75t_L g656 ( 
.A1(n_634),
.A2(n_261),
.A3(n_13),
.B(n_15),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_657),
.B(n_658),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_659),
.B(n_636),
.Y(n_661)
);

XNOR2xp5_ASAP7_75t_L g678 ( 
.A(n_661),
.B(n_666),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_652),
.B(n_625),
.C(n_622),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_662),
.B(n_664),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_641),
.B(n_629),
.C(n_637),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_643),
.Y(n_665)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_665),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_645),
.A2(n_618),
.B1(n_13),
.B2(n_15),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_667),
.B(n_668),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_655),
.A2(n_618),
.B1(n_6),
.B2(n_16),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_1),
.C(n_2),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_669),
.B(n_672),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_670),
.B(n_659),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_649),
.A2(n_5),
.B1(n_17),
.B2(n_16),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g683 ( 
.A1(n_671),
.A2(n_640),
.B1(n_657),
.B2(n_17),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_651),
.B(n_1),
.C(n_2),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_651),
.B(n_1),
.C(n_2),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_674),
.B(n_644),
.C(n_648),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_675),
.B(n_653),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_673),
.A2(n_646),
.B(n_640),
.C(n_647),
.Y(n_676)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_676),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_677),
.B(n_680),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_681),
.B(n_683),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_662),
.B(n_3),
.C(n_5),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g693 ( 
.A(n_684),
.B(n_672),
.C(n_660),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_666),
.A2(n_18),
.B(n_665),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_685),
.A2(n_669),
.B(n_674),
.Y(n_692)
);

AOI21x1_ASAP7_75t_SL g689 ( 
.A1(n_676),
.A2(n_687),
.B(n_661),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_SL g698 ( 
.A1(n_689),
.A2(n_678),
.B(n_681),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_SL g690 ( 
.A1(n_686),
.A2(n_671),
.B1(n_663),
.B2(n_664),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_690),
.B(n_691),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_682),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_692),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_693),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_698),
.B(n_660),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_694),
.A2(n_695),
.B(n_688),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_699),
.A2(n_689),
.B(n_690),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_701),
.A2(n_703),
.B(n_696),
.Y(n_705)
);

AOI322xp5_ASAP7_75t_L g702 ( 
.A1(n_700),
.A2(n_679),
.A3(n_678),
.B1(n_680),
.B2(n_683),
.C1(n_693),
.C2(n_684),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_702),
.Y(n_704)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_705),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_706),
.B(n_697),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_707),
.A2(n_704),
.B(n_18),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_708),
.A2(n_18),
.B(n_700),
.Y(n_709)
);


endmodule