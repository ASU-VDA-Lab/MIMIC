module fake_jpeg_21749_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_17),
.B1(n_22),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_50),
.B1(n_47),
.B2(n_40),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_22),
.B1(n_17),
.B2(n_33),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_85),
.B1(n_89),
.B2(n_96),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_73),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_74),
.B(n_79),
.CI(n_82),
.CON(n_131),
.SN(n_131)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_21),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_32),
.B1(n_27),
.B2(n_22),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_37),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_84),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_32),
.B1(n_27),
.B2(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_32),
.B1(n_33),
.B2(n_27),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_36),
.B1(n_42),
.B2(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_106),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_45),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_41),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_31),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_34),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_35),
.B1(n_33),
.B2(n_36),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_111),
.B1(n_42),
.B2(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_110),
.B1(n_31),
.B2(n_30),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_35),
.B1(n_31),
.B2(n_39),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_130),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_114),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_42),
.B1(n_35),
.B2(n_30),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_98),
.B1(n_76),
.B2(n_86),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_41),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_20),
.B(n_19),
.C(n_18),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_43),
.B1(n_41),
.B2(n_19),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_96),
.B1(n_78),
.B2(n_91),
.Y(n_148)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_71),
.A2(n_43),
.B1(n_41),
.B2(n_20),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_92),
.B1(n_80),
.B2(n_18),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_82),
.B1(n_107),
.B2(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_146),
.B1(n_173),
.B2(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_82),
.B1(n_93),
.B2(n_84),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_166),
.B1(n_169),
.B2(n_134),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_88),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_170),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_84),
.C(n_90),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_158),
.C(n_113),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_165),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_100),
.B(n_87),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_153),
.B(n_171),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_106),
.B(n_28),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_76),
.B1(n_90),
.B2(n_29),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_156),
.B1(n_121),
.B2(n_125),
.Y(n_200)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_18),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_43),
.C(n_83),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

BUFx24_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_163),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_113),
.B(n_28),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_34),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_34),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_121),
.B1(n_124),
.B2(n_115),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_160),
.B1(n_146),
.B2(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_188),
.B1(n_198),
.B2(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_136),
.B1(n_141),
.B2(n_128),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_135),
.B(n_139),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_152),
.B(n_153),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_192),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_149),
.B(n_115),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_137),
.B1(n_124),
.B2(n_134),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_167),
.B1(n_117),
.B2(n_138),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_196),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_125),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_117),
.B1(n_138),
.B2(n_26),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_167),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_209),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_172),
.B(n_171),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_158),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_175),
.B(n_190),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_169),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_223),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_103),
.B(n_75),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_230),
.A2(n_232),
.B1(n_181),
.B2(n_226),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_180),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_188),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_26),
.A3(n_24),
.B1(n_11),
.B2(n_75),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_183),
.A2(n_26),
.B1(n_24),
.B2(n_83),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_227),
.B1(n_203),
.B2(n_230),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_202),
.C(n_193),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_199),
.C(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_199),
.C(n_179),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_194),
.B1(n_185),
.B2(n_177),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_224),
.B1(n_227),
.B2(n_229),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_252),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_197),
.C(n_178),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_215),
.C(n_212),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_248),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_221),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_184),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_182),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_213),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_203),
.C(n_83),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_224),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_270),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_228),
.C(n_225),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_277),
.C(n_245),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_225),
.B(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_253),
.B1(n_220),
.B2(n_242),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_210),
.B1(n_232),
.B2(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_276),
.B1(n_236),
.B2(n_253),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_235),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_208),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_247),
.A2(n_220),
.B1(n_234),
.B2(n_217),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_246),
.C(n_252),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_239),
.B(n_255),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_284),
.B(n_0),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_249),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_283),
.Y(n_294)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_285),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_249),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_239),
.B(n_245),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_254),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_287),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_262),
.B1(n_277),
.B2(n_264),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_11),
.B1(n_1),
.B2(n_3),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_272),
.B1(n_271),
.B2(n_273),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_297),
.B1(n_299),
.B2(n_304),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_276),
.B1(n_262),
.B2(n_275),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_303),
.B1(n_295),
.B2(n_283),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_264),
.B1(n_203),
.B2(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_24),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_292),
.C(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_301),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_284),
.B(n_279),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_4),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_0),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_281),
.C(n_282),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_294),
.B(n_281),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_302),
.B(n_295),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_309),
.B(n_311),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_314),
.B(n_316),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_321),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_310),
.B1(n_5),
.B2(n_6),
.Y(n_324)
);

OAI211xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_5),
.C(n_7),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_8),
.B(n_9),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_8),
.Y(n_330)
);


endmodule