module fake_jpeg_647_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_12),
.B(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_36),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_40),
.B1(n_32),
.B2(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_65),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_59),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_33),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_0),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_32),
.C(n_13),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_14),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_64),
.C(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_71),
.B(n_73),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_89),
.C(n_90),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_59),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_92),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_11),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_15),
.C(n_23),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_10),
.C(n_22),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_82),
.B(n_87),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_86),
.C(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_94),
.Y(n_105)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_85),
.A3(n_16),
.B1(n_18),
.B2(n_29),
.C(n_9),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_4),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_103),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_106),
.B(n_100),
.Y(n_108)
);

NAND4xp25_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_96),
.C(n_6),
.D(n_7),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_5),
.B(n_6),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_7),
.Y(n_111)
);


endmodule