module fake_jpeg_28256_n_262 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_19),
.B1(n_16),
.B2(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_41),
.B1(n_44),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_44)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_54),
.B1(n_58),
.B2(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_51),
.Y(n_70)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_26),
.B1(n_38),
.B2(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_21),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_62),
.B1(n_38),
.B2(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_38),
.B2(n_43),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_42),
.B1(n_40),
.B2(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_79),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_16),
.B1(n_46),
.B2(n_39),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_28),
.C(n_33),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_68),
.C(n_73),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_42),
.B1(n_46),
.B2(n_39),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_50),
.B1(n_47),
.B2(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_99),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_59),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_82),
.B(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_100),
.B1(n_81),
.B2(n_65),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_60),
.B1(n_62),
.B2(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_67),
.Y(n_111)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_62),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_60),
.B1(n_51),
.B2(n_28),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_33),
.C(n_34),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_80),
.C(n_55),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_113),
.C(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_91),
.B1(n_97),
.B2(n_74),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_112),
.B(n_115),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_80),
.C(n_75),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_82),
.B(n_80),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_72),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_102),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_115),
.B(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_77),
.C(n_34),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_18),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_66),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_127),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_129),
.B(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_89),
.B1(n_84),
.B2(n_96),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_139),
.B1(n_140),
.B2(n_69),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_85),
.B(n_12),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_85),
.B(n_12),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_37),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_142),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_74),
.A3(n_71),
.B1(n_12),
.B2(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_109),
.B1(n_103),
.B2(n_104),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_107),
.B1(n_105),
.B2(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_153),
.B1(n_162),
.B2(n_15),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_55),
.C(n_76),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_158),
.C(n_163),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_156),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_55),
.C(n_69),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_0),
.B(n_1),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_15),
.B1(n_13),
.B2(n_25),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_37),
.C(n_23),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_129),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_10),
.B(n_9),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_141),
.B(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_169),
.Y(n_202)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_124),
.B1(n_136),
.B2(n_135),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_173),
.B1(n_177),
.B2(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_124),
.B1(n_131),
.B2(n_125),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_134),
.C(n_138),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_179),
.C(n_183),
.Y(n_190)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_37),
.C(n_23),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_24),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_186),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_37),
.C(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_9),
.C(n_13),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_162),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_24),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_163),
.C(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_180),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_192),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_153),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_160),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_155),
.C(n_152),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_155),
.C(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_154),
.C(n_149),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_154),
.B(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_149),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_167),
.C(n_177),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_0),
.CI(n_1),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_175),
.C(n_169),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_213),
.C(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_172),
.C(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_176),
.B1(n_181),
.B2(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_181),
.C(n_23),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_196),
.B1(n_198),
.B2(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_199),
.B1(n_187),
.B2(n_24),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_224),
.B1(n_0),
.B2(n_1),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_209),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_227),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_24),
.B1(n_22),
.B2(n_9),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_18),
.C(n_22),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_228),
.C(n_2),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_64),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_206),
.C(n_217),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_22),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_0),
.B(n_1),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_237),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_64),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_225),
.B(n_229),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_236),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_228),
.C(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.C(n_3),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_219),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_243),
.B(n_2),
.Y(n_249)
);

AOI31xp33_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_229),
.A3(n_226),
.B(n_238),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_250),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_252),
.B(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_3),
.C(n_4),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_4),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_251),
.A2(n_242),
.B1(n_6),
.B2(n_7),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_253),
.B(n_251),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_8),
.B(n_5),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_5),
.C(n_6),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_5),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_6),
.B1(n_8),
.B2(n_171),
.Y(n_262)
);


endmodule