module fake_jpeg_31071_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_2),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_44),
.B1(n_34),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_23),
.B1(n_30),
.B2(n_9),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_63),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_36),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_43),
.A3(n_41),
.B1(n_35),
.B2(n_24),
.Y(n_67)
);

OR2x4_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_36),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_73),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_3),
.B(n_4),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_31),
.B1(n_20),
.B2(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_5),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_7),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_25),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_26),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_13),
.C(n_14),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_72),
.B1(n_17),
.B2(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_89),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_100),
.B(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_103),
.B1(n_80),
.B2(n_84),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_84),
.B(n_90),
.C(n_80),
.D(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_96),
.B(n_93),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_97),
.B(n_19),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_15),
.C(n_27),
.Y(n_108)
);


endmodule