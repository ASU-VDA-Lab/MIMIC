module fake_jpeg_29375_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_36),
.C(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_18),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_29),
.B1(n_25),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_61),
.B1(n_75),
.B2(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_31),
.B1(n_37),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_70),
.B1(n_77),
.B2(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_31),
.B1(n_37),
.B2(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_66),
.B(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_25),
.B1(n_20),
.B2(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_39),
.A2(n_20),
.B1(n_26),
.B2(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_86),
.Y(n_98)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_24),
.B1(n_26),
.B2(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_27),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_40),
.A2(n_32),
.B1(n_30),
.B2(n_19),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_52),
.B1(n_23),
.B2(n_3),
.Y(n_119)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_101),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_19),
.B1(n_17),
.B2(n_23),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_107),
.Y(n_136)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_17),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_113),
.Y(n_144)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_40),
.B1(n_32),
.B2(n_53),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_53),
.B1(n_49),
.B2(n_32),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_0),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_123),
.Y(n_139)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_1),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_85),
.B1(n_87),
.B2(n_67),
.Y(n_143)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_60),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_128),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_68),
.B(n_63),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_109),
.B(n_110),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_68),
.B(n_11),
.C(n_12),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_131),
.B(n_147),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_15),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_144),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_155),
.B(n_135),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_95),
.A2(n_65),
.B1(n_87),
.B2(n_79),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_141),
.A2(n_161),
.B1(n_162),
.B2(n_97),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_155),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_91),
.A2(n_83),
.B1(n_67),
.B2(n_52),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_128),
.B1(n_100),
.B2(n_111),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_84),
.C(n_85),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_154),
.C(n_108),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_158),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_84),
.C(n_23),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_101),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_23),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_84),
.B1(n_11),
.B2(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_106),
.A2(n_107),
.B1(n_96),
.B2(n_122),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_172),
.B(n_178),
.Y(n_215)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_110),
.B(n_100),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_174),
.B(n_149),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_173),
.B1(n_191),
.B2(n_192),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_181),
.Y(n_205)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_111),
.B1(n_124),
.B2(n_126),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_118),
.B(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_176),
.B(n_179),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_118),
.C(n_92),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_130),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_187),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_140),
.B(n_148),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_90),
.C(n_92),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_137),
.C(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_104),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_175),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_138),
.A2(n_114),
.B1(n_93),
.B2(n_123),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_158),
.B(n_157),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_143),
.B1(n_156),
.B2(n_133),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_121),
.B1(n_116),
.B2(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_146),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_189),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_144),
.C(n_131),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_156),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_209),
.C(n_214),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_207),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_157),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_168),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_210),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_146),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_171),
.B(n_172),
.Y(n_237)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_12),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_10),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_165),
.B(n_10),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_15),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_226),
.B1(n_212),
.B2(n_219),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_229),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_241),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_191),
.B1(n_172),
.B2(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_192),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_237),
.A2(n_197),
.B(n_219),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_170),
.B1(n_179),
.B2(n_166),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_247),
.B1(n_250),
.B2(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_167),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_227),
.C(n_205),
.Y(n_254)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_174),
.B1(n_186),
.B2(n_177),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_248),
.B1(n_245),
.B2(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_184),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_225),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_169),
.B1(n_164),
.B2(n_5),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_255),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_200),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_214),
.C(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_263),
.C(n_268),
.Y(n_285)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_215),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_202),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_259),
.A2(n_261),
.B1(n_264),
.B2(n_271),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_234),
.B1(n_233),
.B2(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_201),
.C(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_234),
.B1(n_233),
.B2(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_212),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_2),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_224),
.B1(n_197),
.B2(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_280),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_251),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_244),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_250),
.B1(n_228),
.B2(n_239),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_268),
.B1(n_273),
.B2(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_283),
.B(n_286),
.Y(n_303)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_237),
.B1(n_247),
.B2(n_252),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_241),
.B1(n_13),
.B2(n_6),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_235),
.C(n_10),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_254),
.C(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

AO221x1_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_7),
.B1(n_8),
.B2(n_14),
.C(n_15),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_16),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_260),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_299),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_264),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_257),
.C(n_14),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_289),
.C(n_281),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_7),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_288),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_314),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_305),
.C(n_293),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_298),
.C(n_291),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_316),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_285),
.B(n_297),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_324),
.B(n_325),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_299),
.B(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_279),
.C(n_277),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_326),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_312),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_329),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_317),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_318),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_308),
.B(n_307),
.C(n_302),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_313),
.C(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_322),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_330),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.C(n_335),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_332),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_328),
.B1(n_277),
.B2(n_325),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_7),
.B(n_2),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_3),
.Y(n_342)
);


endmodule