module fake_jpeg_24948_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_18),
.A2(n_25),
.B1(n_27),
.B2(n_21),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_19),
.B1(n_16),
.B2(n_4),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_52),
.B1(n_20),
.B2(n_19),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_31),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_40),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_22),
.C(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_64),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_50),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_39),
.B1(n_31),
.B2(n_32),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_65),
.B1(n_74),
.B2(n_77),
.Y(n_87)
);

OR2x4_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_69),
.C(n_13),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_68),
.Y(n_89)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_20),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_5),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_1),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_79),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_2),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_41),
.A3(n_50),
.B1(n_45),
.B2(n_10),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_90),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_50),
.B(n_8),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_88),
.C(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_7),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_56),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_8),
.A3(n_11),
.B1(n_13),
.B2(n_57),
.Y(n_93)
);

NOR4xp25_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_56),
.C(n_59),
.D(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_11),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_90),
.B1(n_83),
.B2(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_69),
.B1(n_59),
.B2(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_86),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_104),
.B(n_102),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_109),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_101),
.C(n_113),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_116),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_85),
.B(n_89),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_87),
.B1(n_92),
.B2(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_127),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_126),
.C(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_123),
.C(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_115),
.C(n_105),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_124),
.C(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_103),
.B1(n_112),
.B2(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_120),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_138),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_145),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.C(n_136),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_117),
.B(n_123),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_132),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_132),
.B(n_133),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_139),
.B(n_120),
.Y(n_161)
);

NOR4xp25_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_146),
.C(n_145),
.D(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_159),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_125),
.B1(n_135),
.B2(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_155),
.C(n_156),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_164),
.B(n_165),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_166),
.Y(n_169)
);


endmodule