module fake_jpeg_9837_n_59 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_59);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_40),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_48),
.C(n_47),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_34),
.B1(n_36),
.B2(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_33),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_31),
.B2(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_21),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_29),
.B1(n_22),
.B2(n_26),
.Y(n_58)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_44),
.C(n_35),
.Y(n_59)
);


endmodule