module fake_jpeg_6460_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_1),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_44),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_15),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_1),
.B(n_2),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_43),
.B(n_17),
.C(n_22),
.Y(n_73)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_64)
);

BUFx2_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_20),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_52),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_31),
.B1(n_24),
.B2(n_15),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_57),
.B1(n_89),
.B2(n_90),
.Y(n_119)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_58),
.B(n_68),
.Y(n_122)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx11_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_69),
.Y(n_110)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_77),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_96),
.B(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_23),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_23),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_92),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_19),
.B1(n_32),
.B2(n_26),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_33),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_94),
.B1(n_30),
.B2(n_20),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g94 ( 
.A(n_40),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_24),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_41),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_122),
.B1(n_116),
.B2(n_118),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_21),
.B(n_24),
.C(n_30),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_111),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_108),
.A2(n_7),
.B(n_8),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_51),
.A2(n_24),
.B(n_30),
.C(n_20),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_64),
.B1(n_67),
.B2(n_60),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_164)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_132),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_57),
.B(n_55),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_133),
.B(n_153),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_54),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_54),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_135),
.Y(n_177)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_137),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_52),
.Y(n_138)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_141),
.Y(n_181)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_64),
.B1(n_60),
.B2(n_62),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_31),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_62),
.B1(n_91),
.B2(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_78),
.B1(n_68),
.B2(n_63),
.Y(n_148)
);

OAI22x1_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_63),
.B1(n_24),
.B2(n_31),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_150),
.B1(n_109),
.B2(n_113),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_117),
.B1(n_110),
.B2(n_121),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_6),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_7),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_100),
.B(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_9),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_172),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_109),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_123),
.B1(n_132),
.B2(n_12),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_98),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_98),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_110),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_176),
.B(n_126),
.Y(n_199)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_182),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_101),
.Y(n_176)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_135),
.B1(n_128),
.B2(n_141),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_99),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_134),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_99),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_189),
.Y(n_222)
);

OAI221xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_144),
.B1(n_140),
.B2(n_151),
.C(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_126),
.B(n_143),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_199),
.B(n_166),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

AO221x1_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_178),
.B1(n_158),
.B2(n_176),
.C(n_161),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_147),
.B1(n_125),
.B2(n_121),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_154),
.A3(n_123),
.B1(n_121),
.B2(n_13),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_182),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_207),
.B1(n_165),
.B2(n_168),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_160),
.C(n_167),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_216),
.C(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_213),
.B(n_215),
.Y(n_226)
);

AOI21x1_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_164),
.B(n_171),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_217),
.B(n_219),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_166),
.C(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_175),
.C(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_221),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_165),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_205),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_238),
.B(n_221),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_216),
.C(n_224),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_196),
.C(n_199),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.C(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_205),
.C(n_203),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_206),
.B1(n_207),
.B2(n_191),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_193),
.B1(n_201),
.B2(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_245),
.C(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_247),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_219),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_244),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_222),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_219),
.C(n_209),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_234),
.B1(n_231),
.B2(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_183),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_173),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_229),
.C(n_233),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_248),
.B(n_233),
.Y(n_261)
);

AOI31xp67_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_226),
.A3(n_238),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_232),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_161),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_262),
.B(n_212),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_261),
.A2(n_259),
.B(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_163),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_265),
.B1(n_168),
.B2(n_253),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_266),
.C(n_185),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_258),
.A2(n_251),
.B(n_225),
.Y(n_266)
);

OAI31xp33_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_251),
.A3(n_253),
.B(n_173),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_268),
.Y(n_272)
);


endmodule