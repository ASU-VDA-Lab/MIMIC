module real_jpeg_23448_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_36),
.B1(n_65),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_1),
.A2(n_36),
.B1(n_60),
.B2(n_171),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_3),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_64),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_3),
.A2(n_68),
.B(n_84),
.C(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_3),
.A2(n_65),
.B1(n_68),
.B2(n_172),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_3),
.B(n_29),
.C(n_46),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_3),
.A2(n_41),
.B1(n_43),
.B2(n_172),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_3),
.A2(n_26),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_126),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_5),
.A2(n_41),
.B1(n_43),
.B2(n_62),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_62),
.Y(n_192)
);

INVx8_ASAP7_75t_SL g67 ( 
.A(n_6),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_7),
.A2(n_61),
.B1(n_73),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_7),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_65),
.B1(n_68),
.B2(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_41),
.B1(n_43),
.B2(n_111),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_111),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_10),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_10),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_41),
.B1(n_43),
.B2(n_75),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_10),
.A2(n_65),
.B1(n_68),
.B2(n_75),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_75),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_41),
.B1(n_43),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_51),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_11),
.A2(n_51),
.B1(n_65),
.B2(n_68),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_11),
.A2(n_51),
.B1(n_58),
.B2(n_61),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_12),
.A2(n_65),
.B1(n_68),
.B2(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_12),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_12),
.A2(n_41),
.B1(n_43),
.B2(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_12),
.A2(n_61),
.B1(n_88),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_88),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_13),
.A2(n_65),
.B1(n_68),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_162),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_13),
.A2(n_41),
.B1(n_43),
.B2(n_162),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_162),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_40),
.B1(n_65),
.B2(n_68),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_15),
.A2(n_40),
.B1(n_73),
.B2(n_74),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_180)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_16),
.A2(n_27),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_16),
.A2(n_27),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_353),
.B(n_356),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_348),
.B(n_352),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_335),
.B(n_347),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_137),
.A3(n_151),
.B(n_332),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_115),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_22),
.B(n_115),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.C(n_95),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_23),
.A2(n_79),
.B1(n_80),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_23),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_53),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_24),
.A2(n_25),
.B(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_25),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_54),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_26),
.A2(n_35),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_26),
.A2(n_179),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_26),
.A2(n_32),
.B1(n_100),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_26),
.A2(n_261),
.B(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_27),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_29),
.B1(n_46),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_28),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_33),
.B(n_172),
.Y(n_265)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_39),
.A2(n_44),
.B1(n_52),
.B2(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_43),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_41),
.B(n_253),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_43),
.A2(n_85),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_44),
.A2(n_52),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_44),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_44),
.A2(n_52),
.B1(n_227),
.B2(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_49),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_49),
.A2(n_91),
.B1(n_105),
.B2(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_49),
.B(n_172),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_49),
.A2(n_167),
.B(n_242),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_52),
.B(n_168),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B(n_70),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_57),
.A2(n_63),
.B1(n_112),
.B2(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_58),
.Y(n_171)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g183 ( 
.A(n_59),
.B(n_67),
.C(n_68),
.Y(n_183)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_72),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_63),
.A2(n_112),
.B1(n_134),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_63),
.A2(n_70),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_64),
.A2(n_77),
.B1(n_110),
.B2(n_204),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_64),
.A2(n_77),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_64),
.A2(n_77),
.B1(n_343),
.B2(n_350),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_64),
.A2(n_77),
.B(n_350),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_68),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_65),
.A2(n_69),
.B(n_173),
.C(n_183),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_69),
.B1(n_73),
.B2(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_74),
.B(n_172),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_77),
.A2(n_114),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_94),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_82),
.A2(n_83),
.B1(n_128),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_82),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_82),
.A2(n_201),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_83),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_83),
.A2(n_107),
.B(n_187),
.Y(n_311)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_91),
.A2(n_226),
.B(n_228),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_91),
.A2(n_228),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_95),
.A2(n_96),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.C(n_108),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_97),
.A2(n_98),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_99),
.Y(n_304)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_101),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_101),
.A2(n_235),
.B(n_259),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_106),
.B(n_108),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_118),
.C(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_133),
.B2(n_136),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_126),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_125),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_125),
.A2(n_126),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_126),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_130),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_130),
.B(n_144),
.C(n_148),
.Y(n_346)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_136),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_133),
.B(n_140),
.C(n_143),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_138),
.A2(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_150),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_139),
.B(n_150),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_145),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_149),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_325),
.B(n_331),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_315),
.B(n_324),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_213),
.B(n_298),
.C(n_314),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_196),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_155),
.B(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_174),
.C(n_184),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_156),
.A2(n_157),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_164),
.C(n_169),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_174),
.A2(n_175),
.B1(n_184),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_181),
.B2(n_182),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_181),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_191),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_212),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_197),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.CI(n_202),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_210),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_291),
.B(n_297),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_246),
.B(n_290),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_238),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_218),
.B(n_238),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_237),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_225),
.C(n_229),
.Y(n_296)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.C(n_243),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_284),
.B(n_289),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_274),
.B(n_283),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_262),
.B(n_273),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_257),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_269),
.B(n_272),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_282),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_282),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_288),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_296),
.Y(n_297)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_313),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_313),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_303),
.C(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_310),
.C(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_320),
.C(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_337),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_341),
.B1(n_344),
.B2(n_345),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_339),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_341),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_344),
.C(n_346),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_351),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_354),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_349),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_355),
.B(n_358),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_357),
.Y(n_356)
);


endmodule