module real_aes_507_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_789;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g553 ( .A(n_0), .B(n_193), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_1), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g124 ( .A(n_2), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_3), .B(n_485), .Y(n_484) );
NAND2xp33_ASAP7_75t_SL g539 ( .A(n_4), .B(n_153), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_5), .B(n_133), .Y(n_184) );
INVx1_ASAP7_75t_L g532 ( .A(n_6), .Y(n_532) );
INVx1_ASAP7_75t_L g230 ( .A(n_7), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g771 ( .A(n_8), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_9), .Y(n_244) );
AND2x2_ASAP7_75t_L g482 ( .A(n_10), .B(n_172), .Y(n_482) );
INVx2_ASAP7_75t_L g132 ( .A(n_11), .Y(n_132) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_12), .Y(n_466) );
INVx1_ASAP7_75t_L g194 ( .A(n_13), .Y(n_194) );
AOI221x1_ASAP7_75t_L g535 ( .A1(n_14), .A2(n_158), .B1(n_487), .B2(n_536), .C(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_15), .B(n_485), .Y(n_522) );
INVx1_ASAP7_75t_L g469 ( .A(n_16), .Y(n_469) );
INVx1_ASAP7_75t_L g191 ( .A(n_17), .Y(n_191) );
INVx1_ASAP7_75t_SL g177 ( .A(n_18), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_19), .B(n_144), .Y(n_143) );
AOI33xp33_ASAP7_75t_L g210 ( .A1(n_20), .A2(n_52), .A3(n_121), .B1(n_139), .B2(n_211), .B3(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_21), .A2(n_487), .B(n_488), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_22), .B(n_193), .Y(n_489) );
AOI221xp5_ASAP7_75t_SL g543 ( .A1(n_23), .A2(n_40), .B1(n_485), .B2(n_487), .C(n_544), .Y(n_543) );
AOI22x1_ASAP7_75t_R g751 ( .A1(n_24), .A2(n_36), .B1(n_752), .B2(n_753), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_24), .Y(n_753) );
INVx1_ASAP7_75t_L g238 ( .A(n_25), .Y(n_238) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_26), .A2(n_91), .B(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g134 ( .A(n_26), .B(n_91), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_27), .B(n_196), .Y(n_526) );
INVxp67_ASAP7_75t_L g534 ( .A(n_28), .Y(n_534) );
AND2x2_ASAP7_75t_L g508 ( .A(n_29), .B(n_171), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_30), .B(n_165), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_31), .A2(n_487), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_32), .B(n_196), .Y(n_545) );
AND2x2_ASAP7_75t_L g127 ( .A(n_33), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
AND2x2_ASAP7_75t_L g153 ( .A(n_33), .B(n_124), .Y(n_153) );
OR2x6_ASAP7_75t_L g467 ( .A(n_34), .B(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_35), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_36), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_37), .B(n_165), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_38), .A2(n_118), .B1(n_130), .B2(n_133), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_39), .B(n_150), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_41), .A2(n_82), .B1(n_136), .B2(n_487), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_42), .B(n_144), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_43), .Y(n_761) );
XOR2xp5_ASAP7_75t_L g108 ( .A(n_44), .B(n_109), .Y(n_108) );
AOI22x1_ASAP7_75t_SL g785 ( .A1(n_44), .A2(n_68), .B1(n_786), .B2(n_787), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_44), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_45), .B(n_193), .Y(n_506) );
XNOR2x2_ASAP7_75t_SL g750 ( .A(n_46), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_47), .B(n_155), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_48), .B(n_144), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_49), .Y(n_129) );
AND2x2_ASAP7_75t_L g556 ( .A(n_50), .B(n_171), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_51), .B(n_171), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_53), .B(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_54), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g122 ( .A(n_55), .Y(n_122) );
INVx1_ASAP7_75t_L g146 ( .A(n_55), .Y(n_146) );
AND2x2_ASAP7_75t_L g223 ( .A(n_56), .B(n_171), .Y(n_223) );
AOI221xp5_ASAP7_75t_L g228 ( .A1(n_57), .A2(n_75), .B1(n_136), .B2(n_165), .C(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_58), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_59), .B(n_485), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_60), .B(n_130), .Y(n_246) );
AOI21xp5_ASAP7_75t_SL g160 ( .A1(n_61), .A2(n_136), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g499 ( .A(n_62), .B(n_171), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_63), .B(n_196), .Y(n_554) );
INVx1_ASAP7_75t_L g187 ( .A(n_64), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_65), .B(n_193), .Y(n_497) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_66), .B(n_172), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_67), .A2(n_487), .B(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_68), .Y(n_787) );
INVx1_ASAP7_75t_L g221 ( .A(n_69), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_70), .B(n_196), .Y(n_490) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_71), .B(n_155), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_72), .A2(n_136), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g128 ( .A(n_73), .Y(n_128) );
INVx1_ASAP7_75t_L g148 ( .A(n_73), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_74), .B(n_165), .Y(n_213) );
AND2x2_ASAP7_75t_L g179 ( .A(n_76), .B(n_158), .Y(n_179) );
INVx1_ASAP7_75t_L g188 ( .A(n_77), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_78), .A2(n_136), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_79), .A2(n_136), .B(n_142), .C(n_154), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_80), .B(n_485), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_81), .A2(n_85), .B1(n_165), .B2(n_485), .Y(n_515) );
INVx1_ASAP7_75t_L g470 ( .A(n_83), .Y(n_470) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_84), .B(n_158), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_86), .A2(n_136), .B1(n_208), .B2(n_209), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_87), .B(n_193), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_88), .B(n_193), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_89), .A2(n_104), .B1(n_764), .B2(n_775), .C1(n_793), .C2(n_797), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_89), .A2(n_780), .B1(n_781), .B2(n_790), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_89), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_90), .A2(n_487), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_93), .B(n_196), .Y(n_496) );
AND2x2_ASAP7_75t_L g214 ( .A(n_94), .B(n_158), .Y(n_214) );
OAI22xp33_ASAP7_75t_SL g783 ( .A1(n_95), .A2(n_784), .B1(n_785), .B2(n_788), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_95), .Y(n_788) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_96), .A2(n_236), .B(n_237), .C(n_239), .Y(n_235) );
INVxp67_ASAP7_75t_L g537 ( .A(n_97), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_98), .B(n_485), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_99), .B(n_196), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_100), .A2(n_487), .B(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g772 ( .A(n_101), .Y(n_772) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_101), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_102), .B(n_144), .Y(n_163) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI21xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_750), .B(n_754), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_464), .B1(n_471), .B2(n_473), .Y(n_107) );
INVx1_ASAP7_75t_L g759 ( .A(n_108), .Y(n_759) );
AO22x1_ASAP7_75t_L g781 ( .A1(n_109), .A2(n_782), .B1(n_783), .B2(n_789), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_109), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g109 ( .A(n_110), .B(n_315), .C(n_381), .D(n_444), .Y(n_109) );
NOR2x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_278), .Y(n_110) );
OR3x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_248), .C(n_275), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_180), .B(n_203), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_166), .Y(n_114) );
AND2x2_ASAP7_75t_L g378 ( .A(n_115), .B(n_348), .Y(n_378) );
INVx1_ASAP7_75t_L g451 ( .A(n_115), .Y(n_451) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_156), .Y(n_115) );
INVx2_ASAP7_75t_L g202 ( .A(n_116), .Y(n_202) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_116), .Y(n_266) );
AND2x2_ASAP7_75t_L g270 ( .A(n_116), .B(n_183), .Y(n_270) );
AND2x4_ASAP7_75t_L g286 ( .A(n_116), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g290 ( .A(n_116), .Y(n_290) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_135), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_125), .C(n_129), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g165 ( .A(n_120), .B(n_126), .Y(n_165) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
OR2x6_ASAP7_75t_L g151 ( .A(n_121), .B(n_140), .Y(n_151) );
INVxp33_ASAP7_75t_L g211 ( .A(n_121), .Y(n_211) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g141 ( .A(n_122), .B(n_124), .Y(n_141) );
AND2x4_ASAP7_75t_L g196 ( .A(n_122), .B(n_147), .Y(n_196) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_L g487 ( .A(n_127), .B(n_141), .Y(n_487) );
INVx2_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
AND2x6_ASAP7_75t_L g193 ( .A(n_128), .B(n_145), .Y(n_193) );
INVx4_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_130), .B(n_243), .Y(n_242) );
AOI21x1_ASAP7_75t_L g549 ( .A1(n_130), .A2(n_550), .B(n_556), .Y(n_549) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx4f_ASAP7_75t_L g155 ( .A(n_131), .Y(n_155) );
AND2x4_ASAP7_75t_L g133 ( .A(n_132), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_132), .B(n_134), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_133), .A2(n_160), .B(n_164), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_133), .B(n_152), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_133), .A2(n_484), .B(n_486), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_133), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_133), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_133), .B(n_537), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_133), .B(n_189), .C(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_L g245 ( .A(n_136), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_136), .A2(n_165), .B1(n_531), .B2(n_533), .Y(n_530) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NOR2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_149), .B(n_152), .Y(n_142) );
INVx1_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
AND2x4_ASAP7_75t_L g485 ( .A(n_144), .B(n_153), .Y(n_485) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_151), .A2(n_152), .B(n_162), .C(n_163), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_151), .A2(n_152), .B(n_177), .C(n_178), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_151), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_151), .A2(n_152), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_SL g229 ( .A1(n_151), .A2(n_152), .B(n_230), .C(n_231), .Y(n_229) );
INVxp67_ASAP7_75t_L g236 ( .A(n_151), .Y(n_236) );
INVx1_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_152), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_152), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_152), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_152), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_152), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_152), .A2(n_553), .B(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_153), .Y(n_239) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_154), .A2(n_206), .B(n_214), .Y(n_205) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_154), .A2(n_206), .B(n_214), .Y(n_254) );
AOI21x1_ASAP7_75t_L g513 ( .A1(n_154), .A2(n_514), .B(n_517), .Y(n_513) );
INVx2_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_155), .A2(n_228), .B(n_232), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_155), .A2(n_522), .B(n_523), .Y(n_521) );
AND2x2_ASAP7_75t_L g181 ( .A(n_156), .B(n_182), .Y(n_181) );
INVx4_ASAP7_75t_L g267 ( .A(n_156), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_156), .B(n_257), .Y(n_271) );
INVx2_ASAP7_75t_L g285 ( .A(n_156), .Y(n_285) );
AND2x4_ASAP7_75t_L g289 ( .A(n_156), .B(n_290), .Y(n_289) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_156), .Y(n_324) );
OR2x2_ASAP7_75t_L g330 ( .A(n_156), .B(n_169), .Y(n_330) );
NOR2x1_ASAP7_75t_SL g359 ( .A(n_156), .B(n_183), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_156), .B(n_433), .Y(n_461) );
OR2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx3_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_158), .A2(n_216), .B1(n_235), .B2(n_240), .Y(n_234) );
INVx1_ASAP7_75t_L g247 ( .A(n_165), .Y(n_247) );
AND2x2_ASAP7_75t_L g358 ( .A(n_166), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2x1_ASAP7_75t_L g392 ( .A(n_167), .B(n_182), .Y(n_392) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
INVx2_ASAP7_75t_L g258 ( .A(n_169), .Y(n_258) );
AND2x2_ASAP7_75t_L g281 ( .A(n_169), .B(n_183), .Y(n_281) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_169), .Y(n_308) );
INVx1_ASAP7_75t_L g349 ( .A(n_169), .Y(n_349) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_179), .Y(n_169) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_170), .A2(n_493), .B(n_499), .Y(n_492) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_170), .A2(n_502), .B(n_508), .Y(n_501) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_170), .A2(n_502), .B(n_508), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_171), .A2(n_543), .B(n_547), .Y(n_542) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_198), .Y(n_180) );
AND2x2_ASAP7_75t_L g361 ( .A(n_181), .B(n_256), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_182), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g428 ( .A(n_182), .Y(n_428) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g287 ( .A(n_183), .Y(n_287) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_190), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_189), .B(n_238), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B1(n_194), .B2(n_195), .Y(n_190) );
INVxp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_198), .A2(n_365), .B(n_369), .C(n_375), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_200), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_SL g411 ( .A(n_200), .Y(n_411) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g333 ( .A(n_202), .B(n_287), .Y(n_333) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_224), .Y(n_203) );
AOI32xp33_ASAP7_75t_L g369 ( .A1(n_204), .A2(n_353), .A3(n_370), .B1(n_371), .B2(n_373), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
INVx2_ASAP7_75t_L g295 ( .A(n_205), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_205), .B(n_227), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_213), .Y(n_206) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g307 ( .A(n_215), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_215), .B(n_233), .Y(n_338) );
AND2x2_ASAP7_75t_L g343 ( .A(n_215), .B(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_215), .Y(n_425) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_223), .Y(n_215) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_217), .B(n_223), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
OR2x2_ASAP7_75t_L g326 ( .A(n_224), .B(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g277 ( .A(n_225), .B(n_251), .Y(n_277) );
AND2x2_ASAP7_75t_L g426 ( .A(n_225), .B(n_424), .Y(n_426) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_233), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g263 ( .A(n_227), .Y(n_263) );
AND2x4_ASAP7_75t_L g302 ( .A(n_227), .B(n_303), .Y(n_302) );
INVxp67_ASAP7_75t_L g336 ( .A(n_227), .Y(n_336) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_227), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_227), .B(n_233), .Y(n_353) );
INVx1_ASAP7_75t_L g437 ( .A(n_227), .Y(n_437) );
INVx2_ASAP7_75t_L g274 ( .A(n_233), .Y(n_274) );
INVx1_ASAP7_75t_L g301 ( .A(n_233), .Y(n_301) );
INVx1_ASAP7_75t_L g368 ( .A(n_233), .Y(n_368) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_241), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_245), .B1(n_246), .B2(n_247), .Y(n_241) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OAI32xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_259), .A3(n_264), .B1(n_268), .B2(n_272), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_250), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_251), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g352 ( .A(n_251), .B(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g377 ( .A(n_251), .Y(n_377) );
AND2x2_ASAP7_75t_L g458 ( .A(n_251), .B(n_300), .Y(n_458) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g273 ( .A(n_253), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g372 ( .A(n_253), .B(n_295), .Y(n_372) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_253), .B(n_274), .Y(n_394) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_253), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
INVx1_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
AND2x2_ASAP7_75t_L g342 ( .A(n_254), .B(n_274), .Y(n_342) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g370 ( .A(n_256), .B(n_359), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_256), .B(n_289), .Y(n_440) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_257), .Y(n_409) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_258), .Y(n_391) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_293), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_261), .B(n_377), .Y(n_376) );
NOR2xp67_ASAP7_75t_SL g463 ( .A(n_261), .B(n_401), .Y(n_463) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g320 ( .A(n_263), .B(n_274), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_264), .B(n_330), .Y(n_388) );
INVx2_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_265), .B(n_281), .Y(n_354) );
AND2x4_ASAP7_75t_SL g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2x1_ASAP7_75t_L g313 ( .A(n_267), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g419 ( .A(n_267), .B(n_290), .Y(n_419) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_267), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_268), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g390 ( .A(n_269), .B(n_391), .Y(n_390) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_269), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g379 ( .A(n_270), .B(n_324), .Y(n_379) );
INVxp33_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g293 ( .A(n_273), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g453 ( .A(n_273), .B(n_335), .Y(n_453) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_296), .Y(n_278) );
OAI21xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_282), .B(n_291), .Y(n_279) );
AND2x2_ASAP7_75t_L g414 ( .A(n_281), .B(n_289), .Y(n_414) );
NAND2xp33_ASAP7_75t_R g282 ( .A(n_283), .B(n_288), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g456 ( .A(n_285), .Y(n_456) );
INVx4_ASAP7_75t_L g314 ( .A(n_286), .Y(n_314) );
INVx1_ASAP7_75t_L g433 ( .A(n_287), .Y(n_433) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g427 ( .A(n_289), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_289), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_292), .A2(n_357), .B1(n_461), .B2(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g321 ( .A(n_295), .B(n_307), .Y(n_321) );
AND2x2_ASAP7_75t_L g335 ( .A(n_295), .B(n_336), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_304), .B(n_309), .C(n_312), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g383 ( .A(n_299), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g311 ( .A(n_300), .Y(n_311) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g371 ( .A(n_301), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g380 ( .A(n_301), .B(n_302), .Y(n_380) );
INVx1_ASAP7_75t_L g412 ( .A(n_301), .Y(n_412) );
AND2x4_ASAP7_75t_L g393 ( .A(n_302), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g415 ( .A(n_302), .B(n_306), .Y(n_415) );
AND2x2_ASAP7_75t_L g423 ( .A(n_302), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g398 ( .A(n_306), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_306), .B(n_320), .Y(n_400) );
AND2x2_ASAP7_75t_L g403 ( .A(n_306), .B(n_353), .Y(n_403) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_307), .B(n_368), .Y(n_417) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_333), .Y(n_345) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g441 ( .A(n_311), .B(n_321), .Y(n_441) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_313), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g325 ( .A(n_314), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_314), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_355), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_339), .Y(n_316) );
OAI222xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B1(n_326), .B2(n_328), .C1(n_331), .C2(n_334), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_SL g332 ( .A(n_324), .B(n_333), .Y(n_332) );
OR2x6_ASAP7_75t_L g404 ( .A(n_324), .B(n_374), .Y(n_404) );
NAND5xp2_ASAP7_75t_L g407 ( .A(n_324), .B(n_327), .C(n_343), .D(n_408), .E(n_410), .Y(n_407) );
NAND2x1_ASAP7_75t_L g443 ( .A(n_325), .B(n_329), .Y(n_443) );
INVx2_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
NOR2x1_ASAP7_75t_L g373 ( .A(n_330), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_332), .A2(n_423), .B1(n_426), .B2(n_427), .Y(n_422) );
INVx2_ASAP7_75t_L g374 ( .A(n_333), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_333), .B(n_349), .Y(n_386) );
INVx3_ASAP7_75t_L g421 ( .A(n_334), .Y(n_421) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g366 ( .A(n_335), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g362 ( .A(n_338), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_340), .B(n_351), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B(n_346), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g350 ( .A(n_342), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_345), .A2(n_352), .B1(n_353), .B2(n_354), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_350), .Y(n_346) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_SL g432 ( .A(n_349), .B(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_364), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_379), .B2(n_380), .Y(n_375) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_405), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_387), .C(n_395), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OA21x2_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .B(n_393), .Y(n_387) );
NAND2xp33_ASAP7_75t_SL g389 ( .A(n_390), .B(n_392), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_402), .B(n_404), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_400), .C(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_399), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_429), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_413), .C(n_420), .D(n_422), .Y(n_406) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g418 ( .A(n_409), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g449 ( .A(n_412), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_416), .B2(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_418), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_434), .B(n_438), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_459), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_454), .B2(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22x1_ASAP7_75t_L g755 ( .A1(n_464), .A2(n_756), .B1(n_757), .B2(n_759), .Y(n_755) );
CKINVDCx11_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
AND2x6_ASAP7_75t_SL g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OR2x6_ASAP7_75t_SL g471 ( .A(n_466), .B(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g763 ( .A(n_466), .B(n_467), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_466), .B(n_472), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_467), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
CKINVDCx11_ASAP7_75t_R g758 ( .A(n_471), .Y(n_758) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_474), .Y(n_756) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_672), .Y(n_474) );
NOR3xp33_ASAP7_75t_SL g475 ( .A(n_476), .B(n_596), .C(n_646), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_576), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_518), .B(n_557), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_509), .Y(n_479) );
INVx1_ASAP7_75t_SL g682 ( .A(n_480), .Y(n_682) );
AOI32xp33_ASAP7_75t_L g713 ( .A1(n_480), .A2(n_695), .A3(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_480), .B(n_572), .Y(n_715) );
AND2x4_ASAP7_75t_SL g480 ( .A(n_481), .B(n_491), .Y(n_480) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_481), .Y(n_510) );
INVx5_ASAP7_75t_L g575 ( .A(n_481), .Y(n_575) );
OR2x2_ASAP7_75t_L g582 ( .A(n_481), .B(n_574), .Y(n_582) );
INVx2_ASAP7_75t_L g587 ( .A(n_481), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_481), .B(n_492), .Y(n_599) );
AND2x2_ASAP7_75t_L g604 ( .A(n_481), .B(n_500), .Y(n_604) );
OR2x2_ASAP7_75t_L g611 ( .A(n_481), .B(n_512), .Y(n_611) );
AND2x4_ASAP7_75t_L g620 ( .A(n_481), .B(n_501), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_SL g662 ( .A1(n_481), .A2(n_578), .B(n_613), .C(n_651), .Y(n_662) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx3_ASAP7_75t_SL g612 ( .A(n_491), .Y(n_612) );
AND2x2_ASAP7_75t_L g658 ( .A(n_491), .B(n_575), .Y(n_658) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .Y(n_491) );
AND2x2_ASAP7_75t_L g511 ( .A(n_492), .B(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g589 ( .A(n_492), .B(n_501), .Y(n_589) );
AND2x2_ASAP7_75t_L g593 ( .A(n_492), .B(n_572), .Y(n_593) );
INVx1_ASAP7_75t_L g619 ( .A(n_492), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_492), .B(n_501), .Y(n_641) );
INVx2_ASAP7_75t_L g645 ( .A(n_492), .Y(n_645) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_492), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_492), .B(n_575), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g656 ( .A(n_501), .B(n_512), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .Y(n_502) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g666 ( .A(n_510), .Y(n_666) );
NAND2xp33_ASAP7_75t_SL g691 ( .A(n_510), .B(n_583), .Y(n_691) );
AND2x2_ASAP7_75t_L g733 ( .A(n_511), .B(n_575), .Y(n_733) );
AND2x2_ASAP7_75t_L g644 ( .A(n_512), .B(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g707 ( .A(n_512), .Y(n_707) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_513), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_518), .A2(n_598), .B1(n_700), .B2(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_540), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_519), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_519), .B(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .Y(n_519) );
INVx2_ASAP7_75t_L g563 ( .A(n_520), .Y(n_563) );
OR2x2_ASAP7_75t_L g567 ( .A(n_520), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_520), .B(n_580), .Y(n_585) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_520), .B(n_529), .Y(n_595) );
OR2x2_ASAP7_75t_L g602 ( .A(n_520), .B(n_542), .Y(n_602) );
OR2x2_ASAP7_75t_L g614 ( .A(n_520), .B(n_529), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_520), .B(n_542), .Y(n_628) );
INVx1_ASAP7_75t_L g633 ( .A(n_520), .Y(n_633) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_520), .Y(n_651) );
AND2x2_ASAP7_75t_L g714 ( .A(n_520), .B(n_634), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_520), .Y(n_718) );
OR2x2_ASAP7_75t_L g725 ( .A(n_520), .B(n_615), .Y(n_725) );
OR2x2_ASAP7_75t_L g747 ( .A(n_520), .B(n_748), .Y(n_747) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .Y(n_520) );
AND2x2_ASAP7_75t_L g564 ( .A(n_528), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_528), .B(n_548), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_528), .B(n_624), .Y(n_686) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g583 ( .A(n_529), .Y(n_583) );
AND2x4_ASAP7_75t_L g634 ( .A(n_529), .B(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_529), .B(n_579), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_529), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_529), .B(n_568), .Y(n_727) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AND2x2_ASAP7_75t_L g594 ( .A(n_540), .B(n_595), .Y(n_594) );
AO221x1_ASAP7_75t_L g668 ( .A1(n_540), .A2(n_583), .B1(n_614), .B2(n_669), .C(n_670), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g720 ( .A1(n_540), .A2(n_640), .A3(n_721), .B1(n_723), .B2(n_724), .C1(n_725), .C2(n_726), .Y(n_720) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_548), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g562 ( .A(n_542), .Y(n_562) );
INVx2_ASAP7_75t_L g568 ( .A(n_542), .Y(n_568) );
AND2x2_ASAP7_75t_L g580 ( .A(n_542), .B(n_548), .Y(n_580) );
INVx1_ASAP7_75t_L g625 ( .A(n_542), .Y(n_625) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_542), .Y(n_681) );
INVx1_ASAP7_75t_L g565 ( .A(n_548), .Y(n_565) );
OR2x2_ASAP7_75t_L g615 ( .A(n_548), .B(n_568), .Y(n_615) );
INVx2_ASAP7_75t_L g635 ( .A(n_548), .Y(n_635) );
INVx1_ASAP7_75t_L g688 ( .A(n_548), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_548), .B(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI21xp33_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_566), .B(n_569), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_559), .A2(n_598), .B1(n_600), .B2(n_604), .C(n_605), .Y(n_597) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
NOR2x1p5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g684 ( .A(n_563), .Y(n_684) );
INVx1_ASAP7_75t_SL g603 ( .A(n_564), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g708 ( .A1(n_564), .A2(n_709), .B(n_711), .Y(n_708) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_568), .Y(n_671) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_571), .A2(n_647), .B(n_652), .C(n_663), .Y(n_646) );
OR2x2_ASAP7_75t_L g736 ( .A(n_571), .B(n_641), .Y(n_736) );
AND2x2_ASAP7_75t_L g738 ( .A(n_571), .B(n_604), .Y(n_738) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g578 ( .A(n_572), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g640 ( .A(n_572), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g678 ( .A(n_572), .B(n_645), .Y(n_678) );
OA33x2_ASAP7_75t_L g685 ( .A1(n_572), .A2(n_602), .A3(n_686), .B1(n_687), .B2(n_689), .B3(n_691), .Y(n_685) );
OR2x2_ASAP7_75t_L g696 ( .A(n_572), .B(n_681), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_572), .B(n_620), .Y(n_710) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g598 ( .A(n_574), .B(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_574), .A2(n_604), .B1(n_648), .B2(n_649), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_575), .B(n_655), .C(n_688), .Y(n_687) );
AOI322xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .A3(n_583), .B1(n_584), .B2(n_586), .C1(n_590), .C2(n_594), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g683 ( .A(n_579), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_580), .A2(n_595), .B(n_639), .C(n_642), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_581), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND4xp25_ASAP7_75t_SL g702 ( .A(n_582), .B(n_611), .C(n_703), .D(n_705), .Y(n_702) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g592 ( .A(n_587), .Y(n_592) );
OR2x2_ASAP7_75t_L g637 ( .A(n_587), .B(n_589), .Y(n_637) );
AND2x2_ASAP7_75t_L g706 ( .A(n_588), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g711 ( .A(n_592), .B(n_706), .Y(n_711) );
BUFx2_ASAP7_75t_L g704 ( .A(n_593), .Y(n_704) );
INVx1_ASAP7_75t_SL g734 ( .A(n_594), .Y(n_734) );
AND2x4_ASAP7_75t_L g670 ( .A(n_595), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g723 ( .A(n_595), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_616), .C(n_638), .Y(n_596) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_SL g660 ( .A(n_602), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g728 ( .A1(n_602), .A2(n_729), .B(n_730), .C(n_739), .Y(n_728) );
OR2x2_ASAP7_75t_L g650 ( .A(n_603), .B(n_651), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B1(n_612), .B2(n_613), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_607), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_610), .B(n_667), .Y(n_749) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g724 ( .A(n_611), .B(n_612), .Y(n_724) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g669 ( .A(n_615), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_621), .B1(n_626), .B2(n_630), .C1(n_631), .C2(n_636), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_619), .Y(n_630) );
AND2x2_ASAP7_75t_L g677 ( .A(n_620), .B(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_620), .A2(n_693), .B1(n_698), .B2(n_702), .Y(n_692) );
INVx2_ASAP7_75t_SL g745 ( .A(n_620), .Y(n_745) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g701 ( .A(n_625), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_625), .B(n_688), .Y(n_748) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g661 ( .A(n_629), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_631), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g699 ( .A(n_633), .Y(n_699) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_634), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g742 ( .A(n_634), .B(n_671), .Y(n_742) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g667 ( .A(n_641), .Y(n_667) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g746 ( .A(n_644), .Y(n_746) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_657), .B(n_659), .C(n_662), .Y(n_652) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g697 ( .A(n_659), .Y(n_697) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_712), .C(n_728), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_692), .C(n_708), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B1(n_682), .B2(n_683), .C(n_685), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g721 ( .A(n_707), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g729 ( .A(n_711), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_719), .Y(n_712) );
INVx2_ASAP7_75t_L g735 ( .A(n_714), .Y(n_735) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g726 ( .A(n_717), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B1(n_735), .B2(n_736), .C(n_737), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_743), .B1(n_747), .B2(n_749), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g754 ( .A1(n_750), .A2(n_755), .B(n_760), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
BUFx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_773), .Y(n_766) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_769), .B(n_772), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OR2x2_ASAP7_75t_SL g796 ( .A(n_770), .B(n_772), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_770), .A2(n_799), .B(n_802), .Y(n_798) );
INVx1_ASAP7_75t_SL g792 ( .A(n_773), .Y(n_792) );
BUFx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
BUFx3_ASAP7_75t_L g778 ( .A(n_774), .Y(n_778) );
BUFx2_ASAP7_75t_L g803 ( .A(n_774), .Y(n_803) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI21x1_ASAP7_75t_SL g776 ( .A1(n_777), .A2(n_779), .B(n_791), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g789 ( .A(n_783), .Y(n_789) );
CKINVDCx16_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
CKINVDCx11_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
CKINVDCx8_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
endmodule