module fake_jpeg_9593_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_18),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_28),
.C(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_33),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_23),
.B1(n_19),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_40),
.B1(n_39),
.B2(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_64),
.B1(n_22),
.B2(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_35),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_60),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_39),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_25),
.B1(n_38),
.B2(n_43),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_95),
.B(n_98),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_80),
.Y(n_109)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_88),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_40),
.B(n_26),
.C(n_27),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_91),
.B(n_20),
.C(n_17),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_17),
.B(n_20),
.C(n_31),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_92),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_35),
.B(n_38),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_26),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_97),
.B1(n_65),
.B2(n_54),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_34),
.B1(n_31),
.B2(n_20),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_34),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_31),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_53),
.C(n_54),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_116),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_115),
.B1(n_128),
.B2(n_92),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_118),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_53),
.C(n_44),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

BUFx16f_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_84),
.A2(n_57),
.B1(n_55),
.B2(n_31),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_105),
.B1(n_116),
.B2(n_127),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_91),
.B(n_81),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_132),
.A2(n_142),
.B(n_107),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_138),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_144),
.B1(n_148),
.B2(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_82),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_90),
.B(n_86),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_103),
.B1(n_87),
.B2(n_96),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_69),
.B1(n_101),
.B2(n_96),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_110),
.B1(n_102),
.B2(n_107),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_151),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_71),
.B1(n_79),
.B2(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_98),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_74),
.B1(n_100),
.B2(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_98),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_159),
.C(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_96),
.C(n_85),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_160),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_185),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_108),
.B1(n_124),
.B2(n_119),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_176),
.B1(n_179),
.B2(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_173),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_175),
.C(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_111),
.C(n_131),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_137),
.B1(n_157),
.B2(n_134),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_131),
.B(n_122),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_139),
.B(n_3),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_112),
.B1(n_88),
.B2(n_89),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_155),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_139),
.CI(n_3),
.CON(n_189),
.SN(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_118),
.B1(n_97),
.B2(n_76),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_126),
.C(n_123),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_146),
.B1(n_99),
.B2(n_129),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_20),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_146),
.C(n_99),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_189),
.B(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_196),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_199),
.B(n_202),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_177),
.B(n_182),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_208),
.B1(n_192),
.B2(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_184),
.C(n_175),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_2),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_164),
.B(n_2),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_181),
.B1(n_165),
.B2(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_218),
.C(n_222),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_170),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_189),
.B1(n_204),
.B2(n_198),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_165),
.B1(n_172),
.B2(n_161),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_221),
.B1(n_226),
.B2(n_193),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_172),
.B1(n_162),
.B2(n_180),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_187),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_162),
.C(n_163),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.C(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_163),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_207),
.B1(n_191),
.B2(n_196),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_241),
.B1(n_210),
.B2(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_235),
.C(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_234),
.A2(n_240),
.B(n_215),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_194),
.C(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_190),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_236),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_189),
.B1(n_188),
.B2(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_16),
.C(n_5),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_16),
.C(n_6),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_222),
.C(n_225),
.Y(n_249)
);

AO221x1_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_252),
.Y(n_256)
);

NAND4xp25_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_220),
.C(n_224),
.D(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_250),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_4),
.C(n_9),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_10),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_231),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_247),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_242),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_261),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_248),
.B(n_11),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_10),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_258),
.B1(n_259),
.B2(n_254),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_11),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_273),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C1(n_268),
.C2(n_262),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_268),
.A3(n_274),
.B1(n_12),
.B2(n_13),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_12),
.Y(n_278)
);


endmodule