module fake_jpeg_15420_n_196 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_196);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_7),
.B(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_58),
.B1(n_62),
.B2(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_57),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx2_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_19),
.B1(n_27),
.B2(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_29),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_28),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_71),
.Y(n_105)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_68),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_34),
.B1(n_44),
.B2(n_43),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_48),
.B1(n_45),
.B2(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_74),
.B1(n_84),
.B2(n_85),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_39),
.B1(n_41),
.B2(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_78),
.Y(n_107)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_2),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_5),
.B(n_7),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_43),
.Y(n_108)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_35),
.B1(n_45),
.B2(n_37),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_38),
.B1(n_22),
.B2(n_32),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_30),
.B1(n_3),
.B2(n_5),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_32),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_16),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_38),
.B1(n_35),
.B2(n_33),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_88),
.B1(n_21),
.B2(n_16),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_21),
.B1(n_22),
.B2(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_29),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_99),
.B1(n_101),
.B2(n_104),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_109),
.Y(n_117)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_74),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_7),
.B1(n_8),
.B2(n_33),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_43),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_71),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_126),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_125),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_124),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_89),
.C(n_63),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_94),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_80),
.B(n_67),
.C(n_69),
.D(n_70),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_16),
.CI(n_18),
.CON(n_142),
.SN(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_102),
.B1(n_91),
.B2(n_111),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_69),
.B1(n_85),
.B2(n_66),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_80),
.B1(n_68),
.B2(n_82),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_78),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_99),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_65),
.B1(n_73),
.B2(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_145),
.Y(n_154)
);

NOR4xp25_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_94),
.C(n_97),
.D(n_37),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_81),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_113),
.B(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_90),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_83),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_143),
.A3(n_142),
.B1(n_136),
.B2(n_120),
.C1(n_130),
.C2(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_161),
.B1(n_132),
.B2(n_148),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_133),
.C(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_157),
.C(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_159),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_148),
.B1(n_113),
.B2(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_18),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_169),
.B(n_170),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_142),
.B(n_8),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_18),
.B(n_37),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_151),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_169),
.A2(n_156),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_156),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_167),
.A3(n_163),
.B1(n_171),
.B2(n_12),
.C1(n_9),
.C2(n_11),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_9),
.B(n_10),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_183),
.B(n_180),
.CI(n_175),
.CON(n_188),
.SN(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_188),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_167),
.B(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_182),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_187),
.B(n_182),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_190),
.Y(n_196)
);


endmodule