module fake_jpeg_22302_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_40),
.B1(n_16),
.B2(n_43),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_12),
.B(n_10),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_31),
.C(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_69),
.Y(n_93)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_64),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_27),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_81),
.B1(n_82),
.B2(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_75),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_78),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_85),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_33),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_110),
.C(n_81),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_64),
.B1(n_82),
.B2(n_40),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_105),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_101),
.B(n_112),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_34),
.B1(n_32),
.B2(n_73),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_56),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_109),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_38),
.B1(n_55),
.B2(n_35),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_50),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_55),
.B1(n_35),
.B2(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_0),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_31),
.B(n_19),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_22),
.B(n_17),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_66),
.B(n_36),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_27),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_32),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_124),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_127),
.B1(n_106),
.B2(n_89),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_22),
.B(n_17),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_128),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_84),
.B1(n_58),
.B2(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_34),
.C(n_32),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_137),
.C(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_138),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_90),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_16),
.B1(n_15),
.B2(n_49),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_34),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_112),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_143),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_164),
.B1(n_140),
.B2(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_145),
.B(n_156),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_121),
.A3(n_18),
.B1(n_28),
.B2(n_24),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_92),
.B1(n_97),
.B2(n_89),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_155),
.B1(n_163),
.B2(n_173),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_102),
.B1(n_67),
.B2(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_95),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_116),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_102),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_123),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_87),
.B1(n_49),
.B2(n_86),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_117),
.A2(n_87),
.B1(n_49),
.B2(n_84),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_168),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_86),
.C(n_85),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_171),
.C(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_174),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_36),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_73),
.B(n_23),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_29),
.B(n_28),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_95),
.B1(n_90),
.B2(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_192),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_131),
.B(n_120),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_177),
.A2(n_172),
.B(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_182),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_138),
.B(n_114),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_146),
.B(n_165),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_184),
.C(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_135),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_121),
.B1(n_124),
.B2(n_137),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_191),
.B1(n_202),
.B2(n_172),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_197),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_148),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_194),
.Y(n_215)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_130),
.B1(n_122),
.B2(n_111),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_200),
.B1(n_204),
.B2(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_65),
.C(n_61),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_145),
.A2(n_18),
.A3(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_61),
.C(n_23),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_160),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_157),
.B1(n_153),
.B2(n_163),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_162),
.B(n_29),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_29),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_24),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_155),
.A2(n_30),
.B1(n_25),
.B2(n_28),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_208),
.B(n_213),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_229),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_143),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_218),
.B(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_226),
.B1(n_228),
.B2(n_224),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_175),
.B(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_191),
.A2(n_168),
.B1(n_30),
.B2(n_29),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_202),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_179),
.A2(n_30),
.B1(n_28),
.B2(n_24),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_185),
.B1(n_206),
.B2(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_246),
.B(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_238),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_200),
.B1(n_183),
.B2(n_189),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_242),
.B1(n_245),
.B2(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_203),
.C(n_201),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_250),
.C(n_5),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_184),
.B1(n_192),
.B2(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_207),
.B(n_227),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_211),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_20),
.C(n_4),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_262),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_224),
.B1(n_212),
.B2(n_219),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_6),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_212),
.B1(n_219),
.B2(n_229),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_10),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_3),
.B(n_4),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_236),
.B(n_247),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_20),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_239),
.C(n_241),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_234),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_272),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_280),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_232),
.C(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_233),
.C(n_240),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_275),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_248),
.C(n_234),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_6),
.C(n_8),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_9),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_279),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_255),
.B1(n_265),
.B2(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_285),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_254),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_265),
.B1(n_252),
.B2(n_253),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_263),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_258),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_293),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_282),
.A2(n_272),
.B1(n_257),
.B2(n_253),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_295),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_271),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_264),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_292),
.B(n_290),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_305),
.B(n_293),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_310),
.A3(n_304),
.B1(n_290),
.B2(n_307),
.C(n_9),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_11),
.B(n_12),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_13),
.B(n_14),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_13),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_14),
.Y(n_316)
);


endmodule