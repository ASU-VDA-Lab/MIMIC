module fake_jpeg_31925_n_213 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_46),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_0),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_73),
.B1(n_76),
.B2(n_38),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_69),
.B1(n_83),
.B2(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_30),
.B1(n_25),
.B2(n_19),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_35),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_18),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_SL g80 ( 
.A(n_44),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_42),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_36),
.B(n_4),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_73),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_36),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_80),
.Y(n_125)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_38),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_112),
.B(n_111),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_99),
.B1(n_113),
.B2(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_124),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_91),
.B1(n_96),
.B2(n_90),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_96),
.B1(n_82),
.B2(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_116),
.Y(n_144)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_120),
.Y(n_145)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_109),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_68),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_101),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_63),
.B1(n_91),
.B2(n_68),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_139),
.B1(n_122),
.B2(n_106),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_67),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_79),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_64),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_143),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_61),
.B1(n_64),
.B2(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_143),
.B1(n_129),
.B2(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_105),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_100),
.B1(n_116),
.B2(n_113),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_163),
.B(n_136),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_153),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_162),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_124),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_113),
.B1(n_98),
.B2(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_118),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_164),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_152),
.B(n_160),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.C(n_155),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_177),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_126),
.B(n_125),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_133),
.B(n_134),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_134),
.C(n_130),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_153),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_152),
.B(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_152),
.B1(n_162),
.B2(n_150),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_132),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_186),
.B(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_169),
.C(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_198),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_199),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_181),
.B(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_178),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_194),
.C(n_128),
.Y(n_202)
);

OAI221xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_194),
.B1(n_147),
.B2(n_132),
.C(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_141),
.B(n_132),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_205),
.B(n_141),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_205),
.B(n_119),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_210),
.C(n_119),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_208),
.Y(n_213)
);


endmodule