module real_jpeg_19062_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_3),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_2),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_19),
.B1(n_40),
.B2(n_41),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_19),
.B1(n_44),
.B2(n_45),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_3),
.A2(n_8),
.B1(n_20),
.B2(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_25),
.B(n_28),
.C(n_146),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_97)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_8),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_28),
.B1(n_44),
.B2(n_45),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_9),
.B(n_24),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_21),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_8),
.A2(n_10),
.B(n_45),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_8),
.A2(n_41),
.B(n_50),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_10),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

BUFx3_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_102),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_100),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_85),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_15),
.B(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.C(n_68),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_16),
.B(n_62),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_61),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_17),
.A2(n_61),
.B1(n_87),
.B2(n_98),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_17),
.B(n_117),
.C(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_17),
.A2(n_61),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_17),
.A2(n_61),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_17),
.B(n_230),
.C(n_232),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B(n_26),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_18),
.A2(n_21),
.B1(n_83),
.B2(n_90),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_22),
.B(n_30),
.C(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_22),
.B(n_29),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_23),
.A2(n_49),
.B(n_50),
.C(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_50),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_24),
.A2(n_28),
.B(n_51),
.C(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_27),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_28),
.A2(n_41),
.B(n_42),
.C(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_28),
.B(n_74),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_28),
.B(n_43),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_28),
.B(n_49),
.Y(n_189)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_48),
.B2(n_60),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_34),
.A2(n_35),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_60),
.C(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_46),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_37),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_43),
.B1(n_46),
.B2(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_38),
.A2(n_43),
.B1(n_81),
.B2(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_64),
.B(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_44),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_55),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_56),
.A2(n_67),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_57),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_63),
.B(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_65),
.A2(n_88),
.B1(n_89),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_65),
.B(n_159),
.C(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_65),
.A2(n_142),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_68),
.A2(n_69),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_77),
.B(n_82),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_82),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_70),
.A2(n_78),
.B1(n_107),
.B2(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_72),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_74),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_74),
.A2(n_114),
.B(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_78),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_99),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_88),
.A2(n_89),
.B1(n_117),
.B2(n_153),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_112),
.C(n_117),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_89),
.B(n_142),
.C(n_143),
.Y(n_235)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_95),
.B(n_96),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_121),
.B(n_256),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_118),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_104),
.B(n_118),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_110),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_105),
.B(n_109),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_110),
.A2(n_111),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_112),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_113),
.A2(n_115),
.B1(n_190),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_113),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_115),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_115),
.B(n_147),
.C(n_189),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_115),
.A2(n_190),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_115),
.B(n_208),
.C(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_138),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_117),
.A2(n_128),
.B1(n_129),
.B2(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_117),
.B(n_129),
.C(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_250),
.B(n_255),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_238),
.B(n_249),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_165),
.B(n_222),
.C(n_237),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_149),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_125),
.B(n_149),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_127),
.B(n_137),
.C(n_140),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_129),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_128),
.B(n_133),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_129),
.B(n_174),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_181),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_157),
.B1(n_187),
.B2(n_191),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.C(n_158),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_158),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_221),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_215),
.B(n_220),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_205),
.B(n_214),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_193),
.B(n_204),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_184),
.B(n_192),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_176),
.B(n_183),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B(n_182),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_202),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_235),
.B2(n_236),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.C(n_236),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_235),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_246),
.C(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);


endmodule