module fake_jpeg_3109_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_45),
.B(n_75),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_51),
.Y(n_104)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_72),
.Y(n_94)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_30),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_82),
.Y(n_96)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_85),
.Y(n_108)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_17),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_45),
.B(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_93),
.B(n_127),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_29),
.B1(n_32),
.B2(n_15),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_105),
.A2(n_124),
.B1(n_20),
.B2(n_19),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_51),
.A2(n_19),
.B(n_20),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g144 ( 
.A(n_111),
.B(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_36),
.B1(n_42),
.B2(n_37),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_17),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_86),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_46),
.A2(n_34),
.B1(n_41),
.B2(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_47),
.B(n_37),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_48),
.B(n_44),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_129),
.B(n_70),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_55),
.A2(n_44),
.B1(n_41),
.B2(n_40),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_136),
.B1(n_31),
.B2(n_15),
.Y(n_137)
);

NOR2x1_ASAP7_75t_R g133 ( 
.A(n_58),
.B(n_20),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_50),
.B1(n_64),
.B2(n_66),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_92),
.B1(n_98),
.B2(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_34),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_75),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_65),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_154),
.B1(n_179),
.B2(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_138),
.B(n_152),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_104),
.Y(n_140)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_145),
.Y(n_216)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_156),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_159),
.B(n_169),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_19),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_74),
.B1(n_73),
.B2(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_22),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_164),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_163),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_96),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_69),
.C(n_80),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_168),
.C(n_131),
.Y(n_206)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_95),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_79),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_95),
.B(n_22),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_128),
.A3(n_114),
.B1(n_103),
.B2(n_123),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_49),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_94),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_112),
.A2(n_49),
.B(n_87),
.C(n_84),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_101),
.B(n_122),
.C(n_123),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_107),
.B(n_71),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_177),
.Y(n_218)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_99),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_116),
.A2(n_49),
.B1(n_63),
.B2(n_53),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_113),
.A2(n_71),
.B1(n_63),
.B2(n_53),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_144),
.B(n_173),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_183),
.A2(n_89),
.B(n_1),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_106),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_158),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_89),
.B1(n_98),
.B2(n_97),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_156),
.B1(n_158),
.B2(n_154),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_122),
.CI(n_131),
.CON(n_194),
.SN(n_194)
);

AOI32xp33_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_221),
.A3(n_178),
.B1(n_161),
.B2(n_140),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_198),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_99),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_204),
.C(n_170),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_139),
.A2(n_100),
.B(n_101),
.C(n_16),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_179),
.B1(n_146),
.B2(n_172),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_SL g204 ( 
.A(n_152),
.B(n_100),
.C(n_128),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_168),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_164),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_210),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_159),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_171),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_143),
.B(n_91),
.CI(n_118),
.CON(n_221),
.SN(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_226),
.C(n_245),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_227),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_182),
.B(n_169),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_228),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_235),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_253),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_181),
.B1(n_150),
.B2(n_137),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_148),
.B1(n_160),
.B2(n_118),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_145),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_236),
.B(n_237),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_239),
.B(n_194),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_244),
.Y(n_274)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_243),
.B(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_176),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_219),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_142),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_204),
.C(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_91),
.B1(n_151),
.B2(n_141),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_252),
.B(n_217),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_254),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_186),
.A2(n_191),
.B1(n_183),
.B2(n_184),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_0),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_258),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_187),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_211),
.B(n_208),
.C(n_194),
.D(n_188),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_259),
.A2(n_261),
.B(n_256),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_196),
.B(n_186),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_269),
.C(n_271),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_247),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_272),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_224),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_214),
.C(n_187),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_214),
.C(n_215),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_221),
.B1(n_203),
.B2(n_192),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_285),
.B1(n_3),
.B2(n_4),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_231),
.A2(n_221),
.B1(n_203),
.B2(n_199),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_278),
.B1(n_238),
.B2(n_261),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_215),
.C(n_197),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_287),
.C(n_233),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_216),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_232),
.A2(n_199),
.B1(n_190),
.B2(n_217),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_250),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_248),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_291),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_222),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_315),
.B1(n_285),
.B2(n_262),
.Y(n_333)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_250),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_265),
.Y(n_334)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_284),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_300),
.Y(n_326)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_274),
.A2(n_230),
.B1(n_252),
.B2(n_241),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_313),
.B1(n_275),
.B2(n_283),
.Y(n_342)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_304),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_308),
.Y(n_330)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_264),
.B(n_228),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_257),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_319),
.Y(n_337)
);

OAI211xp5_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_321),
.B(n_281),
.C(n_277),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_314),
.C(n_317),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_274),
.A2(n_241),
.B1(n_242),
.B2(n_254),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_241),
.C(n_216),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_280),
.A2(n_202),
.B1(n_0),
.B2(n_2),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_202),
.C(n_0),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_263),
.B(n_1),
.C(n_2),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_265),
.C(n_282),
.Y(n_339)
);

XOR2x2_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_1),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_287),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_3),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_279),
.B(n_2),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_322),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_293),
.A2(n_270),
.B1(n_260),
.B2(n_278),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_342),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_310),
.A2(n_270),
.B(n_259),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_327),
.A2(n_343),
.B(n_345),
.Y(n_368)
);

NAND2xp33_ASAP7_75t_SL g329 ( 
.A(n_297),
.B(n_289),
.Y(n_329)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_281),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_336),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_334),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_311),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_296),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_296),
.C(n_317),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_4),
.B(n_5),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_4),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_318),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_313),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_328),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_357),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_331),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_362),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_320),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_361),
.Y(n_374)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_342),
.A2(n_312),
.B(n_303),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_325),
.B(n_345),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_326),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_306),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_363),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_364),
.B(n_344),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_343),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_305),
.C(n_319),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_347),
.C(n_323),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_315),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_332),
.Y(n_380)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_371),
.B(n_379),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_359),
.A2(n_337),
.B1(n_323),
.B2(n_341),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_372),
.A2(n_367),
.B1(n_369),
.B2(n_360),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_375),
.B(n_383),
.Y(n_390)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_354),
.B(n_327),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_358),
.C(n_366),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_369),
.B(n_337),
.CI(n_339),
.CON(n_382),
.SN(n_382)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_374),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_341),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_375),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_352),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_388),
.B(n_335),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_393),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_395),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_392),
.A2(n_402),
.B(n_372),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_381),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_360),
.C(n_364),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_396),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_380),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_349),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_399),
.B(n_373),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_368),
.C(n_361),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_391),
.C(n_379),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_371),
.A2(n_365),
.B(n_368),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_403),
.A2(n_414),
.B(n_401),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_394),
.A2(n_386),
.B1(n_376),
.B2(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_408),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_411),
.C(n_348),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_410),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_387),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_384),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_382),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_413),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_382),
.B(n_324),
.Y(n_414)
);

OAI321xp33_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_402),
.A3(n_401),
.B1(n_400),
.B2(n_324),
.C(n_307),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_417),
.A2(n_421),
.B(n_14),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_422),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_8),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_424),
.C(n_405),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_8),
.B(n_9),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_9),
.C(n_11),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_9),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_427),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_408),
.C(n_12),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_11),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_429),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_420),
.B(n_416),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_424),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_436),
.Y(n_438)
);

AOI221xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_437),
.B1(n_433),
.B2(n_434),
.C(n_426),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_419),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);


endmodule