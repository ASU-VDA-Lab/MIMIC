module real_jpeg_13632_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_305, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_305;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_300;
wire n_215;
wire n_288;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_181;
wire n_102;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g107 ( 
.A(n_0),
.Y(n_107)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_3),
.A2(n_41),
.B1(n_45),
.B2(n_112),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_112),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_112),
.Y(n_206)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_6),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_6),
.A2(n_29),
.B1(n_41),
.B2(n_45),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_8),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_8),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_41),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_52),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_10),
.B(n_57),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_44),
.C(n_48),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_10),
.B(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_46),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_24),
.B(n_59),
.C(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_10),
.B(n_20),
.Y(n_185)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_92),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_90),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_82),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_82),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_74),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_16),
.A2(n_17),
.B1(n_68),
.B2(n_76),
.Y(n_300)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B(n_30),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_19),
.A2(n_72),
.B(n_73),
.Y(n_277)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_20),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_20),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_21),
.B(n_24),
.C(n_52),
.Y(n_197)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_23),
.A2(n_24),
.B1(n_59),
.B2(n_60),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_25),
.A2(n_69),
.B(n_72),
.Y(n_87)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_26),
.B(n_197),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_30),
.B(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_31),
.B(n_206),
.Y(n_216)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_53),
.B1(n_54),
.B2(n_66),
.Y(n_36)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_76),
.C(n_77),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_54),
.C(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_37),
.A2(n_66),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_37),
.A2(n_66),
.B1(n_77),
.B2(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_50),
.B(n_51),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_38),
.A2(n_116),
.B(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_39),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_39),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_39),
.B(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_41),
.B(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_45),
.A2(n_52),
.B(n_60),
.Y(n_168)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_46),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_46),
.B(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_46),
.B(n_131),
.Y(n_175)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_48),
.B(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_50),
.A2(n_163),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_62),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_56),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_61),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_57),
.B(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_57),
.A2(n_62),
.B(n_79),
.Y(n_281)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_65),
.Y(n_81)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_61),
.B(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_62),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_63),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_66),
.B(n_203),
.C(n_209),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_68),
.A2(n_76),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_69),
.B(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_71),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_73),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_74),
.A2(n_75),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_77),
.Y(n_294)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_81),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_81),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_84),
.A2(n_88),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_84),
.B(n_222),
.C(n_228),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_284),
.B(n_301),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_267),
.B(n_283),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_246),
.B(n_266),
.Y(n_94)
);

AOI321xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_212),
.A3(n_239),
.B1(n_244),
.B2(n_245),
.C(n_305),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_188),
.B(n_211),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_171),
.B(n_187),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_154),
.B(n_170),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_132),
.B(n_153),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_124),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_124),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_113),
.B1(n_114),
.B2(n_123),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_103),
.B(n_150),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_110),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_107),
.B(n_110),
.Y(n_166)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_107),
.A2(n_150),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_143),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_110),
.A2(n_199),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_116),
.B(n_130),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_121),
.C(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_146),
.B(n_152),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_140),
.B(n_145),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_144),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_149),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_156),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_162),
.C(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_163),
.B(n_175),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_165),
.A2(n_166),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_165),
.A2(n_166),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_263),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_166),
.A2(n_274),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_186),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_186),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_179),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_184),
.C(n_185),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_201),
.B2(n_202),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_194),
.C(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_200),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_233),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_233),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_220),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_221),
.C(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_235),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_243),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_248),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_265),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_261),
.B2(n_262),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_262),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_254),
.C(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_272),
.C(n_279),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_278),
.B2(n_279),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_280),
.B(n_281),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_290),
.B1(n_291),
.B2(n_295),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_288),
.C(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_296),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);


endmodule