module fake_jpeg_13544_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_37),
.B(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_20),
.B1(n_44),
.B2(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_77),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_82),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_64),
.B1(n_53),
.B2(n_61),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_53),
.B1(n_51),
.B2(n_4),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_47),
.C(n_68),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_94),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_57),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_6),
.Y(n_113)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_66),
.B(n_58),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_103),
.B(n_7),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_87),
.B1(n_50),
.B2(n_64),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_102),
.B1(n_85),
.B2(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_2),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_51),
.B1(n_66),
.B2(n_64),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_111),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_3),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_93),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_124),
.B(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_11),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_132),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_21),
.B(n_34),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_19),
.C(n_33),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_130),
.C(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_7),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_8),
.B(n_9),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_17),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_12),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_13),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_32),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_146),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_31),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_121),
.C(n_117),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_145),
.C(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_150),
.B(n_152),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_146),
.B1(n_139),
.B2(n_142),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_131),
.B1(n_118),
.B2(n_127),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_147),
.C(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_153),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_152),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_156),
.Y(n_161)
);


endmodule