module real_aes_538_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_0), .B(n_143), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_1), .A2(n_151), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_2), .B(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_3), .B(n_143), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_4), .B(n_170), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_5), .B(n_170), .Y(n_496) );
INVx1_ASAP7_75t_L g139 ( .A(n_6), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_7), .B(n_170), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_8), .Y(n_105) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_9), .A2(n_99), .B1(n_115), .B2(n_756), .C1(n_766), .C2(n_770), .Y(n_98) );
OAI22xp33_ASAP7_75t_SL g758 ( .A1(n_9), .A2(n_118), .B1(n_748), .B2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_9), .Y(n_759) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_10), .B(n_168), .Y(n_537) );
AND2x2_ASAP7_75t_L g173 ( .A(n_11), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g184 ( .A(n_12), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g130 ( .A(n_13), .Y(n_130) );
AOI221x1_ASAP7_75t_L g481 ( .A1(n_14), .A2(n_25), .B1(n_143), .B2(n_151), .C(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_15), .B(n_170), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_16), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_17), .B(n_143), .Y(n_533) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_18), .A2(n_185), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_19), .B(n_128), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_20), .B(n_170), .Y(n_470) );
AO21x1_ASAP7_75t_L g491 ( .A1(n_21), .A2(n_143), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_22), .B(n_143), .Y(n_226) );
INVx1_ASAP7_75t_L g113 ( .A(n_23), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_24), .A2(n_87), .B1(n_134), .B2(n_143), .Y(n_133) );
NAND2x1_ASAP7_75t_L g512 ( .A(n_26), .B(n_170), .Y(n_512) );
NAND2x1_ASAP7_75t_L g544 ( .A(n_27), .B(n_168), .Y(n_544) );
OR2x2_ASAP7_75t_L g131 ( .A(n_28), .B(n_84), .Y(n_131) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_28), .A2(n_84), .B(n_130), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_29), .B(n_168), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_30), .B(n_170), .Y(n_536) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_31), .A2(n_174), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_32), .B(n_168), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_33), .A2(n_151), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_34), .B(n_170), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_35), .A2(n_151), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g141 ( .A(n_36), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g149 ( .A(n_36), .B(n_139), .Y(n_149) );
INVx1_ASAP7_75t_L g155 ( .A(n_36), .Y(n_155) );
OR2x6_ASAP7_75t_L g111 ( .A(n_37), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_38), .B(n_143), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_39), .B(n_143), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_40), .B(n_170), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_41), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_42), .B(n_168), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_43), .B(n_143), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_44), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_45), .A2(n_151), .B(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_46), .A2(n_151), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_47), .B(n_168), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_48), .B(n_168), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_49), .B(n_143), .Y(n_207) );
INVx1_ASAP7_75t_L g137 ( .A(n_50), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_50), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_51), .B(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g216 ( .A(n_52), .B(n_128), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_53), .B(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_54), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_55), .B(n_170), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_56), .B(n_168), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_57), .A2(n_151), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_58), .B(n_143), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_59), .B(n_143), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_60), .A2(n_151), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g232 ( .A(n_61), .B(n_129), .Y(n_232) );
AO21x1_ASAP7_75t_L g493 ( .A1(n_62), .A2(n_151), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_63), .B(n_143), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_64), .B(n_168), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_65), .B(n_143), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_66), .B(n_168), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_67), .A2(n_91), .B1(n_151), .B2(n_153), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_68), .B(n_170), .Y(n_229) );
AND2x2_ASAP7_75t_L g506 ( .A(n_69), .B(n_129), .Y(n_506) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
INVx1_ASAP7_75t_L g148 ( .A(n_70), .Y(n_148) );
AND2x2_ASAP7_75t_L g547 ( .A(n_71), .B(n_174), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_72), .B(n_168), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_73), .A2(n_151), .B(n_220), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g116 ( .A1(n_74), .A2(n_117), .B1(n_746), .B2(n_747), .C(n_751), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_74), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_75), .A2(n_151), .B(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_76), .A2(n_151), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g242 ( .A(n_77), .B(n_129), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_78), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g114 ( .A(n_79), .Y(n_114) );
AND2x2_ASAP7_75t_L g458 ( .A(n_80), .B(n_174), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_81), .B(n_143), .Y(n_472) );
AND2x2_ASAP7_75t_L g197 ( .A(n_82), .B(n_185), .Y(n_197) );
AND2x2_ASAP7_75t_L g492 ( .A(n_83), .B(n_212), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_85), .B(n_168), .Y(n_471) );
AND2x2_ASAP7_75t_L g515 ( .A(n_86), .B(n_174), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_88), .B(n_170), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_89), .A2(n_151), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_90), .B(n_168), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_92), .A2(n_151), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_93), .B(n_170), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_94), .B(n_170), .Y(n_463) );
BUFx2_ASAP7_75t_L g231 ( .A(n_95), .Y(n_231) );
BUFx2_ASAP7_75t_L g106 ( .A(n_96), .Y(n_106) );
BUFx2_ASAP7_75t_SL g774 ( .A(n_96), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_97), .A2(n_151), .B(n_535), .Y(n_534) );
BUFx4f_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_107), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_SL g769 ( .A(n_104), .B(n_106), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_104), .A2(n_772), .B(n_775), .Y(n_771) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g762 ( .A(n_108), .Y(n_762) );
BUFx2_ASAP7_75t_L g765 ( .A(n_108), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x6_ASAP7_75t_SL g450 ( .A(n_109), .B(n_111), .Y(n_450) );
OR2x6_ASAP7_75t_SL g745 ( .A(n_109), .B(n_110), .Y(n_745) );
OR2x2_ASAP7_75t_L g755 ( .A(n_109), .B(n_111), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_447), .B1(n_451), .B2(n_743), .Y(n_117) );
INVx3_ASAP7_75t_L g748 ( .A(n_118), .Y(n_748) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_372), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_308), .C(n_355), .Y(n_119) );
NAND4xp25_ASAP7_75t_SL g120 ( .A(n_121), .B(n_243), .C(n_261), .D(n_287), .Y(n_120) );
OAI21xp33_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_201), .B(n_202), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_123), .B(n_186), .Y(n_122) );
INVx1_ASAP7_75t_L g423 ( .A(n_123), .Y(n_423) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_158), .Y(n_123) );
INVx2_ASAP7_75t_L g247 ( .A(n_124), .Y(n_247) );
AND2x2_ASAP7_75t_L g267 ( .A(n_124), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g369 ( .A(n_124), .B(n_188), .Y(n_369) );
AND2x2_ASAP7_75t_L g429 ( .A(n_124), .B(n_248), .Y(n_429) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_125), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g313 ( .A(n_126), .B(n_161), .Y(n_313) );
BUFx3_ASAP7_75t_L g323 ( .A(n_126), .Y(n_323) );
AND2x2_ASAP7_75t_L g386 ( .A(n_126), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
AND2x4_ASAP7_75t_L g200 ( .A(n_127), .B(n_132), .Y(n_200) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_128), .A2(n_133), .B(n_150), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_128), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_128), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_128), .A2(n_460), .B(n_461), .Y(n_459) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_128), .A2(n_481), .B(n_485), .Y(n_480) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_128), .A2(n_481), .B(n_485), .Y(n_551) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x4_ASAP7_75t_L g212 ( .A(n_130), .B(n_131), .Y(n_212) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g152 ( .A(n_137), .B(n_139), .Y(n_152) );
AND2x4_ASAP7_75t_L g170 ( .A(n_137), .B(n_147), .Y(n_170) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g151 ( .A(n_141), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
AND2x6_ASAP7_75t_L g168 ( .A(n_142), .B(n_145), .Y(n_168) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
AND2x4_ASAP7_75t_L g153 ( .A(n_152), .B(n_154), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g432 ( .A(n_159), .Y(n_432) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_175), .Y(n_159) );
AND2x2_ASAP7_75t_L g199 ( .A(n_160), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g387 ( .A(n_160), .Y(n_387) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g201 ( .A(n_161), .B(n_190), .Y(n_201) );
AND2x2_ASAP7_75t_L g264 ( .A(n_161), .B(n_175), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_161), .Y(n_269) );
AND2x2_ASAP7_75t_L g271 ( .A(n_161), .B(n_176), .Y(n_271) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_173), .Y(n_161) );
INVx4_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_172), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_168), .B(n_231), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_171), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_171), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_171), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_171), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_171), .A2(n_239), .B(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_171), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_171), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_171), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_171), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_171), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_171), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_171), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_171), .A2(n_544), .B(n_545), .Y(n_543) );
INVx3_ASAP7_75t_L g235 ( .A(n_174), .Y(n_235) );
INVx1_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
INVx2_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
AND2x4_ASAP7_75t_SL g284 ( .A(n_175), .B(n_190), .Y(n_284) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_175), .Y(n_316) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_176), .Y(n_198) );
AOI21x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_184), .Y(n_176) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_177), .A2(n_541), .B(n_547), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_183), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_226), .B(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_199), .Y(n_186) );
AND2x2_ASAP7_75t_L g350 ( .A(n_187), .B(n_295), .Y(n_350) );
INVx2_ASAP7_75t_SL g438 ( .A(n_187), .Y(n_438) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_189), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g358 ( .A(n_189), .B(n_271), .Y(n_358) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
AND2x4_ASAP7_75t_L g248 ( .A(n_190), .B(n_249), .Y(n_248) );
NOR2x1_ASAP7_75t_L g268 ( .A(n_190), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g341 ( .A(n_190), .Y(n_341) );
AND2x2_ASAP7_75t_L g360 ( .A(n_190), .B(n_299), .Y(n_360) );
AND2x2_ASAP7_75t_L g391 ( .A(n_190), .B(n_300), .Y(n_391) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_197), .Y(n_190) );
AND2x2_ASAP7_75t_L g330 ( .A(n_199), .B(n_284), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_199), .B(n_341), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_199), .A2(n_441), .B1(n_443), .B2(n_444), .Y(n_440) );
AND2x2_ASAP7_75t_L g443 ( .A(n_199), .B(n_250), .Y(n_443) );
INVx3_ASAP7_75t_L g296 ( .A(n_200), .Y(n_296) );
AND2x2_ASAP7_75t_L g299 ( .A(n_200), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g315 ( .A(n_201), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g324 ( .A(n_201), .Y(n_324) );
AND2x4_ASAP7_75t_SL g202 ( .A(n_203), .B(n_213), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_203), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g375 ( .A(n_203), .B(n_376), .Y(n_375) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_203), .B(n_337), .C(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g445 ( .A(n_203), .B(n_339), .Y(n_445) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g260 ( .A(n_205), .B(n_224), .Y(n_260) );
INVx1_ASAP7_75t_L g277 ( .A(n_205), .Y(n_277) );
INVx2_ASAP7_75t_L g290 ( .A(n_205), .Y(n_290) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_205), .Y(n_305) );
AND2x2_ASAP7_75t_L g319 ( .A(n_205), .B(n_292), .Y(n_319) );
AND2x2_ASAP7_75t_L g398 ( .A(n_205), .B(n_215), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_212), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_SL g466 ( .A(n_212), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_212), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_212), .A2(n_533), .B(n_534), .Y(n_532) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_213), .A2(n_262), .B1(n_265), .B2(n_272), .C(n_278), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_213), .A2(n_391), .B1(n_392), .B2(n_393), .C(n_394), .Y(n_390) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
INVx2_ASAP7_75t_L g332 ( .A(n_214), .Y(n_332) );
AND2x2_ASAP7_75t_L g392 ( .A(n_214), .B(n_276), .Y(n_392) );
AND2x2_ASAP7_75t_L g402 ( .A(n_214), .B(n_288), .Y(n_402) );
OR2x2_ASAP7_75t_L g442 ( .A(n_214), .B(n_326), .Y(n_442) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_SL g259 ( .A(n_215), .B(n_260), .Y(n_259) );
NAND2x1_ASAP7_75t_L g275 ( .A(n_215), .B(n_224), .Y(n_275) );
INVx4_ASAP7_75t_L g304 ( .A(n_215), .Y(n_304) );
OR2x2_ASAP7_75t_L g346 ( .A(n_215), .B(n_233), .Y(n_346) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g397 ( .A(n_223), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_233), .Y(n_223) );
INVx2_ASAP7_75t_SL g285 ( .A(n_224), .Y(n_285) );
NOR2x1_ASAP7_75t_SL g291 ( .A(n_224), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g306 ( .A(n_224), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g337 ( .A(n_224), .B(n_304), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_224), .B(n_290), .Y(n_344) );
BUFx2_ASAP7_75t_L g378 ( .A(n_224), .Y(n_378) );
AND2x2_ASAP7_75t_L g389 ( .A(n_224), .B(n_304), .Y(n_389) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_232), .Y(n_224) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
AND2x2_ASAP7_75t_L g276 ( .A(n_233), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g307 ( .A(n_233), .Y(n_307) );
AND2x2_ASAP7_75t_L g333 ( .A(n_233), .B(n_289), .Y(n_333) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_242), .Y(n_234) );
AO21x1_ASAP7_75t_SL g292 ( .A1(n_235), .A2(n_236), .B(n_242), .Y(n_292) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_235), .A2(n_500), .B(n_506), .Y(n_499) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_235), .A2(n_509), .B(n_515), .Y(n_508) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_235), .A2(n_509), .B(n_515), .Y(n_521) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_235), .A2(n_500), .B(n_506), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_241), .Y(n_236) );
OAI31xp33_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_248), .A3(n_250), .B(n_254), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g352 ( .A(n_246), .Y(n_352) );
NOR2xp67_ASAP7_75t_L g262 ( .A(n_247), .B(n_263), .Y(n_262) );
AOI322xp5_ASAP7_75t_L g342 ( .A1(n_247), .A2(n_336), .A3(n_343), .B1(n_347), .B2(n_348), .C1(n_350), .C2(n_351), .Y(n_342) );
AND2x2_ASAP7_75t_L g414 ( .A(n_247), .B(n_391), .Y(n_414) );
AOI221xp5_ASAP7_75t_SL g327 ( .A1(n_248), .A2(n_328), .B1(n_330), .B2(n_331), .C(n_334), .Y(n_327) );
INVx2_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_250), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_250), .B(n_343), .Y(n_446) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g321 ( .A(n_251), .B(n_296), .Y(n_321) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g300 ( .A(n_253), .B(n_269), .Y(n_300) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g371 ( .A(n_257), .Y(n_371) );
O2A1O1Ixp5_ASAP7_75t_L g362 ( .A1(n_258), .A2(n_363), .B(n_365), .C(n_367), .Y(n_362) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_259), .A2(n_395), .B1(n_396), .B2(n_399), .Y(n_394) );
OR2x2_ASAP7_75t_L g349 ( .A(n_260), .B(n_346), .Y(n_349) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_266), .B(n_270), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g282 ( .A(n_269), .Y(n_282) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_271), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g325 ( .A(n_275), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_275), .B(n_276), .Y(n_368) );
OR2x2_ASAP7_75t_L g370 ( .A(n_275), .B(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_275), .B(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g286 ( .A(n_277), .Y(n_286) );
NOR4xp25_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .C(n_285), .D(n_286), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g406 ( .A(n_280), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g434 ( .A(n_280), .B(n_283), .Y(n_434) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g364 ( .A(n_282), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_283), .B(n_312), .Y(n_399) );
AOI321xp33_ASAP7_75t_L g401 ( .A1(n_283), .A2(n_402), .A3(n_403), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_401) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_284), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_284), .B(n_323), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_285), .B(n_307), .Y(n_412) );
OR2x2_ASAP7_75t_L g439 ( .A(n_286), .B(n_323), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_293), .B(n_297), .Y(n_287) );
AND2x2_ASAP7_75t_L g328 ( .A(n_288), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g354 ( .A(n_290), .B(n_292), .Y(n_354) );
INVx2_ASAP7_75t_L g339 ( .A(n_291), .Y(n_339) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_294), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g395 ( .A(n_295), .B(n_347), .Y(n_395) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g353 ( .A(n_296), .B(n_354), .Y(n_353) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_296), .B(n_432), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_298), .B(n_301), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g382 ( .A(n_300), .Y(n_382) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NOR2xp67_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_304), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g329 ( .A(n_304), .Y(n_329) );
BUFx2_ASAP7_75t_L g411 ( .A(n_304), .Y(n_411) );
INVxp67_ASAP7_75t_L g419 ( .A(n_307), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_327), .C(n_342), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_317), .B(n_320), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g340 ( .A(n_313), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g393 ( .A(n_314), .Y(n_393) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g408 ( .A(n_316), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_317), .A2(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g326 ( .A(n_319), .Y(n_326) );
AND2x2_ASAP7_75t_L g388 ( .A(n_319), .B(n_389), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_325), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_321), .A2(n_368), .B1(n_369), .B2(n_370), .Y(n_367) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
OR2x2_ASAP7_75t_L g405 ( .A(n_326), .B(n_337), .Y(n_405) );
NOR4xp25_ASAP7_75t_L g437 ( .A(n_329), .B(n_378), .C(n_438), .D(n_439), .Y(n_437) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
OR2x2_ASAP7_75t_L g338 ( .A(n_332), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_332), .B(n_354), .Y(n_436) );
AOI21xp33_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_338), .B(n_340), .Y(n_334) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g425 ( .A(n_337), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g433 ( .A(n_339), .Y(n_433) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVxp67_ASAP7_75t_L g361 ( .A(n_344), .Y(n_361) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g377 ( .A(n_346), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g380 ( .A(n_352), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g426 ( .A(n_354), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B(n_361), .C(n_362), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g420 ( .A(n_363), .Y(n_420) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_400), .C(n_421), .Y(n_372) );
OAI211xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_379), .B(n_383), .C(n_390), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI21xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_423), .B(n_424), .C(n_427), .Y(n_422) );
BUFx2_ASAP7_75t_L g403 ( .A(n_387), .Y(n_403) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_413), .Y(n_400) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_410), .A2(n_416), .B1(n_417), .B2(n_420), .Y(n_415) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g421 ( .A(n_422), .B(n_430), .C(n_440), .D(n_446), .Y(n_421) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_434), .B2(n_435), .C(n_437), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx6p67_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_449), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_SL g750 ( .A(n_451), .Y(n_750) );
NOR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_630), .Y(n_451) );
AO211x2_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_475), .B(n_525), .C(n_598), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
AND3x2_ASAP7_75t_L g679 ( .A(n_455), .B(n_560), .C(n_576), .Y(n_679) );
AND2x4_ASAP7_75t_L g682 ( .A(n_455), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_456), .B(n_539), .Y(n_538) );
INVx4_ASAP7_75t_L g591 ( .A(n_456), .Y(n_591) );
AND2x2_ASAP7_75t_SL g676 ( .A(n_456), .B(n_585), .Y(n_676) );
AND2x2_ASAP7_75t_L g719 ( .A(n_456), .B(n_540), .Y(n_719) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g568 ( .A(n_457), .Y(n_568) );
AND2x2_ASAP7_75t_L g587 ( .A(n_457), .B(n_531), .Y(n_587) );
AND2x2_ASAP7_75t_L g605 ( .A(n_457), .B(n_540), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_457), .B(n_539), .Y(n_665) );
NOR2x1_ASAP7_75t_SL g692 ( .A(n_457), .B(n_465), .Y(n_692) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_465), .B(n_531), .Y(n_530) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_473), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_466), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_466), .A2(n_467), .B(n_473), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
AO21x1_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_507), .B(n_516), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_477), .A2(n_574), .B1(n_578), .B2(n_579), .Y(n_573) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
AND2x2_ASAP7_75t_L g634 ( .A(n_478), .B(n_522), .Y(n_634) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g567 ( .A(n_479), .B(n_550), .Y(n_567) );
AND2x2_ASAP7_75t_L g639 ( .A(n_479), .B(n_524), .Y(n_639) );
AND2x2_ASAP7_75t_L g658 ( .A(n_479), .B(n_624), .Y(n_658) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_480), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_486), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g618 ( .A(n_487), .B(n_519), .Y(n_618) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_499), .Y(n_487) );
AND2x2_ASAP7_75t_L g522 ( .A(n_488), .B(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g555 ( .A(n_488), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_488), .B(n_551), .Y(n_615) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g708 ( .A(n_489), .Y(n_708) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g550 ( .A(n_490), .Y(n_550) );
OAI21x1_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_493), .B(n_497), .Y(n_490) );
INVx1_ASAP7_75t_L g498 ( .A(n_492), .Y(n_498) );
INVx2_ASAP7_75t_L g556 ( .A(n_499), .Y(n_556) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_499), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_501), .B(n_505), .Y(n_500) );
INVx2_ASAP7_75t_L g552 ( .A(n_507), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_507), .B(n_684), .Y(n_710) );
AND2x2_ASAP7_75t_L g729 ( .A(n_507), .B(n_719), .Y(n_729) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_SL g597 ( .A(n_508), .B(n_556), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
AND2x2_ASAP7_75t_SL g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g596 ( .A(n_517), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_517), .B(n_566), .Y(n_601) );
INVx1_ASAP7_75t_SL g728 ( .A(n_517), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_518), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_L g554 ( .A(n_519), .Y(n_554) );
AND2x2_ASAP7_75t_L g740 ( .A(n_519), .B(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g616 ( .A(n_520), .B(n_523), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_520), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g670 ( .A(n_520), .B(n_524), .Y(n_670) );
AND2x2_ASAP7_75t_L g701 ( .A(n_520), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g566 ( .A(n_521), .B(n_524), .Y(n_566) );
INVxp67_ASAP7_75t_L g583 ( .A(n_521), .Y(n_583) );
BUFx3_ASAP7_75t_L g624 ( .A(n_521), .Y(n_624) );
AND2x2_ASAP7_75t_L g644 ( .A(n_522), .B(n_645), .Y(n_644) );
NAND2xp33_ASAP7_75t_L g657 ( .A(n_522), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_523), .B(n_550), .Y(n_613) );
AND2x2_ASAP7_75t_L g702 ( .A(n_523), .B(n_551), .Y(n_702) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g629 ( .A(n_524), .B(n_551), .Y(n_629) );
OR3x1_ASAP7_75t_L g525 ( .A(n_526), .B(n_573), .C(n_588), .Y(n_525) );
OAI321xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_538), .A3(n_548), .B1(n_553), .B2(n_557), .C(n_565), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_530), .Y(n_604) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_530), .Y(n_622) );
OR2x2_ASAP7_75t_L g626 ( .A(n_530), .B(n_538), .Y(n_626) );
BUFx3_ASAP7_75t_L g560 ( .A(n_531), .Y(n_560) );
AND2x2_ASAP7_75t_L g577 ( .A(n_531), .B(n_563), .Y(n_577) );
INVx1_ASAP7_75t_L g594 ( .A(n_531), .Y(n_594) );
INVx2_ASAP7_75t_L g610 ( .A(n_531), .Y(n_610) );
OR2x2_ASAP7_75t_L g649 ( .A(n_531), .B(n_539), .Y(n_649) );
INVx2_ASAP7_75t_L g637 ( .A(n_538), .Y(n_637) );
AND2x2_ASAP7_75t_L g561 ( .A(n_539), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g576 ( .A(n_539), .Y(n_576) );
AND2x4_ASAP7_75t_L g585 ( .A(n_539), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_539), .B(n_562), .Y(n_608) );
AND2x2_ASAP7_75t_L g715 ( .A(n_539), .B(n_610), .Y(n_715) );
INVx4_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
INVx1_ASAP7_75t_L g602 ( .A(n_548), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_552), .Y(n_548) );
AND2x2_ASAP7_75t_L g689 ( .A(n_549), .B(n_616), .Y(n_689) );
INVx1_ASAP7_75t_SL g706 ( .A(n_549), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_549), .B(n_682), .Y(n_735) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
OR2x2_ASAP7_75t_L g578 ( .A(n_550), .B(n_551), .Y(n_578) );
AND2x2_ASAP7_75t_L g671 ( .A(n_552), .B(n_567), .Y(n_671) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_556), .B(n_567), .Y(n_694) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_558), .A2(n_707), .B1(n_712), .B2(n_714), .Y(n_711) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g636 ( .A(n_559), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g731 ( .A(n_559), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g687 ( .A(n_560), .B(n_605), .Y(n_687) );
AND2x4_ASAP7_75t_L g641 ( .A(n_561), .B(n_587), .Y(n_641) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_563), .Y(n_739) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g572 ( .A(n_564), .Y(n_572) );
INVx1_ASAP7_75t_L g586 ( .A(n_564), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .C(n_568), .D(n_569), .Y(n_565) );
AND2x2_ASAP7_75t_L g723 ( .A(n_566), .B(n_708), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_566), .B(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_567), .B(n_643), .Y(n_642) );
OAI322xp33_ASAP7_75t_L g650 ( .A1(n_567), .A2(n_651), .A3(n_655), .B1(n_657), .B2(n_659), .C1(n_661), .C2(n_666), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_567), .B(n_616), .Y(n_666) );
INVx1_ASAP7_75t_L g734 ( .A(n_567), .Y(n_734) );
INVx2_ASAP7_75t_L g580 ( .A(n_568), .Y(n_580) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_571), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_572), .B(n_591), .Y(n_648) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_575), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g621 ( .A(n_576), .Y(n_621) );
AND2x2_ASAP7_75t_L g693 ( .A(n_576), .B(n_604), .Y(n_693) );
AOI31xp33_ASAP7_75t_L g579 ( .A1(n_577), .A2(n_580), .A3(n_581), .B(n_584), .Y(n_579) );
AND2x2_ASAP7_75t_L g590 ( .A(n_577), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g718 ( .A(n_577), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_577), .B(n_605), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_577), .Y(n_726) );
INVx1_ASAP7_75t_SL g684 ( .A(n_578), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_578), .B(n_706), .C(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g612 ( .A(n_583), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
AND2x2_ASAP7_75t_L g593 ( .A(n_585), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g654 ( .A(n_585), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g736 ( .A1(n_585), .A2(n_615), .A3(n_618), .B1(n_737), .B2(n_738), .C1(n_740), .C2(n_742), .Y(n_736) );
AND2x2_ASAP7_75t_L g742 ( .A(n_585), .B(n_591), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B(n_595), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_591), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g737 ( .A(n_591), .B(n_624), .Y(n_737) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g663 ( .A(n_594), .Y(n_663) );
AND2x2_ASAP7_75t_L g691 ( .A(n_594), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g738 ( .A(n_594), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g643 ( .A(n_597), .Y(n_643) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
O2A1O1Ixp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_603), .C(n_606), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g660 ( .A(n_605), .B(n_610), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_611), .B(n_617), .C(n_619), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_607), .A2(n_633), .B1(n_635), .B2(n_638), .C(n_640), .Y(n_632) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g652 ( .A(n_609), .Y(n_652) );
OR2x2_ASAP7_75t_L g672 ( .A(n_609), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g717 ( .A(n_612), .Y(n_717) );
INVx1_ASAP7_75t_L g741 ( .A(n_613), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g623 ( .A(n_615), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_615), .B(n_685), .Y(n_697) );
INVx1_ASAP7_75t_L g677 ( .A(n_616), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B1(n_625), .B2(n_627), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_SL g685 ( .A(n_624), .Y(n_685) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND4xp75_ASAP7_75t_L g630 ( .A(n_631), .B(n_667), .C(n_695), .D(n_720), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g631 ( .A(n_632), .B(n_650), .Y(n_631) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_639), .B(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_644), .B2(n_646), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_643), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g683 ( .A(n_649), .Y(n_683) );
OR2x2_ASAP7_75t_L g698 ( .A(n_649), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g713 ( .A(n_658), .Y(n_713) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_660), .A2(n_705), .B(n_707), .Y(n_704) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_680), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B1(n_675), .B2(n_677), .C(n_678), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OAI21xp33_ASAP7_75t_L g716 ( .A1(n_670), .A2(n_717), .B(n_718), .Y(n_716) );
INVx3_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .A3(n_685), .B1(n_686), .B2(n_688), .C1(n_690), .C2(n_694), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g703 ( .A(n_691), .Y(n_703) );
INVx1_ASAP7_75t_L g699 ( .A(n_692), .Y(n_699) );
AND2x2_ASAP7_75t_L g714 ( .A(n_692), .B(n_715), .Y(n_714) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_709), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_700), .B2(n_703), .C(n_704), .Y(n_696) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
OAI211xp5_ASAP7_75t_SL g709 ( .A1(n_703), .A2(n_710), .B(n_711), .C(n_716), .Y(n_709) );
INVx2_ASAP7_75t_SL g732 ( .A(n_719), .Y(n_732) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_730), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_726), .B2(n_727), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_733), .B(n_735), .C(n_736), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g749 ( .A(n_744), .Y(n_749) );
CKINVDCx11_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_763), .Y(n_757) );
CKINVDCx11_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx2_ASAP7_75t_L g775 ( .A(n_765), .Y(n_775) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
CKINVDCx11_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
CKINVDCx8_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
endmodule