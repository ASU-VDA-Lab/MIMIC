module fake_jpeg_31659_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_14),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_43),
.B1(n_32),
.B2(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_35),
.B1(n_33),
.B2(n_42),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_1),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_18),
.C(n_31),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_72),
.C(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_3),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_17),
.C(n_30),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_16),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_4),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_82),
.B(n_89),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_1),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_4),
.B(n_6),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_15),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_22),
.B1(n_7),
.B2(n_9),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_10),
.C(n_11),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_86),
.C(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_20),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_81),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_92),
.Y(n_104)
);

AOI321xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_96),
.A3(n_93),
.B1(n_85),
.B2(n_27),
.C(n_28),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_87),
.Y(n_106)
);


endmodule