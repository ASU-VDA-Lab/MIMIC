module fake_jpeg_30843_n_487 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_56),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_26),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_79),
.Y(n_122)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_90),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_8),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_16),
.Y(n_139)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_41),
.B1(n_31),
.B2(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_98),
.A2(n_114),
.B1(n_33),
.B2(n_47),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_30),
.B1(n_21),
.B2(n_45),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_30),
.B1(n_21),
.B2(n_45),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_119),
.B1(n_24),
.B2(n_47),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_26),
.B1(n_25),
.B2(n_16),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_41),
.B1(n_36),
.B2(n_43),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_126),
.B1(n_138),
.B2(n_150),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_36),
.B1(n_44),
.B2(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_25),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_144),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_75),
.A2(n_36),
.B1(n_44),
.B2(n_43),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_37),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_SL g142 ( 
.A(n_56),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_49),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_96),
.A2(n_44),
.B1(n_22),
.B2(n_49),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_98),
.A2(n_69),
.B1(n_70),
.B2(n_97),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_111),
.B(n_108),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_61),
.C(n_84),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_154),
.B(n_167),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_155),
.B(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_137),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_33),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_176),
.Y(n_206)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_159),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_165),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_68),
.B1(n_60),
.B2(n_52),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_164),
.A2(n_202),
.B1(n_120),
.B2(n_117),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_89),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_166),
.B(n_172),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_169),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_39),
.B(n_32),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_183),
.Y(n_217)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_171),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_121),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_24),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_31),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_181),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_37),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_182),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_101),
.B(n_54),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_37),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_50),
.C(n_88),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_91),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_200),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_105),
.A2(n_73),
.B1(n_63),
.B2(n_58),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_125),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_190),
.B(n_192),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_37),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_118),
.A2(n_63),
.B1(n_83),
.B2(n_37),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_112),
.B(n_143),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_8),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_195),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_126),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_127),
.A2(n_6),
.B(n_13),
.C(n_2),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_111),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_117),
.B(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_132),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_135),
.A2(n_9),
.B1(n_13),
.B2(n_2),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_238),
.B1(n_245),
.B2(n_164),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_213),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_159),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_179),
.A2(n_135),
.B(n_10),
.C(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_218),
.B(n_15),
.Y(n_274)
);

OAI22x1_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_145),
.B1(n_120),
.B2(n_132),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_153),
.B1(n_185),
.B2(n_131),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_108),
.B(n_107),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_185),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_153),
.B(n_176),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_240),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_200),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_174),
.B(n_112),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_239),
.C(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_177),
.A2(n_106),
.B(n_152),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_165),
.B(n_151),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_195),
.A2(n_145),
.B1(n_151),
.B2(n_131),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_247),
.A2(n_258),
.B1(n_276),
.B2(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_172),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_252),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_251),
.B1(n_253),
.B2(n_216),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_255),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_229),
.A2(n_175),
.B1(n_181),
.B2(n_154),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_156),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_161),
.B1(n_201),
.B2(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_262),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_206),
.A2(n_162),
.A3(n_167),
.B1(n_196),
.B2(n_168),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_155),
.B1(n_158),
.B2(n_199),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_279),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_206),
.B(n_200),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_270),
.Y(n_304)
);

BUFx8_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_194),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_165),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_273),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_236),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_188),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_275),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_215),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_208),
.A2(n_216),
.B1(n_238),
.B2(n_214),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_169),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_187),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_208),
.A2(n_198),
.B1(n_173),
.B2(n_178),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_216),
.A2(n_171),
.B1(n_166),
.B2(n_173),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_240),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_286),
.A2(n_293),
.B1(n_294),
.B2(n_305),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_204),
.B1(n_239),
.B2(n_207),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_208),
.B1(n_237),
.B2(n_217),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_250),
.A2(n_215),
.B(n_220),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_296),
.A2(n_299),
.B(n_284),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_261),
.A2(n_217),
.B1(n_204),
.B2(n_228),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_249),
.A2(n_251),
.B1(n_261),
.B2(n_217),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_247),
.A2(n_205),
.B1(n_230),
.B2(n_241),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_307),
.B1(n_311),
.B2(n_316),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_276),
.A2(n_205),
.B1(n_218),
.B2(n_236),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_228),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_309),
.C(n_310),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_228),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_254),
.B(n_236),
.C(n_240),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_265),
.B(n_224),
.C(n_231),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_318),
.C(n_272),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_262),
.A2(n_218),
.B1(n_203),
.B2(n_245),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_261),
.B(n_231),
.C(n_223),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_256),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_341),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_248),
.Y(n_322)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_339),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_R g325 ( 
.A(n_296),
.B(n_274),
.C(n_262),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_SL g372 ( 
.A(n_325),
.B(n_266),
.C(n_221),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_278),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_347),
.C(n_348),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_277),
.Y(n_327)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_328),
.B(n_333),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_286),
.A2(n_305),
.B1(n_294),
.B2(n_285),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_350),
.B1(n_311),
.B2(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_291),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_335),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_300),
.A2(n_246),
.B1(n_255),
.B2(n_252),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_336),
.A2(n_340),
.B1(n_343),
.B2(n_351),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_246),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_337),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_299),
.B(n_270),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_300),
.A2(n_263),
.B1(n_260),
.B2(n_271),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_317),
.B(n_304),
.C(n_313),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_342),
.A2(n_310),
.B(n_307),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_306),
.A2(n_282),
.B1(n_281),
.B2(n_280),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_314),
.B(n_269),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_344),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_267),
.Y(n_345)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_346),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_283),
.C(n_243),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_243),
.C(n_257),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_352),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_303),
.A2(n_222),
.B1(n_212),
.B2(n_259),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_292),
.B(n_213),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_357),
.B(n_329),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_318),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_360),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_326),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_361),
.A2(n_376),
.B1(n_379),
.B2(n_340),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_336),
.A2(n_320),
.B1(n_302),
.B2(n_301),
.Y(n_364)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_334),
.A2(n_320),
.B1(n_302),
.B2(n_295),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_298),
.C(n_221),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_375),
.C(n_347),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_372),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_266),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_373),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_288),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_342),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_288),
.C(n_210),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_330),
.A2(n_259),
.B1(n_244),
.B2(n_212),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_244),
.B1(n_212),
.B2(n_225),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_329),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_386),
.C(n_388),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_356),
.B(n_338),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_384),
.B(n_385),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_345),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_348),
.C(n_343),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_360),
.B(n_375),
.C(n_366),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_396),
.C(n_399),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_350),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_359),
.A2(n_325),
.B1(n_332),
.B2(n_346),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_394),
.A2(n_397),
.B1(n_376),
.B2(n_377),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_331),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_352),
.B1(n_349),
.B2(n_225),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_380),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_369),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_210),
.C(n_225),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_266),
.B1(n_189),
.B2(n_3),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_400),
.A2(n_365),
.B1(n_368),
.B2(n_362),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_189),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_354),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_189),
.C(n_1),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_374),
.C(n_373),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_363),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_405),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_408),
.A2(n_411),
.B1(n_403),
.B2(n_382),
.Y(n_434)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_394),
.A2(n_361),
.B1(n_369),
.B2(n_357),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_390),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_417),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_416),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_402),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_420),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_10),
.Y(n_438)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_391),
.A2(n_373),
.B(n_368),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_421),
.A2(n_381),
.B(n_362),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_382),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_404),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_423),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_434),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_409),
.A2(n_401),
.B1(n_388),
.B2(n_386),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_411),
.B1(n_410),
.B2(n_408),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_417),
.A2(n_396),
.B(n_383),
.Y(n_430)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

XOR2x1_ASAP7_75t_SL g431 ( 
.A(n_420),
.B(n_395),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_433),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_406),
.A2(n_389),
.B(n_399),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_432),
.A2(n_413),
.B(n_410),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_381),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_437),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_10),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_440),
.C(n_422),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_0),
.C(n_1),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_428),
.C(n_425),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_446),
.A2(n_449),
.B(n_450),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_434),
.C(n_437),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_439),
.B(n_414),
.Y(n_448)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_448),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_423),
.C(n_419),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_414),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_415),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_451),
.A2(n_454),
.B(n_433),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_407),
.B1(n_424),
.B2(n_421),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_453),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_424),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_459),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_453),
.Y(n_459)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_431),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_445),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_446),
.A2(n_427),
.B(n_440),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_463),
.A2(n_465),
.B(n_455),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_464),
.B(n_466),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_444),
.A2(n_438),
.B(n_9),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_4),
.C(n_12),
.Y(n_466)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_467),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_456),
.B(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_470),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_442),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_473),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_462),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_441),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_458),
.Y(n_478)
);

AO21x1_ASAP7_75t_L g481 ( 
.A1(n_478),
.A2(n_471),
.B(n_12),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_459),
.C(n_460),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_474),
.C(n_477),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_480),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_482),
.C(n_475),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_4),
.C(n_13),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_483),
.B(n_13),
.Y(n_485)
);

O2A1O1Ixp33_ASAP7_75t_SL g486 ( 
.A1(n_485),
.A2(n_4),
.B(n_15),
.C(n_451),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_4),
.B(n_15),
.Y(n_487)
);


endmodule