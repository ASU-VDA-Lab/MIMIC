module fake_jpeg_29794_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_49),
.Y(n_134)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_9),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_51),
.B(n_94),
.Y(n_148)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_63),
.Y(n_111)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_29),
.Y(n_147)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_19),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_25),
.B1(n_23),
.B2(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_8),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_97),
.A2(n_113),
.B1(n_122),
.B2(n_123),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_35),
.B1(n_41),
.B2(n_30),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_99),
.A2(n_103),
.B1(n_105),
.B2(n_62),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_41),
.B1(n_30),
.B2(n_44),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_41),
.B1(n_30),
.B2(n_44),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_24),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_22),
.B1(n_44),
.B2(n_30),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_36),
.B1(n_40),
.B2(n_45),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_56),
.A2(n_22),
.B1(n_44),
.B2(n_42),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_57),
.A2(n_30),
.B1(n_22),
.B2(n_32),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_55),
.B(n_45),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_58),
.B(n_40),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_147),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_59),
.B(n_29),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_42),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_156),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_52),
.A2(n_24),
.B(n_32),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_37),
.B(n_39),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_70),
.B(n_26),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_161),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_95),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_160),
.B(n_168),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_73),
.B1(n_91),
.B2(n_71),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_162),
.A2(n_184),
.B1(n_207),
.B2(n_135),
.Y(n_232)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_93),
.B1(n_77),
.B2(n_75),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_166),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_248)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_49),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_192),
.B1(n_199),
.B2(n_211),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_111),
.A2(n_85),
.B1(n_83),
.B2(n_76),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_172),
.A2(n_176),
.B1(n_178),
.B2(n_186),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_173),
.A2(n_113),
.A3(n_145),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_26),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_174),
.B(n_182),
.Y(n_253)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_111),
.A2(n_72),
.B1(n_37),
.B2(n_39),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_114),
.A2(n_37),
.B1(n_39),
.B2(n_10),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_102),
.A2(n_37),
.B1(n_39),
.B2(n_8),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_99),
.A2(n_39),
.B(n_37),
.C(n_2),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_132),
.A2(n_37),
.B1(n_39),
.B2(n_8),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_98),
.B(n_101),
.C(n_104),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_187),
.B(n_206),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_126),
.A2(n_7),
.B(n_15),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_214),
.Y(n_217)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_119),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_190),
.Y(n_264)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_191),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_119),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_192)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_128),
.B(n_17),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_200),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_134),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_198)
);

AOI22x1_ASAP7_75t_L g262 ( 
.A1(n_198),
.A2(n_209),
.B1(n_207),
.B2(n_184),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_17),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_203),
.Y(n_235)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_11),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_116),
.A2(n_12),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_103),
.A2(n_12),
.B(n_3),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_209),
.B(n_210),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_0),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_152),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_215),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_153),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_216),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_152),
.B1(n_135),
.B2(n_146),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_231),
.B1(n_239),
.B2(n_259),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_158),
.A2(n_105),
.B1(n_124),
.B2(n_133),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_262),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_171),
.B(n_124),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_234),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_196),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_166),
.A2(n_133),
.B1(n_115),
.B2(n_145),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_255),
.B1(n_182),
.B2(n_198),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_196),
.A2(n_146),
.B1(n_157),
.B2(n_153),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_259),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_0),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_212),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_193),
.B(n_3),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_206),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_184),
.A2(n_5),
.B1(n_158),
.B2(n_168),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_208),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_261),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_199),
.A2(n_5),
.B1(n_168),
.B2(n_200),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_169),
.A2(n_214),
.B(n_160),
.C(n_159),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_268),
.B(n_276),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_160),
.B1(n_174),
.B2(n_187),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_174),
.B1(n_163),
.B2(n_164),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_161),
.B1(n_210),
.B2(n_194),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_161),
.C(n_215),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_274),
.C(n_237),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_234),
.C(n_257),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_280),
.B1(n_236),
.B2(n_237),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_189),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_210),
.B1(n_181),
.B2(n_213),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

BUFx8_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_278),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_231),
.A2(n_167),
.B1(n_175),
.B2(n_181),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_279),
.A2(n_286),
.B1(n_295),
.B2(n_298),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_219),
.A2(n_216),
.B1(n_191),
.B2(n_165),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_203),
.B1(n_201),
.B2(n_180),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_292),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_288),
.B(n_294),
.Y(n_338)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_289),
.A2(n_299),
.B1(n_305),
.B2(n_308),
.Y(n_349)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_290),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_225),
.A2(n_197),
.B1(n_212),
.B2(n_183),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_179),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_212),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_300),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_235),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_253),
.A2(n_177),
.B1(n_185),
.B2(n_202),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_219),
.A2(n_202),
.B1(n_242),
.B2(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_297),
.A2(n_260),
.B1(n_224),
.B2(n_248),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_253),
.A2(n_202),
.B1(n_262),
.B2(n_265),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_217),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_229),
.B(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_303),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_235),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_302),
.B(n_304),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_217),
.B(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_222),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_307),
.Y(n_335)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_223),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_221),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_274),
.B(n_227),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_314),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_285),
.A2(n_262),
.B1(n_263),
.B2(n_248),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_312),
.A2(n_316),
.B1(n_318),
.B2(n_320),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_227),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_319),
.C(n_325),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_252),
.C(n_246),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_261),
.B1(n_256),
.B2(n_243),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_252),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_244),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_328),
.B(n_332),
.C(n_333),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_297),
.A2(n_243),
.B1(n_244),
.B2(n_238),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_331),
.A2(n_334),
.B1(n_279),
.B2(n_286),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_273),
.B(n_246),
.C(n_224),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_238),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_296),
.A2(n_250),
.B1(n_251),
.B2(n_247),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_292),
.B(n_293),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_337),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_250),
.C(n_247),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_241),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_344),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_282),
.A2(n_258),
.B(n_228),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_346),
.B(n_267),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_251),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_282),
.B(n_228),
.C(n_221),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_345),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_282),
.A2(n_269),
.B(n_285),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_271),
.B(n_287),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_341),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_339),
.Y(n_353)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_L g354 ( 
.A1(n_329),
.A2(n_268),
.B(n_283),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_354),
.Y(n_407)
);

AOI21x1_ASAP7_75t_SL g355 ( 
.A1(n_345),
.A2(n_283),
.B(n_277),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_355),
.A2(n_337),
.B(n_346),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_313),
.A2(n_284),
.B(n_295),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_356),
.A2(n_372),
.B(n_373),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_322),
.B(n_338),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_358),
.A2(n_375),
.B1(n_379),
.B2(n_381),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_336),
.B(n_270),
.Y(n_361)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_330),
.B(n_266),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_363),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_342),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_364),
.Y(n_397)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_366),
.A2(n_376),
.B1(n_349),
.B2(n_305),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_324),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_367),
.Y(n_398)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_368),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_284),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_374),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_313),
.A2(n_304),
.B(n_290),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_326),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_323),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_326),
.B(n_307),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_377),
.B(n_382),
.Y(n_395)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_305),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_334),
.B1(n_331),
.B2(n_323),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_384),
.A2(n_392),
.B1(n_404),
.B2(n_406),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_315),
.C(n_311),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_399),
.C(n_403),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_362),
.A2(n_317),
.B1(n_348),
.B2(n_343),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_390),
.A2(n_396),
.B1(n_402),
.B2(n_368),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_370),
.A2(n_347),
.B1(n_317),
.B2(n_348),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_332),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_362),
.A2(n_319),
.B1(n_325),
.B2(n_328),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_314),
.C(n_333),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_372),
.A2(n_340),
.B1(n_327),
.B2(n_289),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_355),
.A2(n_272),
.B1(n_299),
.B2(n_278),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_308),
.C(n_278),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_369),
.C(n_378),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_353),
.A2(n_278),
.B1(n_308),
.B2(n_374),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_410),
.A2(n_366),
.B1(n_376),
.B2(n_350),
.Y(n_424)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_357),
.C(n_378),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_395),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_380),
.CI(n_359),
.CON(n_416),
.SN(n_416)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_416),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_375),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_420),
.Y(n_437)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_428),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_423),
.C(n_426),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_369),
.C(n_357),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_424),
.A2(n_429),
.B1(n_390),
.B2(n_388),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_361),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_433),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_365),
.C(n_382),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_352),
.B1(n_360),
.B2(n_379),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_427),
.A2(n_405),
.B1(n_410),
.B2(n_407),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_383),
.A2(n_356),
.B(n_373),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_392),
.A2(n_360),
.B1(n_381),
.B2(n_367),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_430),
.A2(n_384),
.B1(n_404),
.B2(n_406),
.Y(n_436)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_387),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_432),
.Y(n_450)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_367),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_391),
.B(n_308),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_434),
.B(n_391),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_436),
.B(n_413),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_447),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_451),
.Y(n_462)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_446),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_385),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_416),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_393),
.C(n_383),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_452),
.C(n_433),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_417),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_426),
.C(n_422),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_455),
.B(n_466),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_412),
.C(n_423),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_463),
.C(n_435),
.Y(n_469)
);

OAI221xp5_ASAP7_75t_L g457 ( 
.A1(n_444),
.A2(n_415),
.B1(n_428),
.B2(n_432),
.C(n_421),
.Y(n_457)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_461),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_459),
.A2(n_445),
.B1(n_442),
.B2(n_444),
.Y(n_471)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_430),
.Y(n_463)
);

AOI21xp33_ASAP7_75t_L g464 ( 
.A1(n_440),
.A2(n_414),
.B(n_420),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_464),
.A2(n_388),
.B(n_450),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_468),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_449),
.B(n_429),
.Y(n_466)
);

BUFx24_ASAP7_75t_SL g467 ( 
.A(n_448),
.Y(n_467)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_467),
.Y(n_475)
);

NOR3xp33_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_397),
.C(n_411),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_470),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_439),
.C(n_447),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_478),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_456),
.A2(n_439),
.B(n_442),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_472),
.B(n_441),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_462),
.A2(n_388),
.B(n_397),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_479),
.A2(n_453),
.B(n_400),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_398),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_480),
.B(n_398),
.Y(n_481)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_483),
.B(n_487),
.Y(n_492)
);

MAJx2_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_462),
.C(n_461),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_485),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_473),
.A2(n_436),
.B1(n_413),
.B2(n_438),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_437),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_488),
.B(n_476),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_486),
.A2(n_474),
.B1(n_479),
.B2(n_471),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_491),
.Y(n_496)
);

INVx11_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_493),
.Y(n_494)
);

OAI321xp33_ASAP7_75t_L g495 ( 
.A1(n_492),
.A2(n_485),
.A3(n_453),
.B1(n_424),
.B2(n_396),
.C(n_400),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_SL g497 ( 
.A1(n_495),
.A2(n_490),
.B(n_489),
.C(n_491),
.Y(n_497)
);

A2O1A1O1Ixp25_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_498),
.B(n_489),
.C(n_469),
.D(n_494),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_496),
.B(n_484),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_499),
.A2(n_475),
.B(n_460),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_394),
.B(n_460),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_501),
.A2(n_394),
.B1(n_393),
.B2(n_463),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_416),
.Y(n_503)
);


endmodule