module fake_netlist_5_1748_n_1878 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1878);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1878;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_48),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_57),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_68),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_45),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_15),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_128),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_7),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_101),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_73),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_69),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_77),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_82),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_43),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_32),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_21),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_24),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_75),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_90),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_8),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_60),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_107),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_16),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_164),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_67),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_51),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_23),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_99),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_28),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_85),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_155),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_58),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_25),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_46),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_39),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_52),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_98),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_48),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_22),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_29),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_153),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_123),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_59),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_53),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_30),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_67),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_93),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_27),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_24),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_53),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_162),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_122),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_43),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_28),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_83),
.Y(n_273)
);

BUFx8_ASAP7_75t_SL g274 ( 
.A(n_140),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_37),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_163),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_94),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_64),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_115),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_17),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_158),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_26),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_38),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_55),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_64),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_110),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_124),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_76),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_21),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_20),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_36),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_31),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_33),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_63),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_32),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_15),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_175),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_60),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_6),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_97),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_165),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_136),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_95),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_154),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_8),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_10),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_61),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_152),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_169),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_40),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_70),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_113),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_168),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_66),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_105),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_86),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_54),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_74),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_61),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_19),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_79),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_104),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_71),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_30),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_5),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_42),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_37),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_33),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_147),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_80),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_14),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_171),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_112),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_14),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_20),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_2),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_116),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_130),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_142),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_29),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_50),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_127),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_50),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_166),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_146),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_159),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_247),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_180),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_274),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_247),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_219),
.B(n_0),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_216),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_223),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_247),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_247),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_200),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_234),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_247),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_201),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_242),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_289),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_249),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_230),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_254),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_247),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_252),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_219),
.B(n_1),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_255),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_252),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_262),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_279),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_200),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_252),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_281),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_290),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_304),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_305),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_176),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_218),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_222),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_226),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_179),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_189),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_252),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_227),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_176),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_231),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_185),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_188),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_252),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_177),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_177),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_252),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_252),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_259),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_236),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_237),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_252),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_243),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_219),
.B(n_1),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_259),
.B(n_3),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_179),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_303),
.B(n_4),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_238),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_181),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_240),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_213),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_246),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_248),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_181),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_182),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_243),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_182),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_250),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_187),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_243),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_225),
.B(n_4),
.Y(n_426)
);

INVxp33_ASAP7_75t_SL g427 ( 
.A(n_184),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_243),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_257),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_243),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_245),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_193),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_187),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_258),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_260),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_261),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_267),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_271),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_278),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_377),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_362),
.B(n_213),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_357),
.B(n_225),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_357),
.B(n_179),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_245),
.Y(n_446)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_375),
.B(n_320),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_320),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_380),
.B(n_245),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_428),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_358),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_377),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_343),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_343),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_353),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_407),
.B(n_183),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_352),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_352),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_356),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_359),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_356),
.B(n_178),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_360),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_380),
.B(n_245),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_361),
.B(n_245),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_427),
.B(n_268),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_361),
.B(n_186),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_363),
.B(n_192),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_365),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_363),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_364),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_396),
.A2(n_333),
.B1(n_269),
.B2(n_264),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_364),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_366),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_366),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_373),
.B(n_322),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_373),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_381),
.B(n_192),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_389),
.B(n_277),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

INVx6_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_370),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_406),
.B(n_194),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_407),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_378),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_404),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_455),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_440),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_470),
.Y(n_523)
);

AND3x4_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_412),
.C(n_322),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

NOR2x1p5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_355),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_478),
.Y(n_527)
);

AOI21x1_ASAP7_75t_L g528 ( 
.A1(n_457),
.A2(n_412),
.B(n_191),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_473),
.B(n_390),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_460),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_460),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_440),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_462),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_462),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_473),
.B(n_379),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_462),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_481),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_446),
.B(n_382),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_491),
.B(n_383),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_446),
.B(n_384),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_453),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_303),
.Y(n_545)
);

BUFx4f_ASAP7_75t_L g546 ( 
.A(n_515),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_481),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_511),
.B(n_198),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_455),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_451),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_483),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_442),
.B(n_446),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_445),
.B(n_386),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_447),
.B(n_385),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_442),
.B(n_411),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_L g558 ( 
.A1(n_502),
.A2(n_396),
.B1(n_233),
.B2(n_266),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_483),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_455),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_486),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_451),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_455),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_508),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_405),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_502),
.B(n_413),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_509),
.B(n_415),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_460),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_444),
.B(n_183),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_509),
.B(n_417),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_484),
.B(n_418),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_487),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_461),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_508),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_466),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_480),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_464),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_488),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_464),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_447),
.B(n_423),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_488),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_511),
.B(n_429),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_461),
.B(n_434),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_515),
.B(n_435),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_492),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_515),
.B(n_436),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_477),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_515),
.B(n_437),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_477),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_477),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_480),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_466),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_492),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_460),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_450),
.B(n_190),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_475),
.B(n_438),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_493),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_510),
.B(n_439),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_515),
.B(n_372),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_494),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_494),
.Y(n_613)
);

AO22x2_ASAP7_75t_L g614 ( 
.A1(n_444),
.A2(n_294),
.B1(n_272),
.B2(n_244),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_450),
.B(n_204),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_482),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_495),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_466),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_460),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_495),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_485),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_496),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_460),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_496),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_466),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_466),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

BUFx4f_ASAP7_75t_L g630 ( 
.A(n_515),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_500),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_485),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_444),
.B(n_183),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_447),
.A2(n_272),
.B1(n_294),
.B2(n_263),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_480),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_447),
.A2(n_209),
.B1(n_275),
.B2(n_315),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_466),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_376),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_450),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_475),
.B(n_506),
.C(n_489),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_510),
.B(n_394),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_445),
.B(n_399),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_501),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_501),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_466),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_501),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_444),
.A2(n_297),
.B1(n_228),
.B2(n_220),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_516),
.B(n_400),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_516),
.B(n_414),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_441),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_471),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_472),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_472),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_472),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_471),
.B(n_313),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_516),
.B(n_419),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_441),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_489),
.B(n_215),
.C(n_207),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_443),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_443),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_463),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_221),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_469),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_484),
.B(n_403),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_448),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_448),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_452),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_452),
.Y(n_668)
);

BUFx8_ASAP7_75t_SL g669 ( 
.A(n_490),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_651),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_554),
.B(n_515),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_587),
.B(n_556),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_650),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_651),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_554),
.B(n_640),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_640),
.B(n_516),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_539),
.B(n_457),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_664),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_664),
.B(n_504),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_543),
.B(n_506),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_589),
.B(n_476),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_576),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_651),
.B(n_444),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_468),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_636),
.B(n_505),
.Y(n_685)
);

INVxp33_ASAP7_75t_SL g686 ( 
.A(n_638),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_634),
.A2(n_497),
.B1(n_371),
.B2(n_433),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_578),
.B(n_498),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_546),
.B(n_504),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_650),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_657),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_606),
.B(n_217),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_652),
.B(n_471),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_606),
.A2(n_497),
.B1(n_424),
.B2(n_422),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_653),
.A2(n_474),
.B1(n_468),
.B2(n_484),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_653),
.A2(n_513),
.B(n_512),
.C(n_514),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_546),
.B(n_504),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_654),
.B(n_518),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_568),
.B(n_514),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_576),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_657),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_568),
.B(n_490),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_666),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_639),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_557),
.B(n_512),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_569),
.B(n_479),
.C(n_498),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_557),
.B(n_512),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_654),
.B(n_468),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_518),
.B(n_468),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_614),
.A2(n_468),
.B1(n_474),
.B2(n_456),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_573),
.B(n_217),
.Y(n_711)
);

AOI22x1_ASAP7_75t_L g712 ( 
.A1(n_614),
.A2(n_474),
.B1(n_513),
.B2(n_459),
.Y(n_712)
);

BUFx5_ASAP7_75t_L g713 ( 
.A(n_531),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_666),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_609),
.A2(n_497),
.B1(n_420),
.B2(n_474),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_519),
.B(n_474),
.Y(n_716)
);

AO221x1_ASAP7_75t_L g717 ( 
.A1(n_614),
.A2(n_558),
.B1(n_195),
.B2(n_300),
.C(n_197),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_571),
.B(n_513),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_639),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_639),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_L g721 ( 
.A1(n_655),
.A2(n_479),
.B1(n_497),
.B2(n_354),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_546),
.B(n_469),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_521),
.B(n_469),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_521),
.B(n_469),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_590),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_524),
.A2(n_212),
.B1(n_214),
.B2(n_235),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_550),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_639),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_550),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_630),
.B(n_469),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_610),
.B(n_497),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_630),
.B(n_549),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_549),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_614),
.A2(n_615),
.B1(n_603),
.B2(n_562),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_575),
.B(n_497),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_552),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_523),
.B(n_469),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_630),
.B(n_499),
.Y(n_738)
);

AND2x4_ASAP7_75t_SL g739 ( 
.A(n_619),
.B(n_367),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_552),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_562),
.B(n_499),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_563),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_529),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_563),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_535),
.B(n_338),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_540),
.B(n_349),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_564),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_590),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_581),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_564),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_668),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_668),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_523),
.B(n_499),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_540),
.B(n_194),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_598),
.B(n_635),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_525),
.B(n_499),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_525),
.B(n_499),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_540),
.B(n_499),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_527),
.B(n_499),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_659),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_603),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_540),
.B(n_503),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_603),
.B(n_503),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_603),
.B(n_503),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_615),
.A2(n_449),
.B1(n_456),
.B2(n_459),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_615),
.B(n_527),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_591),
.B(n_196),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_615),
.B(n_183),
.Y(n_768)
);

HB1xp67_ASAP7_75t_SL g769 ( 
.A(n_641),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_593),
.B(n_196),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_658),
.A2(n_293),
.B(n_299),
.C(n_286),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_538),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_538),
.B(n_503),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_L g774 ( 
.A(n_648),
.B(n_454),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_547),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_545),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_545),
.Y(n_777)
);

AND2x6_ASAP7_75t_L g778 ( 
.A(n_531),
.B(n_183),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_649),
.B(n_656),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_547),
.B(n_503),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_553),
.B(n_503),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_573),
.B(n_217),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_545),
.A2(n_368),
.B1(n_369),
.B2(n_276),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_531),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_553),
.A2(n_265),
.B(n_324),
.C(n_325),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_555),
.B(n_287),
.C(n_280),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_559),
.B(n_561),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_659),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_660),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_559),
.B(n_503),
.Y(n_790)
);

INVx8_ASAP7_75t_L g791 ( 
.A(n_545),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_545),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_662),
.B(n_229),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_561),
.B(n_449),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_660),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_570),
.B(n_449),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_570),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_574),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_574),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_577),
.B(n_585),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_577),
.B(n_449),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_585),
.B(n_449),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_662),
.B(n_232),
.Y(n_803)
);

AND2x4_ASAP7_75t_SL g804 ( 
.A(n_619),
.B(n_224),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_658),
.A2(n_284),
.B(n_330),
.C(n_331),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_588),
.B(n_592),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_595),
.B(n_454),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_588),
.B(n_456),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_592),
.B(n_197),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_601),
.B(n_199),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_601),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_604),
.B(n_456),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_604),
.B(n_456),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_608),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_662),
.A2(n_626),
.B1(n_631),
.B2(n_625),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_608),
.B(n_197),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_619),
.B(n_459),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_612),
.B(n_459),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_612),
.B(n_459),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_613),
.B(n_197),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_613),
.B(n_458),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_617),
.B(n_458),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_665),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_665),
.Y(n_824)
);

AO22x2_ASAP7_75t_L g825 ( 
.A1(n_524),
.A2(n_348),
.B1(n_346),
.B2(n_341),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_667),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_617),
.B(n_621),
.Y(n_827)
);

INVxp33_ASAP7_75t_SL g828 ( 
.A(n_548),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_621),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_620),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_623),
.B(n_507),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_667),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_623),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_625),
.B(n_507),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_626),
.B(n_197),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_642),
.B(n_295),
.C(n_296),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_631),
.B(n_239),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_663),
.B(n_241),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_566),
.B(n_300),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_644),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_680),
.B(n_619),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_755),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_675),
.A2(n_662),
.B(n_644),
.C(n_583),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_672),
.A2(n_662),
.B1(n_524),
.B2(n_526),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_749),
.Y(n_845)
);

AO21x1_ASAP7_75t_L g846 ( 
.A1(n_672),
.A2(n_528),
.B(n_256),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_677),
.B(n_517),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_676),
.A2(n_526),
.B1(n_647),
.B2(n_530),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_718),
.B(n_517),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_683),
.A2(n_572),
.B(n_530),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_679),
.B(n_544),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_704),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_671),
.B(n_566),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_735),
.B(n_517),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_684),
.A2(n_602),
.B(n_572),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_704),
.B(n_620),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_686),
.B(n_580),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_733),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_772),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_184),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_689),
.B(n_620),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_743),
.B(n_566),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_693),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_694),
.B(n_203),
.C(n_202),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_705),
.B(n_536),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_L g866 ( 
.A1(n_745),
.A2(n_292),
.B(n_291),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_736),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_681),
.B(n_580),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_702),
.B(n_206),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_602),
.B(n_624),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_722),
.A2(n_624),
.B(n_618),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_707),
.B(n_536),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_758),
.A2(n_270),
.B(n_251),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_760),
.B(n_536),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_772),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_708),
.A2(n_584),
.B(n_583),
.Y(n_877)
);

AOI21x1_ASAP7_75t_L g878 ( 
.A1(n_730),
.A2(n_594),
.B(n_586),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_742),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_678),
.A2(n_583),
.B(n_584),
.C(n_646),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_709),
.A2(n_584),
.B(n_586),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_730),
.A2(n_738),
.B(n_732),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_689),
.A2(n_594),
.B(n_646),
.C(n_596),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_769),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_775),
.Y(n_885)
);

AO21x1_ASAP7_75t_L g886 ( 
.A1(n_815),
.A2(n_282),
.B(n_273),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_L g887 ( 
.A1(n_745),
.A2(n_211),
.B(n_206),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_697),
.A2(n_596),
.B(n_597),
.C(n_643),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_788),
.B(n_536),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_775),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_738),
.A2(n_624),
.B(n_618),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_732),
.A2(n_627),
.B(n_618),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_693),
.B(n_542),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_789),
.B(n_542),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_693),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_797),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_734),
.A2(n_542),
.B1(n_565),
.B2(n_328),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_725),
.B(n_211),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_716),
.A2(n_607),
.B(n_597),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_695),
.A2(n_565),
.B1(n_542),
.B2(n_327),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_784),
.A2(n_830),
.B(n_764),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_795),
.B(n_565),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_784),
.A2(n_627),
.B(n_618),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_681),
.B(n_580),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_823),
.B(n_565),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_697),
.A2(n_307),
.B(n_288),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_688),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_748),
.B(n_253),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_743),
.A2(n_319),
.B(n_285),
.C(n_306),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_830),
.A2(n_627),
.B(n_628),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_746),
.B(n_580),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_744),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_763),
.A2(n_764),
.B(n_729),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_746),
.A2(n_318),
.B(n_317),
.C(n_316),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_682),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_719),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_727),
.B(n_692),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_766),
.A2(n_627),
.B(n_628),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_719),
.B(n_566),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_824),
.B(n_637),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_797),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_747),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_826),
.B(n_637),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_798),
.Y(n_924)
);

NOR2x1_ASAP7_75t_L g925 ( 
.A(n_779),
.B(n_637),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_766),
.A2(n_628),
.B(n_551),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_700),
.B(n_720),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_685),
.A2(n_607),
.B(n_611),
.C(n_643),
.Y(n_928)
);

AOI21x1_ASAP7_75t_L g929 ( 
.A1(n_758),
.A2(n_611),
.B(n_616),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_791),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_741),
.A2(n_616),
.B(n_622),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_750),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_817),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_771),
.A2(n_805),
.B(n_698),
.C(n_800),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_804),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_832),
.B(n_637),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_706),
.B(n_622),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_SL g938 ( 
.A1(n_787),
.A2(n_548),
.B(n_314),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_798),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_828),
.B(n_645),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_799),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_833),
.B(n_645),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_806),
.B(n_645),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_728),
.B(n_566),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_741),
.A2(n_628),
.B(n_550),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_799),
.B(n_645),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_811),
.B(n_814),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_811),
.B(n_629),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_761),
.B(n_566),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_814),
.B(n_629),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_829),
.B(n_632),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_762),
.A2(n_560),
.B(n_551),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_754),
.B(n_632),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_791),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_673),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_774),
.B(n_520),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_670),
.B(n_520),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_674),
.B(n_522),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_673),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_762),
.A2(n_560),
.B(n_550),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_690),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_810),
.B(n_522),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_791),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_794),
.A2(n_560),
.B(n_550),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_690),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_796),
.A2(n_551),
.B(n_560),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_810),
.B(n_532),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_691),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_754),
.B(n_551),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_787),
.A2(n_567),
.B(n_533),
.C(n_534),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_715),
.B(n_687),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_804),
.B(n_253),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_767),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_713),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_800),
.B(n_827),
.Y(n_975)
);

NOR2x2_ASAP7_75t_L g976 ( 
.A(n_731),
.B(n_669),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_801),
.A2(n_551),
.B(n_560),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_827),
.B(n_533),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_802),
.A2(n_599),
.B(n_661),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_808),
.A2(n_599),
.B(n_661),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_812),
.A2(n_599),
.B(n_661),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_691),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_813),
.A2(n_819),
.B(n_818),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_701),
.B(n_537),
.Y(n_984)
);

BUFx4f_ASAP7_75t_L g985 ( 
.A(n_731),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_739),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_765),
.A2(n_599),
.B(n_661),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_701),
.B(n_703),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_703),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_773),
.A2(n_567),
.B(n_579),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_771),
.A2(n_350),
.B(n_308),
.C(n_351),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_714),
.Y(n_992)
);

OR2x6_ASAP7_75t_SL g993 ( 
.A(n_739),
.B(n_310),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_767),
.A2(n_573),
.B1(n_633),
.B2(n_203),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_714),
.B(n_579),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_751),
.B(n_600),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_751),
.B(n_600),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_752),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_723),
.A2(n_582),
.B(n_633),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_724),
.A2(n_661),
.B(n_605),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_752),
.B(n_600),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_717),
.A2(n_633),
.B1(n_573),
.B2(n_217),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_737),
.A2(n_605),
.B(n_600),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_753),
.A2(n_605),
.B(n_600),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_776),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_712),
.A2(n_633),
.B1(n_573),
.B2(n_217),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_773),
.A2(n_582),
.B(n_573),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_756),
.A2(n_605),
.B(n_600),
.Y(n_1008)
);

AOI22x1_ASAP7_75t_L g1009 ( 
.A1(n_793),
.A2(n_582),
.B1(n_202),
.B2(n_326),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_840),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_770),
.B(n_821),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_831),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_757),
.A2(n_605),
.B(n_300),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_759),
.A2(n_605),
.B(n_300),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_834),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_780),
.A2(n_300),
.B(n_633),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_726),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_781),
.A2(n_790),
.B(n_696),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_777),
.A2(n_326),
.B1(n_208),
.B2(n_210),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_726),
.A2(n_633),
.B1(n_573),
.B2(n_217),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_770),
.B(n_205),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_822),
.B(n_205),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_792),
.B(n_793),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_783),
.B(n_224),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_805),
.A2(n_329),
.B(n_345),
.C(n_340),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_793),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_838),
.A2(n_208),
.B(n_347),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_710),
.A2(n_210),
.B(n_347),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_803),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_711),
.A2(n_337),
.B(n_321),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_973),
.B(n_721),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_841),
.B(n_807),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_841),
.A2(n_731),
.B1(n_803),
.B2(n_837),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_974),
.A2(n_803),
.B(n_782),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_930),
.B(n_726),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_971),
.A2(n_836),
.B(n_786),
.C(n_785),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_859),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_971),
.A2(n_835),
.B(n_809),
.C(n_820),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_845),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_930),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_R g1041 ( 
.A(n_884),
.B(n_768),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1011),
.B(n_825),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_1024),
.B(n_301),
.C(n_302),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_974),
.A2(n_816),
.B(n_835),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_974),
.A2(n_820),
.B(n_816),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_859),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_SL g1047 ( 
.A(n_864),
.B(n_336),
.C(n_311),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_914),
.A2(n_809),
.B(n_839),
.C(n_825),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_930),
.B(n_839),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_990),
.A2(n_713),
.B(n_768),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_914),
.A2(n_825),
.B(n_768),
.C(n_217),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_842),
.B(n_298),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1012),
.B(n_713),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_915),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_876),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_876),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_R g1057 ( 
.A(n_884),
.B(n_768),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_882),
.A2(n_768),
.B(n_778),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_854),
.A2(n_713),
.B(n_335),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1012),
.B(n_713),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_SL g1061 ( 
.A(n_887),
.B(n_345),
.C(n_340),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1015),
.B(n_778),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_863),
.B(n_309),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_895),
.B(n_851),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1015),
.B(n_778),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_907),
.B(n_310),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_868),
.B(n_778),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_934),
.A2(n_975),
.B(n_866),
.C(n_1021),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_868),
.B(n_778),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_933),
.B(n_311),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1017),
.B(n_312),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_870),
.B(n_860),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_898),
.B(n_312),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_885),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_927),
.B(n_329),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_335),
.B(n_309),
.C(n_321),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_983),
.A2(n_337),
.B(n_344),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_917),
.A2(n_323),
.B(n_344),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_847),
.A2(n_342),
.B(n_334),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_927),
.B(n_844),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_890),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_855),
.A2(n_342),
.B(n_334),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_896),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_901),
.A2(n_323),
.B(n_463),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_857),
.B(n_904),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_940),
.A2(n_224),
.B1(n_463),
.B2(n_336),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_909),
.A2(n_339),
.B(n_332),
.C(n_13),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_904),
.B(n_339),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_986),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_969),
.A2(n_332),
.B1(n_103),
.B2(n_172),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_993),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_937),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_969),
.A2(n_463),
.B(n_150),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_895),
.B(n_148),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_972),
.B(n_11),
.C(n_17),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_986),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_857),
.B(n_908),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_843),
.A2(n_463),
.B(n_145),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_985),
.B(n_143),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_930),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_909),
.A2(n_18),
.B(n_19),
.C(n_22),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_L g1103 ( 
.A(n_954),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_953),
.B(n_23),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_954),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_921),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1025),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_947),
.A2(n_967),
.B(n_962),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_935),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_924),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_924),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_886),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_953),
.B(n_34),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1022),
.B(n_35),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_911),
.B(n_36),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_911),
.A2(n_938),
.B(n_985),
.C(n_913),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1019),
.B(n_38),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1010),
.B(n_39),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1025),
.A2(n_40),
.B(n_41),
.C(n_44),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_858),
.B(n_41),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_848),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_1005),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_867),
.B(n_47),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_846),
.A2(n_84),
.B(n_126),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_991),
.A2(n_49),
.B(n_52),
.C(n_54),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_939),
.A2(n_88),
.B1(n_119),
.B2(n_108),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_1005),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1005),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_865),
.A2(n_78),
.B(n_102),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_852),
.B(n_72),
.Y(n_1130)
);

AND2x6_ASAP7_75t_L g1131 ( 
.A(n_861),
.B(n_954),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_869),
.B(n_49),
.Y(n_1132)
);

OAI22x1_ASAP7_75t_L g1133 ( 
.A1(n_1023),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1005),
.Y(n_1134)
);

CKINVDCx8_ASAP7_75t_R g1135 ( 
.A(n_963),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1023),
.B(n_56),
.C(n_62),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_873),
.A2(n_91),
.B(n_96),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_852),
.B(n_63),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_879),
.B(n_65),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_SL g1140 ( 
.A1(n_862),
.A2(n_922),
.B(n_932),
.C(n_912),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1026),
.A2(n_65),
.B1(n_66),
.B2(n_81),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1029),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_941),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_955),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_849),
.A2(n_89),
.B(n_92),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_961),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_852),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_963),
.B(n_141),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_955),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_856),
.A2(n_943),
.B1(n_956),
.B2(n_893),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_893),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_856),
.B(n_893),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_856),
.B(n_968),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_976),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_916),
.B(n_959),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_998),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_963),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_963),
.B(n_916),
.Y(n_1159)
);

AND2x4_ASAP7_75t_SL g1160 ( 
.A(n_982),
.B(n_989),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_991),
.A2(n_897),
.B(n_1018),
.C(n_900),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_992),
.B(n_988),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_906),
.A2(n_994),
.B1(n_925),
.B2(n_1027),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_976),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_992),
.B(n_919),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_957),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1006),
.A2(n_920),
.B1(n_942),
.B2(n_936),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1007),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_948),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_853),
.A2(n_949),
.B(n_944),
.C(n_996),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1020),
.B(n_1028),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1006),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_923),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_850),
.A2(n_877),
.B(n_977),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_928),
.A2(n_918),
.B(n_880),
.C(n_888),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1020),
.B(n_958),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_978),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_949),
.A2(n_853),
.B1(n_944),
.B2(n_919),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_964),
.A2(n_966),
.B(n_881),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1009),
.B(n_1030),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1097),
.B(n_905),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1085),
.A2(n_883),
.B(n_987),
.C(n_926),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1034),
.A2(n_892),
.B(n_910),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1159),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1050),
.A2(n_999),
.B(n_878),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1172),
.A2(n_894),
.B1(n_902),
.B2(n_889),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1034),
.A2(n_903),
.B(n_899),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1179),
.A2(n_952),
.B(n_960),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1108),
.A2(n_872),
.B(n_891),
.Y(n_1189)
);

CKINVDCx6p67_ASAP7_75t_R g1190 ( 
.A(n_1089),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1031),
.A2(n_1002),
.B1(n_950),
.B2(n_951),
.C(n_875),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1068),
.A2(n_970),
.B(n_931),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1039),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1054),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1121),
.A2(n_997),
.B(n_996),
.C(n_1001),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1179),
.A2(n_945),
.B(n_871),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1036),
.A2(n_1016),
.B(n_1002),
.C(n_979),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1088),
.B(n_946),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1146),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1108),
.A2(n_980),
.B(n_981),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1096),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1150),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1072),
.B(n_1070),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1172),
.A2(n_984),
.B1(n_995),
.B2(n_1001),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1038),
.A2(n_1014),
.B(n_1013),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1046),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1135),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1166),
.B(n_1177),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1174),
.A2(n_997),
.B(n_874),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1175),
.A2(n_1000),
.A3(n_1003),
.B(n_1004),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1173),
.B(n_874),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1172),
.A2(n_1008),
.B1(n_1042),
.B2(n_1104),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1152),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1161),
.A2(n_1140),
.B(n_1080),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1121),
.A2(n_1117),
.B(n_1113),
.C(n_1061),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1114),
.A2(n_1095),
.B1(n_1075),
.B2(n_1047),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_1116),
.A2(n_1115),
.B(n_1094),
.C(n_1171),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1172),
.A2(n_1161),
.B(n_1060),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1053),
.A2(n_1033),
.B(n_1180),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1044),
.A2(n_1045),
.B(n_1168),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1164),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1032),
.A2(n_1167),
.B(n_1059),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1099),
.A2(n_1059),
.A3(n_1093),
.B(n_1151),
.Y(n_1223)
);

AOI221x1_ASAP7_75t_L g1224 ( 
.A1(n_1099),
.A2(n_1082),
.B1(n_1093),
.B2(n_1133),
.C(n_1090),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1169),
.B(n_1064),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1058),
.A2(n_1044),
.B(n_1162),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1103),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1103),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1055),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1157),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1043),
.A2(n_1138),
.B1(n_1071),
.B2(n_1112),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1052),
.B(n_1073),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1155),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1176),
.B(n_1118),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1066),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1037),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1067),
.A2(n_1069),
.B(n_1170),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1091),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1092),
.A2(n_1087),
.B(n_1076),
.C(n_1107),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1056),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1074),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1098),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1040),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1035),
.B(n_1142),
.Y(n_1244)
);

AO32x2_ASAP7_75t_L g1245 ( 
.A1(n_1126),
.A2(n_1107),
.A3(n_1119),
.B1(n_1087),
.B2(n_1102),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1084),
.A2(n_1163),
.B(n_1048),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_1137),
.B(n_1129),
.Y(n_1247)
);

BUFx12f_ASAP7_75t_L g1248 ( 
.A(n_1127),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1035),
.B(n_1153),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1136),
.A2(n_1100),
.B1(n_1035),
.B2(n_1123),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1119),
.A2(n_1102),
.B(n_1139),
.C(n_1132),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1154),
.A2(n_1065),
.B(n_1062),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1120),
.B(n_1128),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1147),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1122),
.B(n_1134),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1082),
.A2(n_1129),
.A3(n_1137),
.B(n_1077),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1178),
.A2(n_1156),
.B1(n_1158),
.B2(n_1143),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_1148),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1077),
.A2(n_1078),
.A3(n_1145),
.B(n_1079),
.Y(n_1259)
);

AO21x1_ASAP7_75t_L g1260 ( 
.A1(n_1125),
.A2(n_1051),
.B(n_1048),
.Y(n_1260)
);

AO22x2_ASAP7_75t_L g1261 ( 
.A1(n_1078),
.A2(n_1110),
.B1(n_1111),
.B2(n_1063),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1079),
.A2(n_1083),
.A3(n_1106),
.B(n_1081),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1160),
.A2(n_1130),
.B(n_1165),
.Y(n_1263)
);

AOI221xp5_ASAP7_75t_L g1264 ( 
.A1(n_1125),
.A2(n_1141),
.B1(n_1051),
.B2(n_1109),
.C(n_1086),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1159),
.B(n_1149),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1124),
.A2(n_1148),
.B(n_1049),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1049),
.A2(n_1144),
.B(n_1131),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_SL g1268 ( 
.A1(n_1131),
.A2(n_1124),
.B(n_1127),
.C(n_1057),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1105),
.A2(n_1131),
.A3(n_1041),
.B1(n_1101),
.B2(n_1040),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1131),
.Y(n_1270)
);

AO21x1_ASAP7_75t_L g1271 ( 
.A1(n_1085),
.A2(n_1115),
.B(n_971),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1272)
);

OAI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1172),
.A2(n_1024),
.B1(n_598),
.B2(n_635),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1159),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1097),
.B(n_841),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1068),
.A2(n_1038),
.B(n_1085),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1097),
.B(n_841),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1175),
.A2(n_846),
.A3(n_1174),
.B(n_1179),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1097),
.B(n_841),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1031),
.A2(n_971),
.B1(n_1117),
.B2(n_841),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1175),
.A2(n_846),
.A3(n_1174),
.B(n_1179),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1031),
.A2(n_971),
.B1(n_1117),
.B2(n_841),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1039),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1046),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1097),
.B(n_841),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1097),
.B(n_841),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1174),
.A2(n_1179),
.B(n_1175),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1172),
.A2(n_1085),
.B1(n_636),
.B2(n_971),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1175),
.A2(n_846),
.A3(n_1174),
.B(n_1179),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1039),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1039),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1146),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1097),
.B(n_841),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1097),
.B(n_841),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1050),
.A2(n_929),
.B(n_999),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_1105),
.B(n_676),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1046),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1039),
.Y(n_1302)
);

AO32x2_ASAP7_75t_L g1303 ( 
.A1(n_1033),
.A2(n_844),
.A3(n_1167),
.B1(n_1151),
.B2(n_1090),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1097),
.B(n_841),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1097),
.B(n_841),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1039),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1039),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1039),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1031),
.A2(n_971),
.B1(n_864),
.B2(n_745),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1072),
.B(n_842),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1050),
.A2(n_929),
.B(n_999),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1097),
.B(n_681),
.C(n_841),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1097),
.B(n_841),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_SL g1319 ( 
.A(n_1043),
.B(n_681),
.C(n_841),
.Y(n_1319)
);

O2A1O1Ixp5_ASAP7_75t_L g1320 ( 
.A1(n_1032),
.A2(n_841),
.B(n_971),
.C(n_1180),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1135),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1097),
.B(n_681),
.C(n_841),
.Y(n_1322)
);

AO22x2_ASAP7_75t_L g1323 ( 
.A1(n_1061),
.A2(n_971),
.B1(n_844),
.B2(n_1017),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1135),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1050),
.A2(n_929),
.B(n_999),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1039),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1041),
.B(n_1057),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_SL g1328 ( 
.A(n_1135),
.B(n_749),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1034),
.A2(n_630),
.B(n_546),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1097),
.B(n_841),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1097),
.B(n_686),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1072),
.B(n_842),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1201),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1283),
.A2(n_1285),
.B1(n_1314),
.B2(n_1317),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1283),
.A2(n_1285),
.B1(n_1317),
.B2(n_1322),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1322),
.A2(n_1296),
.B1(n_1307),
.B2(n_1330),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1312),
.Y(n_1337)
);

CKINVDCx6p67_ASAP7_75t_R g1338 ( 
.A(n_1227),
.Y(n_1338)
);

BUFx10_ASAP7_75t_L g1339 ( 
.A(n_1321),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1216),
.A2(n_1231),
.B(n_1331),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1291),
.A2(n_1288),
.B1(n_1275),
.B2(n_1318),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1269),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1278),
.A2(n_1280),
.B1(n_1305),
.B2(n_1289),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1233),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1199),
.Y(n_1345)
);

OAI22x1_ASAP7_75t_SL g1346 ( 
.A1(n_1238),
.A2(n_1293),
.B1(n_1286),
.B2(n_1221),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1291),
.A2(n_1231),
.B1(n_1319),
.B2(n_1297),
.Y(n_1347)
);

NAND2x1p5_ASAP7_75t_L g1348 ( 
.A(n_1328),
.B(n_1267),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1326),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1235),
.A2(n_1232),
.B1(n_1249),
.B2(n_1244),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1277),
.A2(n_1216),
.B1(n_1273),
.B2(n_1260),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1293),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1250),
.A2(n_1234),
.B1(n_1253),
.B2(n_1323),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1202),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1294),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1321),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1311),
.Y(n_1358)
);

INVx3_ASAP7_75t_SL g1359 ( 
.A(n_1321),
.Y(n_1359)
);

BUFx4_ASAP7_75t_SL g1360 ( 
.A(n_1207),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1277),
.A2(n_1323),
.B1(n_1271),
.B2(n_1264),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1184),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1230),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1250),
.A2(n_1225),
.B1(n_1315),
.B2(n_1332),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1269),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1324),
.B(n_1228),
.Y(n_1366)
);

CKINVDCx6p67_ASAP7_75t_R g1367 ( 
.A(n_1248),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1295),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1224),
.A2(n_1198),
.B1(n_1211),
.B2(n_1214),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1246),
.A2(n_1214),
.B1(n_1181),
.B2(n_1290),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1324),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1190),
.Y(n_1372)
);

OAI21xp33_ASAP7_75t_L g1373 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1239),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1236),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1194),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1246),
.A2(n_1258),
.B1(n_1266),
.B2(n_1212),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1191),
.A2(n_1212),
.B1(n_1213),
.B2(n_1222),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1240),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1241),
.A2(n_1242),
.B1(n_1258),
.B2(n_1218),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1193),
.A2(n_1310),
.B1(n_1302),
.B2(n_1254),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1255),
.A2(n_1257),
.B1(n_1287),
.B2(n_1229),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1206),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1301),
.A2(n_1261),
.B1(n_1237),
.B2(n_1184),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1262),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1327),
.A2(n_1274),
.B1(n_1300),
.B2(n_1217),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1262),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1245),
.A2(n_1265),
.B1(n_1300),
.B2(n_1270),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1263),
.A2(n_1261),
.B1(n_1186),
.B2(n_1204),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1243),
.A2(n_1219),
.B1(n_1245),
.B2(n_1204),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1243),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1243),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1247),
.A2(n_1245),
.B1(n_1205),
.B2(n_1303),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1195),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1279),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1268),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1220),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1182),
.A2(n_1197),
.B1(n_1226),
.B2(n_1304),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1192),
.A2(n_1205),
.B1(n_1252),
.B2(n_1187),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1303),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1209),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1192),
.A2(n_1189),
.B1(n_1303),
.B2(n_1298),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1259),
.B(n_1284),
.Y(n_1402)
);

BUFx10_ASAP7_75t_L g1403 ( 
.A(n_1320),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1272),
.A2(n_1282),
.B1(n_1329),
.B2(n_1313),
.Y(n_1404)
);

CKINVDCx14_ASAP7_75t_R g1405 ( 
.A(n_1256),
.Y(n_1405)
);

INVx5_ASAP7_75t_L g1406 ( 
.A(n_1292),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1276),
.A2(n_1281),
.B(n_1309),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1223),
.Y(n_1408)
);

BUFx2_ASAP7_75t_R g1409 ( 
.A(n_1223),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1223),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1306),
.A2(n_1308),
.B1(n_1183),
.B2(n_1196),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1188),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1200),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1210),
.Y(n_1414)
);

CKINVDCx11_ASAP7_75t_R g1415 ( 
.A(n_1210),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1210),
.B(n_1299),
.Y(n_1416)
);

BUFx12f_ASAP7_75t_L g1417 ( 
.A(n_1316),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1325),
.A2(n_1024),
.B1(n_686),
.B2(n_681),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1185),
.A2(n_971),
.B1(n_1285),
.B2(n_1283),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1233),
.Y(n_1420)
);

OAI21xp33_ASAP7_75t_L g1421 ( 
.A1(n_1283),
.A2(n_1285),
.B(n_681),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1283),
.A2(n_971),
.B1(n_1285),
.B2(n_1314),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1321),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1199),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1233),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1199),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1269),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1283),
.A2(n_971),
.B1(n_1285),
.B2(n_1314),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1199),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1233),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1283),
.A2(n_971),
.B1(n_1285),
.B2(n_1314),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1317),
.A2(n_1024),
.B1(n_686),
.B2(n_681),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1233),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1293),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1317),
.A2(n_1024),
.B1(n_686),
.B2(n_681),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1199),
.Y(n_1436)
);

BUFx10_ASAP7_75t_L g1437 ( 
.A(n_1321),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1283),
.A2(n_971),
.B1(n_1285),
.B2(n_1314),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1283),
.A2(n_971),
.B1(n_1285),
.B2(n_1314),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1199),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1283),
.A2(n_1285),
.B1(n_1024),
.B2(n_1172),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_1321),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1233),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1233),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1275),
.B(n_1278),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1199),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1312),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1233),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1317),
.A2(n_1024),
.B1(n_686),
.B2(n_681),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_SL g1450 ( 
.A(n_1221),
.Y(n_1450)
);

CKINVDCx11_ASAP7_75t_R g1451 ( 
.A(n_1233),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1199),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1269),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1417),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1399),
.B(n_1342),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1345),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1342),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1432),
.A2(n_1449),
.B1(n_1435),
.B2(n_1352),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1407),
.A2(n_1369),
.B(n_1441),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1369),
.A2(n_1441),
.B(n_1397),
.Y(n_1460)
);

INVxp33_ASAP7_75t_L g1461 ( 
.A(n_1447),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1344),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1355),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1393),
.A2(n_1421),
.B(n_1416),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1352),
.A2(n_1428),
.B1(n_1439),
.B2(n_1438),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1387),
.A2(n_1388),
.B(n_1412),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1351),
.A2(n_1395),
.B1(n_1389),
.B2(n_1336),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1396),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1406),
.B(n_1400),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1358),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1356),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1350),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1353),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1430),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1401),
.A2(n_1361),
.B(n_1398),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1384),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1401),
.A2(n_1361),
.B(n_1398),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1402),
.B(n_1394),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1386),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1399),
.B(n_1365),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1343),
.B(n_1445),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1434),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1422),
.A2(n_1431),
.B1(n_1438),
.B2(n_1439),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1363),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1340),
.B(n_1349),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1422),
.A2(n_1431),
.B1(n_1428),
.B2(n_1334),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1348),
.Y(n_1487)
);

AO21x1_ASAP7_75t_SL g1488 ( 
.A1(n_1334),
.A2(n_1335),
.B(n_1373),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1341),
.B(n_1364),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1425),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1341),
.B(n_1364),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1374),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1365),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1378),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1387),
.A2(n_1381),
.B(n_1354),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1365),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1365),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1370),
.B(n_1427),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1427),
.B(n_1453),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1427),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1453),
.B(n_1405),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1348),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1453),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1453),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1380),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1347),
.B(n_1335),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1347),
.A2(n_1418),
.B(n_1377),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1414),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1368),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1405),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1424),
.Y(n_1511)
);

AOI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1426),
.A2(n_1429),
.B(n_1446),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1413),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1436),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1440),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1395),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1377),
.A2(n_1419),
.B(n_1376),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1370),
.B(n_1419),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1395),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1452),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1375),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1415),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1408),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1409),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1381),
.A2(n_1379),
.B1(n_1346),
.B2(n_1385),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1392),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1383),
.A2(n_1379),
.B(n_1382),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1410),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1403),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1337),
.B(n_1333),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1403),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1383),
.B(n_1362),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1458),
.A2(n_1371),
.B1(n_1423),
.B2(n_1359),
.C(n_1433),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1485),
.B(n_1443),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1455),
.B(n_1411),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1455),
.B(n_1404),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1507),
.A2(n_1366),
.B(n_1391),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_SL g1538 ( 
.A(n_1495),
.B(n_1460),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1517),
.A2(n_1423),
.B(n_1359),
.C(n_1444),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1481),
.B(n_1366),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1448),
.Y(n_1541)
);

OAI211xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1505),
.A2(n_1451),
.B(n_1360),
.C(n_1338),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1488),
.A2(n_1420),
.B1(n_1450),
.B2(n_1357),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1471),
.B(n_1357),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1461),
.B(n_1450),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1498),
.B(n_1367),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1457),
.Y(n_1547)
);

OAI21xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1525),
.A2(n_1390),
.B(n_1339),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1506),
.B(n_1473),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1486),
.A2(n_1339),
.B(n_1437),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1465),
.A2(n_1437),
.B(n_1442),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1482),
.B(n_1372),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1498),
.B(n_1372),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1480),
.B(n_1499),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1484),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1468),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1480),
.B(n_1499),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1509),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1515),
.Y(n_1559)
);

BUFx4f_ASAP7_75t_SL g1560 ( 
.A(n_1474),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1457),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1454),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1483),
.A2(n_1489),
.B(n_1491),
.C(n_1460),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1487),
.B(n_1502),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1460),
.A2(n_1469),
.B(n_1459),
.Y(n_1565)
);

AND2x4_ASAP7_75t_SL g1566 ( 
.A(n_1519),
.B(n_1516),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1510),
.B(n_1478),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1472),
.B(n_1530),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1488),
.A2(n_1467),
.B1(n_1528),
.B2(n_1522),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1487),
.B(n_1502),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1495),
.A2(n_1524),
.B1(n_1475),
.B2(n_1477),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1528),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1476),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1513),
.B(n_1470),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1501),
.B(n_1510),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1501),
.B(n_1526),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1513),
.B(n_1456),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1479),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1479),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_SL g1580 ( 
.A1(n_1525),
.A2(n_1523),
.B(n_1522),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.B(n_1493),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1523),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1495),
.A2(n_1459),
.B1(n_1475),
.B2(n_1477),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1462),
.B(n_1490),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1512),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1512),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1469),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1524),
.A2(n_1518),
.B(n_1523),
.C(n_1522),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1469),
.B(n_1529),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1492),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1459),
.A2(n_1518),
.B1(n_1513),
.B2(n_1532),
.C(n_1529),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1516),
.A2(n_1519),
.B1(n_1531),
.B2(n_1475),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1527),
.A2(n_1516),
.B(n_1531),
.C(n_1519),
.Y(n_1595)
);

AND2x4_ASAP7_75t_SL g1596 ( 
.A(n_1590),
.B(n_1562),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1533),
.A2(n_1475),
.B1(n_1477),
.B2(n_1532),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1559),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1500),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1556),
.B(n_1564),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1538),
.A2(n_1477),
.B1(n_1466),
.B2(n_1519),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1558),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1580),
.A2(n_1466),
.B1(n_1519),
.B2(n_1516),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1554),
.B(n_1503),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1564),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1573),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1557),
.B(n_1503),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1580),
.A2(n_1466),
.B1(n_1502),
.B2(n_1464),
.Y(n_1610)
);

OAI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1593),
.A2(n_1520),
.B(n_1514),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1592),
.B(n_1464),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1567),
.B(n_1478),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1579),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1568),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1563),
.A2(n_1520),
.B1(n_1514),
.B2(n_1511),
.C(n_1463),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1591),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1577),
.B(n_1494),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1579),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1547),
.Y(n_1621)
);

AND2x4_ASAP7_75t_SL g1622 ( 
.A(n_1590),
.B(n_1454),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1570),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1575),
.B(n_1504),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1571),
.B(n_1494),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1556),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1575),
.B(n_1508),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1591),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1561),
.Y(n_1629)
);

BUFx8_ASAP7_75t_SL g1630 ( 
.A(n_1552),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1622),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1618),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1597),
.A2(n_1539),
.B(n_1543),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1614),
.B(n_1583),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1604),
.B(n_1583),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1599),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1617),
.B(n_1589),
.C(n_1569),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1602),
.B(n_1576),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1611),
.A2(n_1546),
.B1(n_1536),
.B2(n_1553),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1621),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1597),
.A2(n_1549),
.B1(n_1565),
.B2(n_1540),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1608),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1611),
.A2(n_1548),
.B1(n_1595),
.B2(n_1582),
.C(n_1572),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.B(n_1607),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1628),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1617),
.A2(n_1536),
.B1(n_1553),
.B2(n_1548),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1598),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1619),
.B(n_1538),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1603),
.A2(n_1537),
.B1(n_1576),
.B2(n_1551),
.Y(n_1653)
);

NOR2xp67_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1586),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1598),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1602),
.B(n_1535),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1619),
.B(n_1581),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1602),
.B(n_1535),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1629),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1616),
.A2(n_1550),
.B1(n_1534),
.B2(n_1542),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1622),
.A2(n_1594),
.B1(n_1587),
.B2(n_1566),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1598),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1622),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1651),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1651),
.B(n_1626),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1633),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1633),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1637),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1635),
.B(n_1612),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1613),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1655),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1631),
.B(n_1663),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1654),
.B(n_1613),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1654),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1644),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1639),
.A2(n_1645),
.B1(n_1653),
.B2(n_1642),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1662),
.B(n_1626),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1662),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1656),
.B(n_1600),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1644),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1646),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1663),
.B(n_1623),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1656),
.B(n_1606),
.Y(n_1690)
);

AOI21xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1639),
.A2(n_1584),
.B(n_1541),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1606),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1632),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1632),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1632),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1658),
.B(n_1609),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1632),
.B(n_1609),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1636),
.B(n_1620),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1687),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1683),
.A2(n_1645),
.B(n_1634),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1683),
.B(n_1638),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1687),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1694),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1691),
.B(n_1630),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_1636),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1677),
.B(n_1663),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1686),
.B(n_1659),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1699),
.B(n_1635),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1677),
.B(n_1648),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1668),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1699),
.B(n_1652),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1692),
.B(n_1641),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1668),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1665),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1716)
);

AOI32xp33_ASAP7_75t_L g1717 ( 
.A1(n_1677),
.A2(n_1653),
.A3(n_1650),
.B1(n_1661),
.B2(n_1660),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1686),
.B(n_1640),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1689),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1690),
.B(n_1640),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1665),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1668),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1677),
.B(n_1663),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1677),
.B(n_1648),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1677),
.B(n_1689),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1689),
.B(n_1698),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1669),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1665),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1664),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1665),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1692),
.B(n_1641),
.Y(n_1731)
);

NAND2x1_ASAP7_75t_L g1732 ( 
.A(n_1689),
.B(n_1632),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1669),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1690),
.B(n_1693),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1669),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1689),
.B(n_1632),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1674),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1670),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1679),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1670),
.Y(n_1740)
);

AOI322xp5_ASAP7_75t_L g1741 ( 
.A1(n_1691),
.A2(n_1625),
.A3(n_1610),
.B1(n_1647),
.B2(n_1664),
.C1(n_1605),
.C2(n_1624),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1689),
.B(n_1698),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1701),
.A2(n_1689),
.B1(n_1681),
.B2(n_1676),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1711),
.Y(n_1744)
);

AND3x2_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1739),
.C(n_1679),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1725),
.B(n_1675),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1702),
.B(n_1691),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1741),
.B(n_1690),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1717),
.B(n_1693),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1719),
.B(n_1710),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1714),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1700),
.B(n_1634),
.C(n_1694),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1707),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1693),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1714),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1727),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1732),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1727),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1733),
.Y(n_1761)
);

AOI211x1_ASAP7_75t_SL g1762 ( 
.A1(n_1706),
.A2(n_1696),
.B(n_1695),
.C(n_1694),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1732),
.A2(n_1667),
.B(n_1692),
.Y(n_1763)
);

NOR3xp33_ASAP7_75t_L g1764 ( 
.A(n_1703),
.B(n_1545),
.C(n_1544),
.Y(n_1764)
);

OAI21xp33_ASAP7_75t_L g1765 ( 
.A1(n_1709),
.A2(n_1671),
.B(n_1667),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1709),
.B(n_1697),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1725),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1734),
.B(n_1671),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1712),
.B(n_1697),
.Y(n_1769)
);

NAND2x1_ASAP7_75t_L g1770 ( 
.A(n_1725),
.B(n_1675),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1710),
.B(n_1697),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1712),
.B(n_1697),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1733),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1736),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1724),
.B(n_1695),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1716),
.B(n_1698),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1736),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1718),
.B(n_1720),
.Y(n_1779)
);

AND3x1_ASAP7_75t_L g1780 ( 
.A(n_1747),
.B(n_1742),
.C(n_1726),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1751),
.B(n_1707),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1751),
.B(n_1707),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1748),
.A2(n_1750),
.B1(n_1770),
.B2(n_1758),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1743),
.A2(n_1723),
.B1(n_1742),
.B2(n_1726),
.C(n_1703),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1758),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1753),
.A2(n_1723),
.B(n_1678),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1745),
.B(n_1729),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1755),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1749),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1763),
.A2(n_1765),
.B1(n_1778),
.B2(n_1775),
.C(n_1767),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1749),
.Y(n_1791)
);

OAI322xp33_ASAP7_75t_L g1792 ( 
.A1(n_1768),
.A2(n_1723),
.A3(n_1731),
.B1(n_1713),
.B2(n_1671),
.C1(n_1735),
.C2(n_1738),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1755),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1754),
.B(n_1704),
.Y(n_1794)
);

AOI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1754),
.A2(n_1695),
.B(n_1696),
.C(n_1704),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1752),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1746),
.A2(n_1676),
.B1(n_1681),
.B2(n_1675),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1746),
.A2(n_1676),
.B1(n_1681),
.B2(n_1675),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1774),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1752),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1756),
.Y(n_1801)
);

AOI321xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1762),
.A2(n_1671),
.A3(n_1713),
.B1(n_1731),
.B2(n_1698),
.C(n_1740),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1771),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1746),
.A2(n_1676),
.B1(n_1681),
.B2(n_1675),
.Y(n_1804)
);

AO21x1_ASAP7_75t_L g1805 ( 
.A1(n_1756),
.A2(n_1735),
.B(n_1722),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1789),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1789),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1780),
.A2(n_1770),
.B1(n_1764),
.B2(n_1776),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1781),
.B(n_1771),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1791),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1791),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1800),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1794),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1790),
.B(n_1779),
.Y(n_1814)
);

A2O1A1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1786),
.A2(n_1777),
.B(n_1768),
.C(n_1695),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1783),
.A2(n_1744),
.B(n_1759),
.C(n_1757),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1781),
.B(n_1774),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1800),
.Y(n_1818)
);

OAI322xp33_ASAP7_75t_L g1819 ( 
.A1(n_1802),
.A2(n_1766),
.A3(n_1773),
.B1(n_1761),
.B2(n_1769),
.C1(n_1772),
.C2(n_1760),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1787),
.B(n_1776),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1803),
.B(n_1761),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1795),
.B(n_1704),
.C(n_1773),
.Y(n_1822)
);

O2A1O1Ixp5_ASAP7_75t_L g1823 ( 
.A1(n_1792),
.A2(n_1696),
.B(n_1730),
.C(n_1728),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1782),
.B(n_1696),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1801),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1809),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1821),
.Y(n_1827)
);

AOI32xp33_ASAP7_75t_L g1828 ( 
.A1(n_1814),
.A2(n_1809),
.A3(n_1817),
.B1(n_1784),
.B2(n_1820),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1817),
.B(n_1785),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1813),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1824),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1816),
.B(n_1785),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1815),
.B(n_1799),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1815),
.B(n_1803),
.Y(n_1834)
);

XOR2xp5_ASAP7_75t_L g1835 ( 
.A(n_1808),
.B(n_1797),
.Y(n_1835)
);

OA21x2_ASAP7_75t_L g1836 ( 
.A1(n_1822),
.A2(n_1805),
.B(n_1801),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1821),
.Y(n_1837)
);

OAI31xp33_ASAP7_75t_L g1838 ( 
.A1(n_1833),
.A2(n_1794),
.A3(n_1782),
.B(n_1813),
.Y(n_1838)
);

AO21x1_ASAP7_75t_L g1839 ( 
.A1(n_1832),
.A2(n_1807),
.B(n_1806),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1828),
.A2(n_1819),
.B1(n_1823),
.B2(n_1825),
.C(n_1810),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1826),
.B(n_1829),
.Y(n_1841)
);

AOI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1834),
.A2(n_1818),
.B1(n_1812),
.B2(n_1811),
.C(n_1805),
.Y(n_1842)
);

AO21x1_ASAP7_75t_L g1843 ( 
.A1(n_1827),
.A2(n_1794),
.B(n_1796),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1836),
.A2(n_1824),
.B(n_1793),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1835),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1830),
.B(n_1831),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1840),
.A2(n_1836),
.B1(n_1837),
.B2(n_1804),
.C(n_1798),
.Y(n_1847)
);

O2A1O1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1842),
.A2(n_1793),
.B(n_1788),
.C(n_1737),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1845),
.Y(n_1849)
);

AOI321xp33_ASAP7_75t_L g1850 ( 
.A1(n_1846),
.A2(n_1788),
.A3(n_1737),
.B1(n_1730),
.B2(n_1728),
.C(n_1721),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1838),
.B(n_1704),
.Y(n_1851)
);

NAND3xp33_ASAP7_75t_SL g1852 ( 
.A(n_1849),
.B(n_1843),
.C(n_1839),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1847),
.A2(n_1844),
.B(n_1841),
.C(n_1704),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_L g1854 ( 
.A(n_1851),
.B(n_1721),
.C(n_1715),
.Y(n_1854)
);

NAND3xp33_ASAP7_75t_SL g1855 ( 
.A(n_1848),
.B(n_1560),
.C(n_1715),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_SL g1856 ( 
.A(n_1850),
.B(n_1678),
.C(n_1574),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1849),
.A2(n_1675),
.B1(n_1676),
.B2(n_1681),
.Y(n_1857)
);

NOR2x1p5_ASAP7_75t_L g1858 ( 
.A(n_1852),
.B(n_1562),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1855),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1857),
.Y(n_1860)
);

NAND4xp75_ASAP7_75t_L g1861 ( 
.A(n_1853),
.B(n_1678),
.C(n_1684),
.D(n_1666),
.Y(n_1861)
);

NOR3xp33_ASAP7_75t_L g1862 ( 
.A(n_1854),
.B(n_1562),
.C(n_1675),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1860),
.B(n_1856),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1860),
.A2(n_1688),
.B1(n_1670),
.B2(n_1673),
.C(n_1680),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1858),
.B(n_1672),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1865),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1866),
.Y(n_1867)
);

OAI22x1_ASAP7_75t_SL g1868 ( 
.A1(n_1867),
.A2(n_1859),
.B1(n_1866),
.B2(n_1863),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1867),
.Y(n_1869)
);

NAND2x1p5_ASAP7_75t_L g1870 ( 
.A(n_1869),
.B(n_1861),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1868),
.A2(n_1862),
.B1(n_1864),
.B2(n_1676),
.Y(n_1871)
);

OA21x2_ASAP7_75t_L g1872 ( 
.A1(n_1871),
.A2(n_1685),
.B(n_1674),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1870),
.A2(n_1674),
.B1(n_1685),
.B2(n_1682),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1872),
.B(n_1674),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1874),
.B(n_1873),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1875),
.A2(n_1676),
.B1(n_1681),
.B2(n_1673),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1876),
.A2(n_1673),
.B1(n_1688),
.B2(n_1680),
.C(n_1685),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1454),
.B(n_1688),
.C(n_1680),
.Y(n_1878)
);


endmodule