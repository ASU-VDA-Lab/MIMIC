module fake_jpeg_23477_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_24),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_18),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_5),
.B(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_16),
.B(n_14),
.Y(n_31)
);

FAx1_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_17),
.CI(n_16),
.CON(n_29),
.SN(n_29)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_29),
.A2(n_31),
.B(n_25),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_19),
.B1(n_15),
.B2(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_35),
.B1(n_28),
.B2(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_15),
.B1(n_11),
.B2(n_2),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_33),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_21),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_6),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_57),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_29),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_56),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_29),
.B1(n_38),
.B2(n_25),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_34),
.C(n_30),
.Y(n_64)
);

BUFx12f_ASAP7_75t_SL g59 ( 
.A(n_58),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_7),
.Y(n_66)
);

OAI322xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_44),
.A3(n_45),
.B1(n_42),
.B2(n_46),
.C1(n_34),
.C2(n_30),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_7),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.C(n_60),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_54),
.C(n_8),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_59),
.B(n_9),
.C(n_62),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_54),
.B(n_68),
.C(n_65),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_71),
.Y(n_74)
);


endmodule