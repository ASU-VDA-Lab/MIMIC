module fake_jpeg_23302_n_75 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_20),
.Y(n_22)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_19),
.B1(n_21),
.B2(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_R g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_21),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_13),
.B1(n_12),
.B2(n_19),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_11),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_11),
.B(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_29),
.C(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_50),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_53),
.B(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_8),
.B1(n_43),
.B2(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_8),
.B1(n_15),
.B2(n_4),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_59),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_47),
.C(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_43),
.C(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_40),
.C(n_52),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_64),
.B(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.C(n_67),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_41),
.B1(n_53),
.B2(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_61),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_41),
.A3(n_62),
.B1(n_39),
.B2(n_15),
.C1(n_5),
.C2(n_4),
.Y(n_73)
);

OAI321xp33_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_72),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_1),
.Y(n_75)
);


endmodule