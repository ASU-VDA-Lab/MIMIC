module fake_jpeg_14187_n_546 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_546);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_7),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_58),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_59),
.B(n_114),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_66),
.Y(n_180)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_67),
.Y(n_195)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_74),
.Y(n_189)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_42),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_78),
.B(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_21),
.B(n_0),
.CON(n_85),
.SN(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_1),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_96),
.A2(n_43),
.B1(n_34),
.B2(n_37),
.Y(n_187)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_106),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_4),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_117),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_31),
.B(n_4),
.Y(n_117)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_122),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_22),
.A2(n_4),
.B(n_5),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_24),
.B(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_50),
.Y(n_141)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_31),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_126),
.B(n_156),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_25),
.B1(n_49),
.B2(n_31),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_128),
.A2(n_164),
.B(n_201),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_60),
.A2(n_29),
.B1(n_33),
.B2(n_46),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_130),
.A2(n_172),
.B1(n_200),
.B2(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_141),
.B(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_50),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_106),
.C(n_94),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_153),
.B(n_165),
.C(n_137),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_38),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_38),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_161),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_62),
.B(n_24),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_160),
.B(n_186),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_63),
.B(n_40),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_61),
.A2(n_25),
.B1(n_49),
.B2(n_65),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_64),
.A2(n_49),
.B1(n_46),
.B2(n_45),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_167),
.A2(n_187),
.B1(n_196),
.B2(n_17),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_168),
.B(n_13),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_66),
.B(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_206),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_73),
.A2(n_45),
.B1(n_43),
.B2(n_33),
.Y(n_172)
);

INVx6_ASAP7_75t_SL g184 ( 
.A(n_72),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_96),
.B(n_41),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_74),
.A2(n_31),
.B1(n_37),
.B2(n_34),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_78),
.B(n_41),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_76),
.A2(n_40),
.B1(n_35),
.B2(n_42),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_79),
.A2(n_31),
.B(n_8),
.C(n_9),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_83),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_204),
.B1(n_128),
.B2(n_164),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_88),
.B(n_10),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_132),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_208),
.B(n_263),
.Y(n_315)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_210),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_121),
.B1(n_112),
.B2(n_111),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_213),
.A2(n_215),
.B1(n_218),
.B2(n_248),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_229),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_107),
.B1(n_100),
.B2(n_13),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_216),
.A2(n_231),
.B1(n_255),
.B2(n_266),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_131),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_225),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_226),
.Y(n_324)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_228),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_138),
.Y(n_229)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

BUFx24_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_232),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_135),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_234),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_130),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_238),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_145),
.Y(n_240)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_157),
.Y(n_242)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_135),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_243),
.A2(n_247),
.B1(n_249),
.B2(n_253),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_134),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_244),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_280)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_152),
.A2(n_202),
.B1(n_193),
.B2(n_185),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_125),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_167),
.A2(n_18),
.B1(n_165),
.B2(n_137),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_SL g310 ( 
.A(n_254),
.B(n_236),
.Y(n_310)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_256),
.Y(n_329)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_168),
.A2(n_146),
.B1(n_177),
.B2(n_140),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_258),
.A2(n_237),
.B(n_259),
.Y(n_326)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_142),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_152),
.A2(n_176),
.B1(n_202),
.B2(n_193),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_264),
.B1(n_268),
.B2(n_277),
.Y(n_294)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_150),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_185),
.A2(n_155),
.B1(n_174),
.B2(n_189),
.Y(n_264)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_266),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_267),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_171),
.A2(n_174),
.B1(n_181),
.B2(n_189),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_134),
.A2(n_140),
.B1(n_177),
.B2(n_192),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_139),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_171),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_148),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_180),
.A2(n_181),
.B1(n_190),
.B2(n_144),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_273),
.B(n_275),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_170),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_147),
.A2(n_154),
.B1(n_166),
.B2(n_180),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_154),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_283),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_224),
.A2(n_147),
.B1(n_175),
.B2(n_247),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_282),
.A2(n_295),
.B1(n_216),
.B2(n_249),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_220),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_254),
.B(n_220),
.CI(n_265),
.CON(n_290),
.SN(n_290)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_290),
.B(n_314),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_218),
.B(n_258),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_291),
.B(n_317),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_224),
.A2(n_217),
.B1(n_213),
.B2(n_215),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_216),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_319),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_211),
.B(n_246),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_321),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_210),
.C(n_275),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_260),
.B(n_246),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_251),
.B(n_221),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_212),
.B(n_208),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_230),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_326),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_288),
.A2(n_216),
.B1(n_241),
.B2(n_232),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_331),
.A2(n_349),
.B1(n_352),
.B2(n_359),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_333),
.A2(n_330),
.B1(n_301),
.B2(n_305),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_279),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_335),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_239),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_341),
.C(n_347),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_276),
.B(n_263),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_353),
.B(n_358),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_257),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_351),
.C(n_293),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_225),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_356),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_227),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_357),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_284),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_354),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_245),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_288),
.A2(n_250),
.B1(n_219),
.B2(n_223),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_313),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_350),
.B(n_365),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_209),
.C(n_226),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_295),
.A2(n_228),
.B1(n_252),
.B2(n_271),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_315),
.A2(n_262),
.B(n_272),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_286),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_302),
.A2(n_307),
.B1(n_322),
.B2(n_290),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_355),
.A2(n_362),
.B(n_369),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_287),
.B(n_256),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_317),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_315),
.A2(n_240),
.B(n_242),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_322),
.A2(n_280),
.B1(n_294),
.B2(n_311),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_306),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_364),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_325),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_371),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_325),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_299),
.A2(n_303),
.B(n_285),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_363),
.A2(n_367),
.B(n_323),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_296),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_303),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_281),
.B(n_292),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_347),
.C(n_342),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_312),
.A2(n_297),
.B(n_294),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_316),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_296),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_327),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_363),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_372),
.B(n_340),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_381),
.B1(n_387),
.B2(n_400),
.Y(n_408)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_361),
.Y(n_378)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_339),
.A2(n_296),
.B(n_301),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_385),
.B(n_397),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_355),
.A2(n_330),
.B1(n_305),
.B2(n_328),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_333),
.A2(n_332),
.B1(n_343),
.B2(n_362),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_331),
.A2(n_316),
.B1(n_327),
.B2(n_300),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_389),
.A2(n_401),
.B1(n_364),
.B2(n_370),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_289),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_391),
.B(n_386),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_332),
.B(n_293),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_402),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_398),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_339),
.A2(n_304),
.B(n_320),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_399),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_345),
.A2(n_298),
.B1(n_304),
.B2(n_320),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_298),
.B1(n_329),
.B2(n_323),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_341),
.B(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_337),
.A2(n_324),
.B1(n_345),
.B2(n_346),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_404),
.A2(n_344),
.B1(n_357),
.B2(n_349),
.Y(n_410)
);

OA22x2_ASAP7_75t_L g407 ( 
.A1(n_383),
.A2(n_339),
.B1(n_357),
.B2(n_367),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_412),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_383),
.A2(n_350),
.B1(n_338),
.B2(n_352),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_409),
.A2(n_417),
.B1(n_419),
.B2(n_392),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_410),
.A2(n_415),
.B1(n_427),
.B2(n_385),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_379),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_375),
.C(n_336),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_420),
.C(n_428),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_377),
.A2(n_353),
.B(n_358),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_425),
.Y(n_434)
);

OAI22x1_ASAP7_75t_L g415 ( 
.A1(n_372),
.A2(n_351),
.B1(n_344),
.B2(n_356),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_383),
.A2(n_338),
.B1(n_351),
.B2(n_344),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_366),
.C(n_360),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_421),
.B(n_384),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_373),
.B(n_340),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_432),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_424),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_377),
.A2(n_348),
.B(n_369),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_324),
.B1(n_369),
.B2(n_381),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_369),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_373),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_372),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_379),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_430),
.B(n_400),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_431),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_395),
.B(n_384),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_402),
.C(n_378),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_426),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_437),
.B(n_433),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_440),
.Y(n_463)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_450),
.C(n_428),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_409),
.A2(n_404),
.B1(n_376),
.B2(n_392),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_443),
.A2(n_444),
.B1(n_449),
.B2(n_458),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_422),
.B(n_386),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_447),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_424),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_448),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_408),
.A2(n_388),
.B1(n_393),
.B2(n_389),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_388),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_452),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_398),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_390),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_454),
.Y(n_479)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_411),
.Y(n_454)
);

OAI221xp5_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_391),
.B1(n_390),
.B2(n_399),
.C(n_392),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_457),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_401),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_456),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_417),
.A2(n_392),
.B1(n_380),
.B2(n_389),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_408),
.B1(n_432),
.B2(n_427),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_459),
.A2(n_405),
.B1(n_410),
.B2(n_411),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_462),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_429),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_454),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_420),
.C(n_415),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_476),
.C(n_436),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_468),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_451),
.B(n_405),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_472),
.Y(n_488)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_439),
.B(n_425),
.CI(n_414),
.CON(n_471),
.SN(n_471)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_474),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_406),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_406),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_480),
.Y(n_491)
);

FAx1_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_380),
.CI(n_407),
.CON(n_475),
.SN(n_475)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_458),
.B(n_456),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_407),
.C(n_397),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_407),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_482),
.A2(n_487),
.B(n_467),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_435),
.Y(n_483)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_435),
.B1(n_443),
.B2(n_444),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_484),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_493),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_463),
.A2(n_439),
.B1(n_453),
.B2(n_445),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_468),
.Y(n_500)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_495),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_449),
.C(n_437),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_492),
.B(n_494),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_460),
.B(n_441),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_374),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_469),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_481),
.A2(n_463),
.B1(n_473),
.B2(n_476),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_498),
.A2(n_499),
.B1(n_506),
.B2(n_509),
.Y(n_511)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_492),
.B(n_475),
.CI(n_471),
.CON(n_499),
.SN(n_499)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_487),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_489),
.Y(n_505)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_481),
.A2(n_467),
.B1(n_475),
.B2(n_471),
.Y(n_506)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_508),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_486),
.A2(n_477),
.B1(n_401),
.B2(n_480),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_516),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_485),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_514),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_494),
.C(n_485),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_493),
.C(n_491),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_515),
.B(n_465),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_491),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_488),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_519),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_488),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_518),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_522),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_505),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_503),
.C(n_507),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_527),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_502),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_528),
.B(n_529),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_500),
.B1(n_419),
.B2(n_472),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_511),
.Y(n_531)
);

AOI31xp33_ASAP7_75t_L g539 ( 
.A1(n_531),
.A2(n_532),
.A3(n_534),
.B(n_517),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_526),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_524),
.B(n_516),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_523),
.C(n_524),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_538),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_530),
.A2(n_533),
.B(n_499),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_537),
.A2(n_539),
.B(n_519),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_499),
.B(n_523),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_461),
.B(n_470),
.Y(n_542)
);

OAI321xp33_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_540),
.A3(n_461),
.B1(n_374),
.B2(n_396),
.C(n_423),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_543),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_423),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_382),
.Y(n_546)
);


endmodule