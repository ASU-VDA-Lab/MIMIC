module fake_jpeg_14727_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_33),
.B1(n_17),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_42),
.B1(n_23),
.B2(n_33),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_56),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_42),
.C(n_37),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_33),
.B1(n_23),
.B2(n_18),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_68),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_42),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_86),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_32),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_82),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_25),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_80),
.B1(n_95),
.B2(n_26),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_77),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_31),
.B1(n_32),
.B2(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_78),
.Y(n_99)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_92),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_18),
.B1(n_23),
.B2(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_27),
.Y(n_81)
);

XOR2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_32),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_59),
.B1(n_34),
.B2(n_35),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_19),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_21),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_36),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_31),
.B1(n_36),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_45),
.A2(n_31),
.B1(n_21),
.B2(n_26),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_122),
.B1(n_19),
.B2(n_22),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_26),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_95),
.B1(n_65),
.B2(n_89),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_62),
.B1(n_92),
.B2(n_88),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_139),
.B1(n_105),
.B2(n_113),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_87),
.B1(n_74),
.B2(n_62),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_93),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_130),
.C(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_69),
.C(n_66),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_144),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_78),
.B(n_66),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_136),
.B(n_140),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_94),
.B(n_91),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_22),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_22),
.B(n_2),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_116),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_1),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_98),
.B(n_14),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_1),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_11),
.C(n_10),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_101),
.B(n_120),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_159),
.B(n_163),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_122),
.B(n_99),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_96),
.B1(n_108),
.B2(n_117),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_154),
.B1(n_151),
.B2(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_115),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_119),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_146),
.B1(n_144),
.B2(n_133),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_137),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_179),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_186),
.Y(n_194)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_126),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_124),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_150),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_123),
.B1(n_131),
.B2(n_125),
.C(n_140),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_184),
.B(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_174),
.A2(n_153),
.B1(n_163),
.B2(n_150),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_199),
.B1(n_200),
.B2(n_3),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_179),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_160),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_176),
.C(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_197),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_198),
.B(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_165),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_153),
.B(n_149),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_164),
.B1(n_169),
.B2(n_131),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_164),
.B1(n_147),
.B2(n_121),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_182),
.C(n_178),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_205),
.B(n_210),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_203),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_172),
.C(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_121),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_2),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_212),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_3),
.C(n_4),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_191),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_211),
.A2(n_192),
.B1(n_198),
.B2(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

XNOR2x2_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_216),
.B1(n_206),
.B2(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_210),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_214),
.B(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_211),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_224),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_209),
.C(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_215),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_9),
.B(n_6),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_222),
.B(n_226),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_219),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_4),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_234),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_227),
.Y(n_238)
);


endmodule