module fake_jpeg_27657_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_30),
.B1(n_23),
.B2(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_54),
.B1(n_33),
.B2(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_30),
.B1(n_23),
.B2(n_15),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_35),
.B1(n_36),
.B2(n_28),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_29),
.B1(n_21),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_22),
.B1(n_19),
.B2(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_21),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_69),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_34),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_61),
.B(n_31),
.Y(n_85)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_34),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_67),
.B1(n_72),
.B2(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_74),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_14),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_35),
.B1(n_28),
.B2(n_16),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_77),
.B1(n_84),
.B2(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_44),
.B1(n_45),
.B2(n_41),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_89),
.B(n_92),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_92),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_44),
.B1(n_61),
.B2(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_57),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_52),
.B(n_53),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_73),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_69),
.C(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_63),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_79),
.B1(n_84),
.B2(n_91),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_52),
.B1(n_53),
.B2(n_16),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_121),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_84),
.A3(n_89),
.B1(n_79),
.B2(n_16),
.C1(n_14),
.C2(n_82),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_120),
.B(n_115),
.C(n_95),
.D(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_98),
.Y(n_129)
);

AO221x1_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_96),
.B1(n_104),
.B2(n_75),
.C(n_52),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_133),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_119),
.A3(n_121),
.B1(n_116),
.B2(n_114),
.C(n_110),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_129),
.Y(n_136)
);

NAND4xp25_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_97),
.C(n_99),
.D(n_102),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_135),
.B1(n_3),
.B2(n_4),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_106),
.C(n_97),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_110),
.C(n_116),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_140),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_136),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_75),
.C(n_53),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_8),
.C(n_9),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_13),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_125),
.B(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_144),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_128),
.C(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_156),
.B1(n_148),
.B2(n_5),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_12),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_151),
.A2(n_133),
.B1(n_125),
.B2(n_9),
.Y(n_156)
);

NAND2x1_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

OAI221xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_4),
.B1(n_5),
.B2(n_12),
.C(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_154),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_155),
.C(n_4),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_161),
.Y(n_167)
);


endmodule