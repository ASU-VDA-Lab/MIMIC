module real_jpeg_27907_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_286;
wire n_288;
wire n_292;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_0),
.A2(n_40),
.B1(n_47),
.B2(n_51),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_77),
.B1(n_78),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_1),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_125),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_1),
.A2(n_47),
.B1(n_51),
.B2(n_125),
.Y(n_229)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_2),
.A2(n_112),
.B(n_170),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_4),
.A2(n_77),
.B1(n_78),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_4),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_153),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_4),
.A2(n_47),
.B1(n_51),
.B2(n_153),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_44),
.B1(n_47),
.B2(n_51),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_44),
.B1(n_77),
.B2(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_164)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_8),
.A2(n_11),
.B(n_47),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_38),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_9),
.A2(n_38),
.B1(n_47),
.B2(n_51),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_47),
.B1(n_51),
.B2(n_58),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_11),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_27),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_27),
.B(n_194),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_151),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_11),
.B(n_119),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_11),
.A2(n_89),
.B1(n_90),
.B2(n_242),
.Y(n_244)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_15),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_15),
.A2(n_77),
.B1(n_78),
.B2(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_15),
.A2(n_47),
.B1(n_51),
.B2(n_147),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_101),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_60),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_25),
.B(n_70),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_25),
.A2(n_30),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_25),
.A2(n_30),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_25),
.A2(n_30),
.B1(n_179),
.B2(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_27),
.A2(n_28),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_27),
.B(n_74),
.Y(n_167)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_28),
.A2(n_81),
.B1(n_150),
.B2(n_167),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_28),
.A2(n_32),
.A3(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_30),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_30)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_31),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_31),
.B(n_33),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_33),
.B1(n_50),
.B2(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_33),
.A2(n_50),
.B(n_151),
.C(n_221),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_37),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_42),
.A2(n_55),
.B(n_202),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_55),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_46),
.A2(n_55),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_46),
.A2(n_53),
.B(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_46),
.A2(n_55),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_46),
.A2(n_55),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_46),
.A2(n_55),
.B1(n_201),
.B2(n_219),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_46),
.B(n_151),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_90),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_51),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_55),
.A2(n_64),
.B(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_67),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_67),
.A2(n_69),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_83),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_72),
.A2(n_123),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_72),
.B(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_72),
.A2(n_123),
.B1(n_124),
.B2(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.C(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_73),
.A2(n_80),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_78),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_78),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_94),
.B(n_98),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_98),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_88),
.A2(n_95),
.B1(n_105),
.B2(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_92),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_89),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_89),
.A2(n_90),
.B1(n_138),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_89),
.A2(n_114),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_89),
.A2(n_91),
.B1(n_234),
.B2(n_242),
.Y(n_241)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_90),
.B(n_151),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_93),
.A2(n_140),
.B(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_102),
.B(n_106),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_107),
.A2(n_108),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.C(n_121),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_109),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_110),
.B(n_116),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_115),
.A2(n_191),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_118),
.Y(n_291)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_297),
.B(n_302),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_284),
.B(n_296),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_183),
.B(n_265),
.C(n_283),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_171),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_133),
.B(n_171),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_154),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_135),
.B(n_141),
.C(n_154),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_136),
.B(n_137),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_149),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_156),
.B(n_161),
.C(n_165),
.Y(n_281)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_164),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_168),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_172),
.A2(n_173),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_181),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_207),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_264),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_257),
.B(n_263),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_212),
.B(n_256),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_203),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_187),
.B(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.C(n_199),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_189),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_204),
.B(n_210),
.C(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_250),
.B(n_255),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_230),
.B(n_249),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_238),
.B(n_248),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_236),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_243),
.B(n_247),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_281),
.B2(n_282),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_273),
.C(n_282),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_276),
.C(n_279),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_295),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_293),
.C(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);


endmodule