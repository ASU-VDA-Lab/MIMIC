module fake_jpeg_29148_n_48 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_48);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx12_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_25),
.B1(n_0),
.B2(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_27),
.B(n_2),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_25),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_21),
.B(n_19),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_21),
.C(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_39),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_21),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_32),
.B1(n_38),
.B2(n_6),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_3),
.Y(n_44)
);

NOR2xp67_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_41),
.C(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_6),
.Y(n_48)
);


endmodule