module fake_netlist_5_343_n_1567 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1567);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1567;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_92),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_20),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_33),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_61),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_117),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_46),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_67),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_54),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_68),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_32),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_88),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_45),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_25),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_19),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_77),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_97),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_105),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_62),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_76),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_144),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_94),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_120),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_147),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_17),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_122),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_126),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_151),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_12),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_53),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_34),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_20),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_111),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_87),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_9),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_22),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_29),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_38),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_145),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_91),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_27),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_139),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_52),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_137),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_32),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_84),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_29),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_25),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_6),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_71),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_90),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_119),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_85),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_127),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_51),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_86),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_24),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_134),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_79),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_10),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_8),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_72),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_60),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_30),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_37),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_133),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_65),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_103),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_150),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_82),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_140),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_96),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_39),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_19),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_18),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_108),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_12),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_48),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_35),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_93),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_7),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_109),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_40),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_143),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_23),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_74),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_78),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_63),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_3),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_115),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_22),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_135),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_104),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_80),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_98),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_21),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_41),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_159),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_201),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_159),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_167),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_305),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_305),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_155),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_153),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_236),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_167),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_169),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_233),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_156),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_233),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_172),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_229),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_237),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_172),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_172),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_166),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_221),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_161),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_174),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_231),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_179),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_170),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_221),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_170),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_231),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_192),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_231),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_152),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_194),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_152),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_205),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_162),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_221),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_205),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_194),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_163),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_280),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_168),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_299),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_203),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_210),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_192),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_171),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_180),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_216),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_173),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_214),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_217),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_176),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_192),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_249),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_279),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_291),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_307),
.Y(n_379)
);

NOR2x1_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_154),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_308),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_316),
.B(n_294),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_314),
.B(n_241),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_327),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_310),
.A2(n_160),
.B1(n_218),
.B2(n_234),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_177),
.Y(n_393)
);

BUFx12f_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_315),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_340),
.B(n_178),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_325),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_154),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_331),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_181),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_309),
.B(n_289),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_345),
.B(n_182),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_332),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_324),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_311),
.Y(n_416)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_368),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_335),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_346),
.B(n_175),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_351),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_356),
.Y(n_429)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_346),
.B(n_175),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_196),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_183),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_329),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_350),
.A2(n_164),
.B(n_158),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_362),
.B(n_184),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_359),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_394),
.Y(n_448)
);

INVx11_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_437),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_378),
.B(n_364),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_402),
.B(n_280),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_378),
.B(n_157),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_437),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_378),
.B(n_406),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_378),
.A2(n_297),
.B1(n_300),
.B2(n_292),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_406),
.B(n_369),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_386),
.B(n_365),
.Y(n_464)
);

INVx4_ASAP7_75t_SL g465 ( 
.A(n_417),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_384),
.B(n_157),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_393),
.B(n_373),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_381),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_384),
.B(n_157),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_424),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_334),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_192),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_388),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_186),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_397),
.B(n_187),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_397),
.B(n_188),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_435),
.B(n_157),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_440),
.B(n_336),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_440),
.B(n_165),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_396),
.B(n_399),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_404),
.B(n_185),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_334),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_404),
.B(n_190),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_412),
.Y(n_502)
);

CKINVDCx6p67_ASAP7_75t_R g503 ( 
.A(n_394),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_412),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_405),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_408),
.B(n_380),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_383),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_409),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_432),
.A2(n_352),
.B1(n_341),
.B2(n_313),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_426),
.B(n_338),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

AND3x2_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_320),
.C(n_319),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_408),
.B(n_189),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_380),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_413),
.B(n_191),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_392),
.B(n_321),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_382),
.B(n_193),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_415),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_383),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_428),
.B(n_320),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_382),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_429),
.B(n_372),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_430),
.B(n_417),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_382),
.B(n_195),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_416),
.B(n_323),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_427),
.B(n_208),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_427),
.B(n_212),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_418),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_427),
.B(n_219),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_431),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_382),
.B(n_198),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_382),
.B(n_339),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_436),
.B(n_192),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_422),
.B(n_160),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_392),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_439),
.B(n_372),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_423),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_423),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_436),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_414),
.B(n_342),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_414),
.B(n_421),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_414),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_431),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_434),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_434),
.B(n_377),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_414),
.B(n_199),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_414),
.B(n_200),
.Y(n_572)
);

INVx8_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_421),
.B(n_347),
.Y(n_574)
);

AO21x2_ASAP7_75t_L g575 ( 
.A1(n_439),
.A2(n_302),
.B(n_225),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_421),
.B(n_239),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_438),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_442),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_442),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_436),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_421),
.B(n_202),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_385),
.A2(n_247),
.B1(n_242),
.B2(n_264),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_421),
.B(n_355),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_385),
.B(n_390),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_563),
.A2(n_400),
.B(n_439),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_450),
.B(n_357),
.Y(n_588)
);

BUFx5_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_458),
.B(n_400),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_456),
.B(n_192),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_456),
.B(n_192),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_578),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_457),
.B(n_375),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_443),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_578),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_560),
.Y(n_597)
);

NOR2x1p5_ASAP7_75t_L g598 ( 
.A(n_503),
.B(n_197),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_468),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_443),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_478),
.A2(n_447),
.B1(n_451),
.B2(n_464),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_499),
.B(n_278),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_537),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_569),
.B(n_262),
.C(n_261),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_536),
.B(n_567),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_499),
.B(n_290),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_460),
.B(n_478),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_536),
.B(n_400),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_536),
.B(n_400),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_567),
.B(n_400),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_551),
.A2(n_562),
.B1(n_584),
.B2(n_574),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_206),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_579),
.Y(n_617)
);

BUFx5_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_517),
.B(n_204),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_567),
.B(n_433),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_452),
.A2(n_270),
.B1(n_223),
.B2(n_226),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_467),
.B(n_433),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_540),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_509),
.B(n_433),
.Y(n_624)
);

AND2x6_ASAP7_75t_SL g625 ( 
.A(n_491),
.B(n_375),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_557),
.A2(n_252),
.B1(n_244),
.B2(n_235),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_444),
.B(n_220),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_535),
.B(n_507),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_509),
.B(n_433),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_548),
.B(n_433),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_568),
.B(n_445),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_R g632 ( 
.A(n_452),
.B(n_207),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_481),
.B(n_441),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_489),
.A2(n_273),
.B1(n_211),
.B2(n_222),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_482),
.B(n_441),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_502),
.B(n_376),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_486),
.B(n_441),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_559),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_456),
.B(n_248),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_565),
.B(n_376),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_523),
.B(n_224),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_555),
.A2(n_252),
.B1(n_234),
.B2(n_218),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_534),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_566),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_557),
.A2(n_235),
.B1(n_244),
.B2(n_266),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_521),
.B(n_577),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_463),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_480),
.B(n_377),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_463),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_489),
.B(n_245),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_580),
.B(n_441),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_549),
.B(n_248),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_490),
.A2(n_390),
.B(n_420),
.C(n_403),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_459),
.A2(n_441),
.B(n_420),
.C(n_403),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_556),
.B(n_490),
.C(n_515),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_454),
.B(n_436),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_469),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_549),
.B(n_395),
.Y(n_658)
);

NAND2x1_ASAP7_75t_L g659 ( 
.A(n_549),
.B(n_395),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_557),
.A2(n_476),
.B1(n_494),
.B2(n_500),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_570),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_547),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_476),
.A2(n_401),
.B(n_398),
.C(n_246),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_549),
.B(n_248),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_494),
.B(n_253),
.Y(n_665)
);

NOR2xp67_ASAP7_75t_L g666 ( 
.A(n_538),
.B(n_398),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_500),
.B(n_256),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_585),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_540),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_564),
.B(n_248),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_487),
.B(n_401),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_487),
.B(n_213),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_530),
.B(n_228),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_484),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_471),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_473),
.B(n_257),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_473),
.B(n_498),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_520),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_539),
.B(n_230),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_484),
.B(n_232),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_550),
.B(n_238),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_571),
.B(n_240),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_243),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_475),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_582),
.B(n_250),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_484),
.B(n_251),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_466),
.B(n_254),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_528),
.Y(n_689)
);

CKINVDCx16_ASAP7_75t_R g690 ( 
.A(n_448),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_473),
.A2(n_265),
.B1(n_255),
.B2(n_304),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_472),
.B(n_263),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_485),
.B(n_272),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_556),
.B(n_258),
.Y(n_694)
);

OAI221xp5_ASAP7_75t_L g695 ( 
.A1(n_583),
.A2(n_285),
.B1(n_259),
.B2(n_260),
.C(n_268),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_473),
.B(n_306),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_485),
.B(n_286),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_498),
.B(n_269),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_498),
.B(n_366),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_542),
.B(n_287),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_485),
.B(n_284),
.Y(n_701)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_576),
.A2(n_446),
.B(n_453),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_455),
.B(n_298),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_461),
.B(n_276),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_449),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_498),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_448),
.B(n_366),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_474),
.B(n_296),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_576),
.B(n_544),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_557),
.A2(n_277),
.B1(n_295),
.B2(n_274),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_477),
.B(n_303),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_479),
.B(n_275),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_483),
.B(n_282),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_493),
.B(n_248),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_495),
.B(n_248),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_492),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_496),
.B(n_248),
.Y(n_717)
);

AO221x1_ASAP7_75t_L g718 ( 
.A1(n_497),
.A2(n_301),
.B1(n_229),
.B2(n_354),
.C(n_353),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_504),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_564),
.B(n_229),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_501),
.B(n_288),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_504),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_544),
.B(n_271),
.Y(n_723)
);

AND2x2_ASAP7_75t_SL g724 ( 
.A(n_553),
.B(n_360),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_516),
.B(n_283),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_546),
.B(n_281),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_448),
.B(n_503),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_505),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_546),
.B(n_301),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_564),
.B(n_301),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_505),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_518),
.B(n_360),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_522),
.B(n_358),
.Y(n_733)
);

INVxp33_ASAP7_75t_L g734 ( 
.A(n_466),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_575),
.A2(n_358),
.B1(n_354),
.B2(n_4),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_526),
.B(n_148),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_533),
.B(n_142),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_448),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_488),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_525),
.A2(n_141),
.B1(n_138),
.B2(n_130),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_545),
.B(n_0),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_575),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_488),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_607),
.Y(n_744)
);

BUFx12f_ASAP7_75t_L g745 ( 
.A(n_705),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_679),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_610),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_SL g748 ( 
.A1(n_642),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_646),
.B(n_531),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_SL g750 ( 
.A1(n_626),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_631),
.B(n_531),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_597),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_645),
.A2(n_541),
.B1(n_506),
.B2(n_511),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_690),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_602),
.B(n_465),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_665),
.A2(n_541),
.B(n_511),
.C(n_506),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_601),
.Y(n_757)
);

OAI21xp33_ASAP7_75t_L g758 ( 
.A1(n_645),
.A2(n_470),
.B(n_508),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_594),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_743),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_604),
.B(n_465),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_614),
.B(n_465),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_647),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_743),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_638),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_606),
.A2(n_573),
.B(n_586),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_644),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_599),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_735),
.A2(n_527),
.B1(n_513),
.B2(n_519),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_600),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_593),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_628),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_596),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_609),
.B(n_529),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_636),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_662),
.B(n_462),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_655),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_622),
.B(n_668),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_676),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_662),
.B(n_497),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_662),
.Y(n_781)
);

BUFx12f_ASAP7_75t_SL g782 ( 
.A(n_588),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_709),
.A2(n_665),
.B1(n_667),
.B2(n_597),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_603),
.B(n_513),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_590),
.B(n_519),
.Y(n_785)
);

AND2x6_ASAP7_75t_L g786 ( 
.A(n_678),
.B(n_709),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_649),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_667),
.A2(n_525),
.B1(n_462),
.B2(n_514),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_603),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_616),
.B(n_514),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_627),
.B(n_543),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

AND2x6_ASAP7_75t_SL g793 ( 
.A(n_650),
.B(n_16),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_735),
.A2(n_543),
.B1(n_524),
.B2(n_552),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_661),
.B(n_581),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_615),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_627),
.B(n_552),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_657),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_623),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_694),
.B(n_16),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_743),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_669),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_739),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_743),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_605),
.B(n_561),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_640),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_648),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_640),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_727),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_616),
.B(n_514),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_608),
.B(n_497),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_608),
.B(n_510),
.Y(n_812)
);

OR2x2_ASAP7_75t_SL g813 ( 
.A(n_617),
.B(n_561),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_643),
.B(n_21),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_716),
.Y(n_815)
);

AND2x2_ASAP7_75t_SL g816 ( 
.A(n_626),
.B(n_742),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_731),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_658),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_699),
.B(n_581),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_732),
.Y(n_820)
);

CKINVDCx11_ASAP7_75t_R g821 ( 
.A(n_625),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_675),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_724),
.B(n_532),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_724),
.B(n_532),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_674),
.B(n_510),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_632),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_729),
.A2(n_650),
.B(n_723),
.C(n_726),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_R g828 ( 
.A(n_700),
.B(n_59),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_675),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_733),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_589),
.B(n_586),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_689),
.B(n_23),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_660),
.A2(n_525),
.B1(n_586),
.B2(n_573),
.Y(n_833)
);

INVx5_ASAP7_75t_L g834 ( 
.A(n_707),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_641),
.B(n_28),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_619),
.B(n_641),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_721),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_651),
.Y(n_838)
);

AND2x6_ASAP7_75t_SL g839 ( 
.A(n_677),
.B(n_696),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_725),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_739),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_632),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_624),
.B(n_525),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_659),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_719),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_660),
.A2(n_525),
.B1(n_573),
.B2(n_34),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_629),
.B(n_573),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_633),
.B(n_58),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_635),
.B(n_66),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_706),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_729),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_SL g852 ( 
.A1(n_742),
.A2(n_695),
.B1(n_726),
.B2(n_723),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_637),
.B(n_83),
.Y(n_853)
);

CKINVDCx6p67_ASAP7_75t_R g854 ( 
.A(n_720),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_598),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_620),
.B(n_722),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_652),
.A2(n_31),
.B1(n_36),
.B2(n_42),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_728),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_677),
.B(n_42),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_696),
.B(n_698),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_702),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_698),
.B(n_43),
.Y(n_862)
);

INVx6_ASAP7_75t_L g863 ( 
.A(n_589),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_671),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_589),
.B(n_57),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_630),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_654),
.A2(n_43),
.B(n_44),
.C(n_73),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_672),
.Y(n_868)
);

INVx5_ASAP7_75t_L g869 ( 
.A(n_718),
.Y(n_869)
);

BUFx5_ASAP7_75t_L g870 ( 
.A(n_618),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_618),
.B(n_44),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_R g872 ( 
.A(n_706),
.B(n_738),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_618),
.B(n_613),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_653),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_670),
.A2(n_591),
.B1(n_592),
.B2(n_639),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_730),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_714),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_618),
.B(n_686),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_621),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_634),
.B(n_734),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_618),
.B(n_612),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_715),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_717),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_652),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_741),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_618),
.B(n_680),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_664),
.B(n_741),
.C(n_663),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_611),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_673),
.B(n_682),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_664),
.A2(n_670),
.B1(n_591),
.B2(n_592),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_710),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_683),
.B(n_684),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_666),
.B(n_692),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_656),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_691),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_587),
.A2(n_639),
.B(n_688),
.C(n_704),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_703),
.B(n_711),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_708),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_693),
.A2(n_697),
.B(n_701),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_712),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_736),
.A2(n_737),
.B(n_713),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_681),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_687),
.B(n_740),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_595),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_599),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_646),
.B(n_622),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_SL g907 ( 
.A(n_695),
.B(n_556),
.C(n_452),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_614),
.A2(n_609),
.B1(n_602),
.B2(n_458),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_594),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_789),
.B(n_772),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_SL g911 ( 
.A(n_816),
.B(n_745),
.Y(n_911)
);

BUFx8_ASAP7_75t_L g912 ( 
.A(n_768),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_799),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_744),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_878),
.A2(n_886),
.B(n_906),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_802),
.Y(n_916)
);

OAI33xp33_ASAP7_75t_L g917 ( 
.A1(n_750),
.A2(n_748),
.A3(n_759),
.B1(n_747),
.B2(n_767),
.B3(n_765),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_760),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_779),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_809),
.B(n_808),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_906),
.A2(n_881),
.B(n_873),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_827),
.B(n_836),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_772),
.B(n_909),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_L g924 ( 
.A1(n_862),
.A2(n_835),
.B(n_851),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_860),
.B(n_775),
.Y(n_925)
);

O2A1O1Ixp5_ASAP7_75t_L g926 ( 
.A1(n_790),
.A2(n_810),
.B(n_762),
.C(n_901),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_783),
.A2(n_908),
.B1(n_852),
.B2(n_875),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_900),
.A2(n_892),
.B(n_846),
.C(n_887),
.Y(n_928)
);

XOR2xp5_ASAP7_75t_L g929 ( 
.A(n_826),
.B(n_842),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_873),
.A2(n_881),
.B(n_893),
.Y(n_930)
);

CKINVDCx8_ASAP7_75t_R g931 ( 
.A(n_839),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_864),
.B(n_784),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_806),
.B(n_880),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_757),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_864),
.B(n_778),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_760),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_SL g937 ( 
.A1(n_750),
.A2(n_748),
.B1(n_879),
.B2(n_891),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_859),
.A2(n_885),
.B(n_800),
.C(n_876),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_905),
.B(n_807),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_852),
.A2(n_890),
.B1(n_824),
.B2(n_823),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_818),
.B(n_820),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_792),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_903),
.A2(n_830),
.B(n_837),
.C(n_840),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_887),
.A2(n_884),
.B(n_758),
.C(n_903),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_898),
.B(n_749),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_782),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_866),
.B(n_868),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_796),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_847),
.A2(n_899),
.B(n_896),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_847),
.A2(n_831),
.B(n_785),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_822),
.B(n_829),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_758),
.A2(n_907),
.B(n_902),
.C(n_877),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_746),
.B(n_806),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_850),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_L g955 ( 
.A1(n_901),
.A2(n_897),
.B(n_755),
.C(n_871),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_785),
.A2(n_833),
.B(n_849),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_882),
.A2(n_883),
.B(n_838),
.C(n_848),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_823),
.A2(n_824),
.B1(n_834),
.B2(n_863),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_SL g959 ( 
.A1(n_895),
.A2(n_754),
.B1(n_832),
.B2(n_857),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_839),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_867),
.A2(n_811),
.B(n_812),
.C(n_770),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_848),
.A2(n_853),
.B(n_849),
.C(n_791),
.Y(n_962)
);

AND2x6_ASAP7_75t_SL g963 ( 
.A(n_821),
.B(n_793),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_760),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_854),
.B(n_771),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_834),
.A2(n_863),
.B1(n_797),
.B2(n_752),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_853),
.A2(n_888),
.B(n_874),
.C(n_805),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_803),
.A2(n_766),
.B(n_776),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_781),
.B(n_855),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_786),
.B(n_889),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_754),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_786),
.B(n_819),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_894),
.A2(n_756),
.B(n_773),
.C(n_843),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_752),
.A2(n_841),
.B1(n_753),
.B2(n_788),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_894),
.A2(n_843),
.B(n_865),
.C(n_774),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_814),
.B(n_813),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_763),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_777),
.A2(n_872),
.B(n_817),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_764),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_869),
.B(n_825),
.Y(n_980)
);

BUFx4_ASAP7_75t_SL g981 ( 
.A(n_793),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_764),
.B(n_801),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_777),
.A2(n_904),
.B1(n_787),
.B2(n_798),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_764),
.B(n_801),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_801),
.B(n_869),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_815),
.A2(n_751),
.B(n_845),
.C(n_858),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_804),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_804),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_828),
.Y(n_989)
);

OA21x2_ASAP7_75t_L g990 ( 
.A1(n_861),
.A2(n_865),
.B(n_856),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_869),
.B(n_780),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_844),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_769),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_844),
.A2(n_761),
.B1(n_870),
.B2(n_825),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_870),
.A2(n_456),
.B(n_606),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_870),
.B(n_827),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_870),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_816),
.A2(n_852),
.B1(n_862),
.B2(n_836),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_827),
.A2(n_836),
.B(n_783),
.C(n_862),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_906),
.B(n_864),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_827),
.A2(n_862),
.B(n_789),
.C(n_835),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_906),
.B(n_864),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_827),
.A2(n_862),
.B(n_789),
.C(n_835),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_827),
.B(n_457),
.C(n_614),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_816),
.A2(n_852),
.B1(n_827),
.B2(n_786),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_827),
.A2(n_836),
.B(n_783),
.C(n_862),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_906),
.B(n_864),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_827),
.B(n_602),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_781),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_760),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_906),
.B(n_864),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_878),
.A2(n_456),
.B(n_606),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_827),
.B(n_602),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_827),
.B(n_447),
.C(n_386),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_SL g1015 ( 
.A(n_816),
.B(n_457),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_789),
.B(n_457),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_906),
.B(n_864),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_906),
.B(n_864),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_827),
.A2(n_783),
.B1(n_816),
.B2(n_906),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_744),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_827),
.A2(n_862),
.B(n_789),
.C(n_835),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_906),
.B(n_864),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_760),
.Y(n_1023)
);

AO32x1_ASAP7_75t_L g1024 ( 
.A1(n_769),
.A2(n_794),
.A3(n_874),
.B1(n_784),
.B2(n_860),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_809),
.B(n_808),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_760),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_906),
.B(n_864),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_799),
.B(n_416),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_795),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_799),
.B(n_416),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_953),
.B(n_948),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1016),
.B(n_910),
.Y(n_1032)
);

OA21x2_ASAP7_75t_L g1033 ( 
.A1(n_949),
.A2(n_956),
.B(n_955),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_927),
.A2(n_1019),
.B1(n_1014),
.B2(n_922),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1015),
.B(n_1007),
.Y(n_1036)
);

INVx5_ASAP7_75t_L g1037 ( 
.A(n_936),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_999),
.A2(n_1006),
.B(n_1013),
.C(n_1008),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1011),
.B(n_1017),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_914),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_995),
.A2(n_968),
.B(n_950),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_930),
.A2(n_967),
.B(n_962),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_998),
.A2(n_1005),
.B(n_924),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_912),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_SL g1045 ( 
.A1(n_928),
.A2(n_952),
.B(n_957),
.C(n_944),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1001),
.A2(n_1021),
.B(n_1003),
.C(n_924),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_1004),
.A2(n_938),
.B(n_943),
.C(n_933),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_987),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_935),
.B(n_1018),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_915),
.A2(n_996),
.B(n_921),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1022),
.B(n_1027),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_939),
.Y(n_1052)
);

AOI32xp33_ASAP7_75t_L g1053 ( 
.A1(n_911),
.A2(n_976),
.A3(n_978),
.B1(n_937),
.B2(n_940),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_932),
.B(n_941),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1012),
.A2(n_926),
.B(n_997),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_945),
.B(n_925),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_L g1057 ( 
.A1(n_985),
.A2(n_991),
.B(n_917),
.C(n_974),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_975),
.A2(n_961),
.B(n_973),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1020),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_993),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_990),
.A2(n_970),
.B(n_972),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_986),
.A2(n_994),
.B(n_990),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_947),
.B(n_923),
.Y(n_1063)
);

BUFx8_ASAP7_75t_L g1064 ( 
.A(n_946),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_SL g1065 ( 
.A1(n_983),
.A2(n_994),
.B(n_958),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1024),
.A2(n_980),
.B(n_982),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_912),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1024),
.A2(n_984),
.B(n_992),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_951),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_954),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1024),
.A2(n_992),
.B(n_1029),
.Y(n_1071)
);

AOI221x1_ASAP7_75t_L g1072 ( 
.A1(n_978),
.A2(n_959),
.B1(n_965),
.B2(n_942),
.C(n_919),
.Y(n_1072)
);

BUFx10_ASAP7_75t_L g1073 ( 
.A(n_913),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_920),
.B(n_1025),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_934),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_936),
.Y(n_1076)
);

AO31x2_ASAP7_75t_L g1077 ( 
.A1(n_977),
.A2(n_1009),
.A3(n_988),
.B(n_931),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_920),
.A2(n_1025),
.B(n_960),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_988),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_918),
.A2(n_979),
.B(n_1026),
.Y(n_1080)
);

CKINVDCx14_ASAP7_75t_R g1081 ( 
.A(n_1028),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1026),
.A2(n_987),
.B(n_1023),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1030),
.B(n_916),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_987),
.A2(n_969),
.B(n_1023),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_951),
.B(n_1023),
.Y(n_1085)
);

AOI221x1_ASAP7_75t_L g1086 ( 
.A1(n_964),
.A2(n_1010),
.B1(n_963),
.B2(n_981),
.C(n_969),
.Y(n_1086)
);

NAND3x1_ASAP7_75t_L g1087 ( 
.A(n_929),
.B(n_953),
.C(n_971),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_964),
.A2(n_1010),
.B(n_953),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_1010),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_915),
.A2(n_996),
.B(n_456),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_949),
.A2(n_1006),
.B(n_999),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_996),
.B(n_456),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_927),
.A2(n_999),
.A3(n_1006),
.B(n_1019),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1016),
.B(n_1015),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_998),
.A2(n_827),
.B1(n_816),
.B2(n_999),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_914),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_912),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_954),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_936),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_939),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_914),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_998),
.A2(n_827),
.B1(n_816),
.B2(n_999),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_1009),
.B(n_781),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_936),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.C(n_1014),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_912),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_914),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_949),
.A2(n_956),
.B(n_955),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_1014),
.B(n_827),
.C(n_447),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1015),
.B(n_308),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_SL g1119 ( 
.A(n_989),
.B(n_1000),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.C(n_1014),
.Y(n_1120)
);

AO32x2_ASAP7_75t_L g1121 ( 
.A1(n_927),
.A2(n_1019),
.A3(n_852),
.B1(n_940),
.B2(n_750),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.C(n_1014),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_927),
.A2(n_999),
.A3(n_1006),
.B(n_1019),
.Y(n_1123)
);

BUFx10_ASAP7_75t_L g1124 ( 
.A(n_1016),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_927),
.A2(n_999),
.A3(n_1006),
.B(n_1019),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_SL g1127 ( 
.A(n_912),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_998),
.A2(n_816),
.B1(n_852),
.B2(n_924),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1130)
);

AOI211x1_ASAP7_75t_L g1131 ( 
.A1(n_1014),
.A2(n_924),
.B(n_978),
.C(n_927),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_998),
.A2(n_827),
.B1(n_816),
.B2(n_999),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_912),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1014),
.A2(n_862),
.B1(n_1005),
.B2(n_556),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_1000),
.Y(n_1137)
);

INVx5_ASAP7_75t_L g1138 ( 
.A(n_936),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_SL g1139 ( 
.A(n_966),
.B(n_781),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_SL g1140 ( 
.A1(n_998),
.A2(n_852),
.B1(n_937),
.B2(n_924),
.C(n_645),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_999),
.A2(n_827),
.B(n_1006),
.C(n_1014),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_915),
.A2(n_996),
.B(n_456),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_914),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_914),
.Y(n_1145)
);

AO21x1_ASAP7_75t_L g1146 ( 
.A1(n_927),
.A2(n_922),
.B(n_1019),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_914),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_L g1149 ( 
.A1(n_922),
.A2(n_827),
.B(n_1006),
.C(n_999),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_995),
.A2(n_968),
.B(n_949),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1116),
.B(n_1053),
.C(n_1140),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1052),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_SL g1156 ( 
.A1(n_1129),
.A2(n_1128),
.B(n_1096),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1103),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1098),
.B(n_1107),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1059),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1049),
.B(n_1137),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1127),
.B(n_1100),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1114),
.A2(n_1142),
.B(n_1118),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1090),
.A2(n_1092),
.B(n_1143),
.Y(n_1163)
);

INVxp33_ASAP7_75t_L g1164 ( 
.A(n_1032),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1065),
.A2(n_1146),
.B(n_1047),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1046),
.A2(n_1122),
.B(n_1120),
.C(n_1110),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1056),
.B(n_1034),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1113),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1039),
.B(n_1051),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1141),
.A2(n_1132),
.B(n_1135),
.C(n_1134),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1150),
.A2(n_1151),
.B(n_1041),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1094),
.A2(n_1117),
.B1(n_1148),
.B2(n_1106),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1078),
.B(n_1037),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1097),
.B(n_1125),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1131),
.B(n_1043),
.Y(n_1175)
);

OAI222xp33_ASAP7_75t_L g1176 ( 
.A1(n_1121),
.A2(n_1036),
.B1(n_1130),
.B2(n_1152),
.C1(n_1054),
.C2(n_1063),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1048),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1038),
.A2(n_1149),
.B(n_1057),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1035),
.A2(n_1121),
.B1(n_1091),
.B2(n_1081),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1045),
.A2(n_1042),
.B(n_1091),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1042),
.A2(n_1055),
.B(n_1033),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1064),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1066),
.A2(n_1068),
.B(n_1071),
.Y(n_1183)
);

AO21x1_ASAP7_75t_SL g1184 ( 
.A1(n_1060),
.A2(n_1085),
.B(n_1079),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1070),
.B(n_1147),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1037),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1119),
.A2(n_1136),
.B1(n_1035),
.B2(n_1124),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1061),
.A2(n_1033),
.B(n_1115),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1104),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1115),
.A2(n_1084),
.B(n_1060),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1072),
.A2(n_1145),
.B(n_1144),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_SL g1192 ( 
.A1(n_1079),
.A2(n_1145),
.B(n_1075),
.C(n_1121),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1074),
.B(n_1101),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1080),
.A2(n_1082),
.B(n_1088),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1040),
.Y(n_1195)
);

OAI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1069),
.A2(n_1099),
.B1(n_1031),
.B2(n_1083),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1064),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1037),
.B(n_1138),
.Y(n_1198)
);

AO22x2_ASAP7_75t_L g1199 ( 
.A1(n_1093),
.A2(n_1126),
.B1(n_1123),
.B2(n_1086),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1139),
.A2(n_1126),
.B(n_1123),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1108),
.A2(n_1089),
.B(n_1087),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1044),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1073),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1077),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1112),
.A2(n_1067),
.B1(n_1133),
.B2(n_1073),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1076),
.A2(n_998),
.B1(n_816),
.B2(n_626),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1102),
.A2(n_1105),
.B(n_1095),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1102),
.A2(n_1105),
.B(n_1095),
.Y(n_1208)
);

AO221x2_ASAP7_75t_L g1209 ( 
.A1(n_1109),
.A2(n_750),
.B1(n_937),
.B2(n_1136),
.C(n_1107),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1109),
.A2(n_1105),
.B(n_1095),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_L g1211 ( 
.A1(n_1098),
.A2(n_998),
.B1(n_1132),
.B2(n_1107),
.C(n_1140),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1129),
.A2(n_816),
.B1(n_750),
.B2(n_1098),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1037),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1116),
.A2(n_827),
.B(n_1014),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1058),
.A2(n_1050),
.B(n_1062),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1049),
.B(n_1137),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1059),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1117),
.A2(n_623),
.B1(n_669),
.B2(n_383),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1059),
.Y(n_1222)
);

AO21x2_ASAP7_75t_L g1223 ( 
.A1(n_1050),
.A2(n_1092),
.B(n_1090),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1129),
.A2(n_642),
.B(n_626),
.Y(n_1225)
);

AO21x2_ASAP7_75t_L g1226 ( 
.A1(n_1050),
.A2(n_1092),
.B(n_1090),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1129),
.A2(n_816),
.B1(n_750),
.B2(n_1098),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1098),
.A2(n_1132),
.B1(n_1107),
.B2(n_927),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1032),
.B(n_1014),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1231)
);

BUFx2_ASAP7_75t_R g1232 ( 
.A(n_1044),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1032),
.B(n_1049),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1078),
.B(n_781),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1052),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1096),
.A2(n_827),
.B(n_1006),
.C(n_999),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_SL g1238 ( 
.A1(n_1065),
.A2(n_1146),
.B(n_1047),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1037),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1049),
.B(n_1137),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1058),
.A2(n_1050),
.B(n_1062),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1064),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1096),
.A2(n_827),
.B(n_1006),
.C(n_999),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_SL g1244 ( 
.A1(n_1110),
.A2(n_827),
.B(n_1006),
.C(n_999),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1058),
.A2(n_1050),
.B(n_1062),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1058),
.A2(n_1050),
.B(n_1062),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1081),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1058),
.A2(n_1050),
.B(n_1062),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1032),
.B(n_1014),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1095),
.A2(n_1111),
.B(n_1105),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1129),
.A2(n_998),
.B1(n_816),
.B2(n_626),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1170),
.A2(n_1166),
.B(n_1156),
.C(n_1237),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1160),
.B(n_1218),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1240),
.B(n_1172),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1185),
.B(n_1155),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1236),
.B(n_1167),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1169),
.B(n_1174),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1229),
.B(n_1250),
.Y(n_1260)
);

O2A1O1Ixp5_ASAP7_75t_L g1261 ( 
.A1(n_1158),
.A2(n_1215),
.B(n_1176),
.C(n_1237),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1220),
.B(n_1222),
.Y(n_1262)
);

O2A1O1Ixp5_ASAP7_75t_L g1263 ( 
.A1(n_1158),
.A2(n_1176),
.B(n_1243),
.C(n_1178),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1225),
.A2(n_1253),
.B(n_1243),
.C(n_1244),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1229),
.B(n_1250),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1170),
.A2(n_1166),
.B(n_1211),
.C(n_1153),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1175),
.B(n_1209),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1175),
.B(n_1209),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1244),
.A2(n_1180),
.B(n_1226),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1187),
.B(n_1168),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1157),
.B(n_1211),
.Y(n_1271)
);

CKINVDCx11_ASAP7_75t_R g1272 ( 
.A(n_1182),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1206),
.A2(n_1165),
.B(n_1238),
.C(n_1196),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1190),
.A2(n_1200),
.B(n_1171),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1179),
.B(n_1193),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1213),
.B(n_1227),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1200),
.A2(n_1154),
.B(n_1251),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1223),
.A2(n_1163),
.B(n_1228),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1198),
.A2(n_1239),
.B(n_1214),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1228),
.B(n_1195),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1182),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1221),
.A2(n_1205),
.B1(n_1173),
.B2(n_1232),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1198),
.A2(n_1214),
.B(n_1239),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1191),
.B(n_1204),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1205),
.A2(n_1232),
.B1(n_1199),
.B2(n_1234),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1162),
.A2(n_1252),
.B(n_1212),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1217),
.A2(n_1230),
.B(n_1247),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1214),
.A2(n_1239),
.B(n_1186),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1242),
.A2(n_1192),
.B(n_1161),
.C(n_1177),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1191),
.B(n_1201),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1183),
.B(n_1194),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1216),
.A2(n_1249),
.B(n_1245),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1202),
.A2(n_1197),
.B1(n_1248),
.B2(n_1203),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1219),
.A2(n_1231),
.B(n_1235),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1241),
.A2(n_1245),
.B1(n_1246),
.B2(n_1210),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1241),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1241),
.B(n_1245),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1246),
.B(n_1207),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1208),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1224),
.B(n_1189),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1155),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1160),
.B(n_1218),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1213),
.A2(n_998),
.B1(n_1227),
.B2(n_816),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1213),
.A2(n_998),
.B1(n_1227),
.B2(n_816),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1160),
.B(n_1218),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1213),
.A2(n_998),
.B1(n_1227),
.B2(n_816),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1213),
.A2(n_998),
.B1(n_1227),
.B2(n_816),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1164),
.B(n_1233),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1160),
.B(n_1218),
.Y(n_1309)
);

AND2x2_ASAP7_75t_SL g1310 ( 
.A(n_1213),
.B(n_816),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1159),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1170),
.A2(n_827),
.B(n_1050),
.Y(n_1312)
);

NOR2x1_ASAP7_75t_SL g1313 ( 
.A(n_1184),
.B(n_1158),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1170),
.A2(n_1166),
.B(n_827),
.C(n_816),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1181),
.A2(n_1188),
.B(n_1180),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1300),
.B(n_1291),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1300),
.B(n_1298),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1290),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1297),
.B(n_1296),
.Y(n_1319)
);

AO21x2_ASAP7_75t_L g1320 ( 
.A1(n_1269),
.A2(n_1292),
.B(n_1278),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1295),
.A2(n_1263),
.B(n_1312),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1284),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1280),
.B(n_1315),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1274),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1277),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1261),
.A2(n_1263),
.B(n_1266),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1299),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1299),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1277),
.B(n_1256),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1258),
.B(n_1257),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1314),
.A2(n_1254),
.B(n_1266),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1311),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1262),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1303),
.A2(n_1304),
.B1(n_1306),
.B2(n_1307),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1286),
.A2(n_1287),
.B(n_1294),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1314),
.A2(n_1254),
.B(n_1273),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1270),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1261),
.B(n_1275),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1287),
.Y(n_1339)
);

AND2x2_ASAP7_75t_SL g1340 ( 
.A(n_1321),
.B(n_1310),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1329),
.B(n_1301),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1316),
.B(n_1313),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1323),
.B(n_1268),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1323),
.B(n_1267),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1323),
.B(n_1265),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1319),
.B(n_1260),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1316),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1318),
.B(n_1305),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1339),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1316),
.B(n_1308),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1329),
.B(n_1255),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1329),
.B(n_1309),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1332),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1316),
.B(n_1317),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1322),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1324),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1331),
.Y(n_1357)
);

OAI211xp5_ASAP7_75t_L g1358 ( 
.A1(n_1326),
.A2(n_1264),
.B(n_1276),
.C(n_1271),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1358),
.A2(n_1334),
.B1(n_1326),
.B2(n_1310),
.Y(n_1359)
);

NOR3xp33_ASAP7_75t_SL g1360 ( 
.A(n_1358),
.B(n_1281),
.C(n_1326),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1355),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1348),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1348),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1348),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_SL g1366 ( 
.A(n_1358),
.B(n_1328),
.C(n_1334),
.Y(n_1366)
);

AOI31xp33_ASAP7_75t_L g1367 ( 
.A1(n_1351),
.A2(n_1328),
.A3(n_1338),
.B(n_1327),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1355),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1347),
.Y(n_1369)
);

NAND4xp25_ASAP7_75t_L g1370 ( 
.A(n_1357),
.B(n_1259),
.C(n_1302),
.D(n_1338),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1340),
.A2(n_1331),
.B1(n_1336),
.B2(n_1338),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1346),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1340),
.A2(n_1331),
.B1(n_1336),
.B2(n_1282),
.Y(n_1373)
);

AOI221xp5_ASAP7_75t_L g1374 ( 
.A1(n_1357),
.A2(n_1331),
.B1(n_1336),
.B2(n_1285),
.C(n_1318),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1350),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1341),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1340),
.A2(n_1328),
.B1(n_1327),
.B2(n_1337),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1340),
.A2(n_1327),
.B1(n_1337),
.B2(n_1330),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1341),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1353),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1340),
.A2(n_1331),
.B1(n_1336),
.B2(n_1337),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1353),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1347),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1347),
.Y(n_1384)
);

AO21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1351),
.A2(n_1329),
.B(n_1333),
.Y(n_1385)
);

OAI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1357),
.A2(n_1330),
.B1(n_1293),
.B2(n_1289),
.C(n_1333),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1354),
.B(n_1317),
.Y(n_1387)
);

INVx4_ASAP7_75t_SL g1388 ( 
.A(n_1375),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1384),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1364),
.B(n_1345),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1367),
.A2(n_1335),
.B(n_1320),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1363),
.B(n_1351),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1361),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1362),
.B(n_1365),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1385),
.B(n_1383),
.Y(n_1395)
);

INVx4_ASAP7_75t_SL g1396 ( 
.A(n_1375),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1361),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1380),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1383),
.Y(n_1399)
);

INVxp67_ASAP7_75t_L g1400 ( 
.A(n_1386),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1368),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1385),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1382),
.A2(n_1356),
.B(n_1349),
.Y(n_1403)
);

OAI31xp33_ASAP7_75t_L g1404 ( 
.A1(n_1359),
.A2(n_1337),
.A3(n_1352),
.B(n_1342),
.Y(n_1404)
);

BUFx8_ASAP7_75t_L g1405 ( 
.A(n_1369),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1374),
.A2(n_1324),
.B(n_1325),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1376),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_SL g1408 ( 
.A(n_1402),
.B(n_1377),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1392),
.B(n_1390),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1392),
.B(n_1363),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1394),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1397),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1388),
.B(n_1396),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1399),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1388),
.B(n_1347),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_SL g1416 ( 
.A(n_1404),
.B(n_1366),
.C(n_1370),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1397),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1400),
.B(n_1345),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1388),
.B(n_1387),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1388),
.B(n_1387),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1388),
.B(n_1354),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1402),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1400),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1399),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1403),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1398),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1407),
.B(n_1272),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1399),
.Y(n_1428)
);

NOR3xp33_ASAP7_75t_L g1429 ( 
.A(n_1389),
.B(n_1357),
.C(n_1378),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1396),
.B(n_1372),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1396),
.B(n_1379),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1404),
.B(n_1343),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1405),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1405),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1398),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1402),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1393),
.B(n_1401),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1406),
.B(n_1343),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1398),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1423),
.B(n_1344),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1428),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_SL g1442 ( 
.A(n_1436),
.B(n_1402),
.Y(n_1442)
);

AOI21xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1427),
.A2(n_1406),
.B(n_1272),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1426),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1428),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1413),
.B(n_1396),
.Y(n_1446)
);

NOR4xp25_ASAP7_75t_L g1447 ( 
.A(n_1411),
.B(n_1424),
.C(n_1422),
.D(n_1417),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1425),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1426),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1413),
.B(n_1396),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1424),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1435),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1435),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1416),
.A2(n_1360),
.B1(n_1373),
.B2(n_1371),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1425),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1418),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_1395),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1409),
.B(n_1401),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1408),
.B(n_1395),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1414),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1419),
.B(n_1395),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1436),
.B(n_1402),
.Y(n_1462)
);

AOI21xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1433),
.A2(n_1434),
.B(n_1429),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1432),
.A2(n_1406),
.B(n_1391),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1436),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1439),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1431),
.A2(n_1422),
.B(n_1430),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1439),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1425),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1431),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1422),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1437),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1471),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1441),
.B(n_1409),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1471),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1444),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1442),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1447),
.B(n_1412),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1462),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1457),
.B(n_1419),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1444),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1441),
.B(n_1410),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1445),
.Y(n_1483)
);

OAI21xp33_ASAP7_75t_L g1484 ( 
.A1(n_1454),
.A2(n_1381),
.B(n_1438),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1410),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1449),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1460),
.B(n_1412),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1457),
.B(n_1420),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1454),
.A2(n_1422),
.B(n_1433),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1417),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1459),
.B(n_1420),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1449),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1452),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1460),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1462),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1452),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1450),
.B(n_1415),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1480),
.B(n_1446),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1473),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1473),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1483),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1494),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1482),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1479),
.B(n_1465),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1480),
.B(n_1488),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1488),
.B(n_1446),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1478),
.A2(n_1459),
.B(n_1465),
.Y(n_1507)
);

AOI332xp33_ASAP7_75t_L g1508 ( 
.A1(n_1486),
.A2(n_1472),
.A3(n_1451),
.B1(n_1453),
.B2(n_1468),
.B3(n_1466),
.C1(n_1450),
.C2(n_1469),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1482),
.Y(n_1509)
);

AOI321xp33_ASAP7_75t_L g1510 ( 
.A1(n_1489),
.A2(n_1484),
.A3(n_1464),
.B1(n_1491),
.B2(n_1443),
.C(n_1497),
.Y(n_1510)
);

NOR2xp67_ASAP7_75t_L g1511 ( 
.A(n_1477),
.B(n_1470),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1491),
.B(n_1450),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1490),
.A2(n_1443),
.B(n_1463),
.C(n_1467),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1479),
.A2(n_1463),
.B(n_1451),
.C(n_1462),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1497),
.A2(n_1434),
.B1(n_1450),
.B2(n_1402),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1499),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1500),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1500),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1514),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1514),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1498),
.A2(n_1497),
.B1(n_1357),
.B2(n_1442),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1503),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1511),
.B(n_1495),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1503),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1513),
.A2(n_1485),
.B1(n_1474),
.B2(n_1402),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1526),
.A2(n_1510),
.B1(n_1515),
.B2(n_1516),
.C(n_1502),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1524),
.A2(n_1507),
.B(n_1518),
.Y(n_1528)
);

OAI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1518),
.A2(n_1508),
.B(n_1507),
.C(n_1501),
.Y(n_1529)
);

NOR3xp33_ASAP7_75t_SL g1530 ( 
.A(n_1517),
.B(n_1501),
.C(n_1504),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1519),
.B(n_1509),
.Y(n_1531)
);

OAI322xp33_ASAP7_75t_L g1532 ( 
.A1(n_1523),
.A2(n_1509),
.A3(n_1487),
.B1(n_1474),
.B2(n_1495),
.C1(n_1493),
.C2(n_1492),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1525),
.A2(n_1505),
.B1(n_1506),
.B2(n_1498),
.C(n_1512),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1520),
.A2(n_1506),
.B(n_1512),
.C(n_1505),
.Y(n_1534)
);

OAI211xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1522),
.A2(n_1475),
.B(n_1487),
.C(n_1485),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1530),
.A2(n_1462),
.B1(n_1402),
.B2(n_1521),
.Y(n_1536)
);

OAI21xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1533),
.A2(n_1461),
.B(n_1472),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1534),
.B(n_1461),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1527),
.A2(n_1529),
.B1(n_1528),
.B2(n_1535),
.C(n_1532),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1531),
.A2(n_1415),
.B1(n_1406),
.B2(n_1481),
.Y(n_1540)
);

NOR2x1_ASAP7_75t_L g1541 ( 
.A(n_1536),
.B(n_1538),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1537),
.B(n_1421),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1539),
.B(n_1476),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1540),
.B(n_1476),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1536),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1539),
.B(n_1481),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_R g1547 ( 
.A(n_1545),
.B(n_1496),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1542),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1543),
.A2(n_1496),
.B1(n_1440),
.B2(n_1458),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1546),
.B(n_1458),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1541),
.Y(n_1551)
);

AND4x2_ASAP7_75t_L g1552 ( 
.A(n_1551),
.B(n_1544),
.C(n_1448),
.D(n_1469),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1548),
.B(n_1415),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1550),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1552),
.Y(n_1555)
);

AO22x2_ASAP7_75t_L g1556 ( 
.A1(n_1555),
.A2(n_1554),
.B1(n_1553),
.B2(n_1549),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1556),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1557),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1558),
.A2(n_1547),
.B1(n_1455),
.B2(n_1469),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1559),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1560),
.A2(n_1455),
.B(n_1448),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1560),
.B(n_1448),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1562),
.B(n_1561),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1562),
.A2(n_1455),
.B(n_1453),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1563),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1565),
.A2(n_1564),
.B1(n_1468),
.B2(n_1466),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_L g1567 ( 
.A1(n_1566),
.A2(n_1288),
.B(n_1279),
.C(n_1283),
.Y(n_1567)
);


endmodule