module real_aes_9025_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g433 ( .A(n_0), .Y(n_433) );
INVx1_ASAP7_75t_L g500 ( .A(n_1), .Y(n_500) );
INVx1_ASAP7_75t_L g249 ( .A(n_2), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_3), .A2(n_38), .B1(n_168), .B2(n_528), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g156 ( .A1(n_4), .A2(n_157), .B(n_158), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_5), .B(n_155), .Y(n_477) );
AND2x6_ASAP7_75t_L g130 ( .A(n_6), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_7), .A2(n_225), .B(n_226), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_8), .B(n_39), .Y(n_434) );
INVx1_ASAP7_75t_L g165 ( .A(n_9), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_10), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g127 ( .A(n_11), .Y(n_127) );
INVx1_ASAP7_75t_L g496 ( .A(n_12), .Y(n_496) );
INVx1_ASAP7_75t_L g231 ( .A(n_13), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_14), .B(n_133), .Y(n_534) );
AOI222xp33_ASAP7_75t_SL g445 ( .A1(n_15), .A2(n_446), .B1(n_447), .B2(n_456), .C1(n_744), .C2(n_745), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_16), .B(n_123), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_17), .A2(n_104), .B1(n_437), .B2(n_444), .C1(n_748), .C2(n_753), .Y(n_103) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_17), .B(n_106), .Y(n_105) );
AO32x2_ASAP7_75t_L g525 ( .A1(n_17), .A2(n_122), .A3(n_155), .B1(n_488), .B2(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_18), .B(n_168), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_19), .B(n_176), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_20), .B(n_123), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_21), .A2(n_50), .B1(n_168), .B2(n_528), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_22), .B(n_157), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_23), .A2(n_77), .B1(n_133), .B2(n_168), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_24), .B(n_168), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_25), .B(n_153), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_26), .A2(n_448), .B1(n_449), .B2(n_455), .Y(n_447) );
INVx1_ASAP7_75t_L g455 ( .A(n_26), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_27), .A2(n_229), .B(n_230), .C(n_232), .Y(n_228) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_28), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_29), .B(n_170), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_30), .B(n_163), .Y(n_250) );
INVx1_ASAP7_75t_L g141 ( .A(n_31), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_32), .B(n_170), .Y(n_522) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_34), .B(n_168), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_35), .B(n_170), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_36), .A2(n_42), .B1(n_111), .B2(n_112), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_36), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_37), .A2(n_130), .B(n_142), .C(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g139 ( .A(n_40), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_41), .B(n_163), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_42), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_43), .B(n_168), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_44), .A2(n_87), .B1(n_193), .B2(n_528), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_45), .B(n_168), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_46), .B(n_168), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_47), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_48), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_49), .B(n_157), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_51), .A2(n_60), .B1(n_133), .B2(n_168), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_52), .A2(n_133), .B1(n_136), .B2(n_142), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_53), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_54), .B(n_168), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_55), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_56), .B(n_168), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_57), .A2(n_162), .B(n_164), .C(n_167), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_58), .Y(n_206) );
INVx1_ASAP7_75t_L g159 ( .A(n_59), .Y(n_159) );
INVx1_ASAP7_75t_L g131 ( .A(n_61), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_62), .B(n_168), .Y(n_501) );
INVx1_ASAP7_75t_L g126 ( .A(n_63), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_64), .Y(n_440) );
AO32x2_ASAP7_75t_L g545 ( .A1(n_65), .A2(n_155), .A3(n_211), .B1(n_488), .B2(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g485 ( .A(n_66), .Y(n_485) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_67), .A2(n_109), .B1(n_110), .B2(n_113), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_67), .Y(n_113) );
INVx1_ASAP7_75t_L g517 ( .A(n_68), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_69), .A2(n_167), .B(n_176), .C(n_177), .Y(n_175) );
INVxp67_ASAP7_75t_L g178 ( .A(n_70), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_71), .B(n_133), .Y(n_518) );
INVx1_ASAP7_75t_L g443 ( .A(n_72), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_73), .Y(n_150) );
INVx1_ASAP7_75t_L g199 ( .A(n_74), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_75), .A2(n_101), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_75), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_76), .B(n_436), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_78), .A2(n_130), .B(n_142), .C(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_79), .B(n_528), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_80), .B(n_133), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_81), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_83), .B(n_176), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_84), .B(n_133), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_85), .A2(n_130), .B(n_142), .C(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g430 ( .A(n_86), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g459 ( .A(n_86), .B(n_432), .Y(n_459) );
INVx2_ASAP7_75t_L g743 ( .A(n_86), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_88), .A2(n_102), .B1(n_133), .B2(n_134), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_89), .B(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_90), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_91), .A2(n_130), .B(n_142), .C(n_214), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_92), .Y(n_221) );
INVx1_ASAP7_75t_L g174 ( .A(n_93), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_94), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_95), .B(n_189), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_96), .A2(n_450), .B1(n_451), .B2(n_452), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_96), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_97), .B(n_133), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_98), .B(n_155), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_99), .A2(n_157), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_100), .B(n_443), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_101), .Y(n_454) );
OAI21x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_427), .B(n_435), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_108), .B1(n_114), .B2(n_115), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_114), .A2(n_457), .B1(n_460), .B2(n_740), .Y(n_456) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_115), .A2(n_457), .B1(n_746), .B2(n_747), .Y(n_745) );
AND3x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_352), .C(n_401), .Y(n_115) );
NOR3xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_259), .C(n_297), .Y(n_116) );
OAI222xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_180), .B1(n_234), .B2(n_240), .C1(n_254), .C2(n_257), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_151), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_119), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_119), .B(n_302), .Y(n_393) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g270 ( .A(n_120), .B(n_171), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_120), .B(n_152), .Y(n_278) );
AND2x2_ASAP7_75t_L g313 ( .A(n_120), .B(n_290), .Y(n_313) );
OR2x2_ASAP7_75t_L g337 ( .A(n_120), .B(n_152), .Y(n_337) );
OR2x2_ASAP7_75t_L g345 ( .A(n_120), .B(n_244), .Y(n_345) );
AND2x2_ASAP7_75t_L g348 ( .A(n_120), .B(n_171), .Y(n_348) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g242 ( .A(n_121), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g256 ( .A(n_121), .B(n_171), .Y(n_256) );
AND2x2_ASAP7_75t_L g306 ( .A(n_121), .B(n_244), .Y(n_306) );
AND2x2_ASAP7_75t_L g319 ( .A(n_121), .B(n_152), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_121), .B(n_405), .Y(n_426) );
AO21x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_128), .B(n_149), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_122), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g194 ( .A(n_122), .Y(n_194) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_122), .A2(n_245), .B(n_252), .Y(n_244) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_124), .B(n_125), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI22xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B1(n_145), .B2(n_146), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_129), .A2(n_159), .B(n_160), .C(n_161), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_129), .A2(n_160), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_129), .A2(n_160), .B(n_227), .C(n_228), .Y(n_226) );
INVx4_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_130), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g157 ( .A(n_130), .B(n_147), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_130), .A2(n_469), .B(n_472), .Y(n_468) );
BUFx3_ASAP7_75t_L g488 ( .A(n_130), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_130), .A2(n_495), .B(n_499), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_130), .A2(n_516), .B(n_519), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_130), .A2(n_532), .B(n_536), .Y(n_531) );
INVx2_ASAP7_75t_L g251 ( .A(n_133), .Y(n_251) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_139), .B1(n_140), .B2(n_141), .Y(n_136) );
INVx2_ASAP7_75t_L g140 ( .A(n_137), .Y(n_140) );
INVx4_ASAP7_75t_L g229 ( .A(n_137), .Y(n_229) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
AND2x2_ASAP7_75t_L g147 ( .A(n_138), .B(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_138), .Y(n_163) );
INVx3_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
INVx1_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
INVx5_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
BUFx3_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx1_ASAP7_75t_L g528 ( .A(n_143), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_146), .A2(n_199), .B(n_200), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_146), .A2(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g475 ( .A(n_148), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_151), .A2(n_345), .B(n_346), .C(n_349), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_151), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_151), .B(n_289), .Y(n_411) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_171), .Y(n_151) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_152), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g269 ( .A(n_152), .Y(n_269) );
AND2x2_ASAP7_75t_L g296 ( .A(n_152), .B(n_290), .Y(n_296) );
INVx1_ASAP7_75t_SL g304 ( .A(n_152), .Y(n_304) );
AND2x2_ASAP7_75t_L g327 ( .A(n_152), .B(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g405 ( .A(n_152), .Y(n_405) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_169), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_SL g195 ( .A(n_154), .B(n_196), .Y(n_195) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_154), .B(n_488), .C(n_507), .Y(n_506) );
AO21x1_ASAP7_75t_L g551 ( .A1(n_154), .A2(n_507), .B(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_155), .A2(n_172), .B(n_179), .Y(n_171) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_155), .A2(n_468), .B(n_477), .Y(n_467) );
BUFx2_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g484 ( .A1(n_162), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_162), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g217 ( .A(n_163), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_163), .A2(n_476), .B1(n_508), .B2(n_509), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_163), .A2(n_476), .B1(n_527), .B2(n_529), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g546 ( .A1(n_163), .A2(n_166), .B1(n_547), .B2(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_166), .B(n_178), .Y(n_177) );
INVx5_ASAP7_75t_L g189 ( .A(n_166), .Y(n_189) );
O2A1O1Ixp5_ASAP7_75t_SL g516 ( .A1(n_167), .A2(n_189), .B(n_517), .C(n_518), .Y(n_516) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVx1_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
INVx2_ASAP7_75t_L g211 ( .A(n_170), .Y(n_211) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_170), .A2(n_224), .B(n_233), .Y(n_223) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_170), .A2(n_515), .B(n_522), .Y(n_514) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_170), .A2(n_531), .B(n_539), .Y(n_530) );
BUFx2_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
INVx1_ASAP7_75t_L g303 ( .A(n_171), .Y(n_303) );
INVx3_ASAP7_75t_L g328 ( .A(n_171), .Y(n_328) );
INVx1_ASAP7_75t_L g535 ( .A(n_176), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_180), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_208), .Y(n_180) );
INVx1_ASAP7_75t_L g324 ( .A(n_181), .Y(n_324) );
OAI32xp33_ASAP7_75t_L g330 ( .A1(n_181), .A2(n_269), .A3(n_331), .B1(n_332), .B2(n_333), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_181), .A2(n_335), .B1(n_338), .B2(n_343), .Y(n_334) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g272 ( .A(n_182), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g350 ( .A(n_182), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g420 ( .A(n_182), .B(n_366), .Y(n_420) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_197), .Y(n_182) );
AND2x2_ASAP7_75t_L g235 ( .A(n_183), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g265 ( .A(n_183), .Y(n_265) );
INVx1_ASAP7_75t_L g284 ( .A(n_183), .Y(n_284) );
OR2x2_ASAP7_75t_L g292 ( .A(n_183), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g299 ( .A(n_183), .B(n_273), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_183), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g320 ( .A(n_183), .B(n_238), .Y(n_320) );
INVx3_ASAP7_75t_L g342 ( .A(n_183), .Y(n_342) );
AND2x2_ASAP7_75t_L g367 ( .A(n_183), .B(n_239), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_183), .B(n_332), .Y(n_415) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_195), .Y(n_183) );
AOI21xp5_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_186), .B(n_194), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B(n_191), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_189), .A2(n_249), .B(n_250), .C(n_251), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_189), .A2(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g476 ( .A(n_189), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_189), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_191), .A2(n_202), .B(n_203), .Y(n_201) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
INVx1_ASAP7_75t_L g204 ( .A(n_194), .Y(n_204) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_194), .A2(n_480), .B(n_489), .Y(n_479) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_194), .A2(n_494), .B(n_502), .Y(n_493) );
INVx2_ASAP7_75t_L g239 ( .A(n_197), .Y(n_239) );
AND2x2_ASAP7_75t_L g371 ( .A(n_197), .B(n_209), .Y(n_371) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_204), .B(n_205), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_207), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_207), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g413 ( .A(n_208), .Y(n_413) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_222), .Y(n_208) );
INVx1_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_209), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_209), .B(n_239), .Y(n_293) );
AND2x2_ASAP7_75t_L g351 ( .A(n_209), .B(n_274), .Y(n_351) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g237 ( .A(n_210), .Y(n_237) );
AND2x2_ASAP7_75t_L g264 ( .A(n_210), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g273 ( .A(n_210), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_210), .B(n_239), .Y(n_339) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_219), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_218), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_222), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g286 ( .A(n_222), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_222), .B(n_239), .Y(n_332) );
AND2x2_ASAP7_75t_L g341 ( .A(n_222), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g366 ( .A(n_222), .Y(n_366) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g238 ( .A(n_223), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g274 ( .A(n_223), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_229), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g498 ( .A(n_229), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_229), .A2(n_520), .B(n_521), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_234), .A2(n_244), .B1(n_403), .B2(n_406), .Y(n_402) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_236), .A2(n_347), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_237), .B(n_342), .Y(n_359) );
INVx1_ASAP7_75t_L g384 ( .A(n_237), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_238), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g311 ( .A(n_238), .B(n_264), .Y(n_311) );
INVx2_ASAP7_75t_L g267 ( .A(n_239), .Y(n_267) );
INVx1_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_240), .A2(n_392), .B1(n_409), .B2(n_412), .C(n_414), .Y(n_408) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g279 ( .A(n_241), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_241), .B(n_290), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_242), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g333 ( .A(n_242), .B(n_279), .Y(n_333) );
INVx3_ASAP7_75t_SL g374 ( .A(n_242), .Y(n_374) );
AND2x2_ASAP7_75t_L g318 ( .A(n_243), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g347 ( .A(n_243), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_243), .B(n_256), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_243), .B(n_302), .Y(n_388) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_244), .A2(n_316), .A3(n_338), .B1(n_386), .B2(n_388), .C1(n_389), .C2(n_390), .Y(n_385) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_251), .A2(n_496), .B(n_497), .C(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_255), .A2(n_258), .B(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_SL g335 ( .A(n_256), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g357 ( .A(n_256), .B(n_269), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_256), .B(n_296), .Y(n_372) );
INVxp67_ASAP7_75t_L g323 ( .A(n_258), .Y(n_323) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_258), .A2(n_330), .B(n_334), .C(n_344), .Y(n_329) );
OAI221xp5_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_268), .B1(n_271), .B2(n_275), .C(n_280), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g283 ( .A(n_267), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g400 ( .A(n_267), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_268), .A2(n_417), .B1(n_422), .B2(n_423), .C(n_425), .Y(n_416) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_269), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g316 ( .A(n_269), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_269), .B(n_347), .Y(n_354) );
AND2x2_ASAP7_75t_L g396 ( .A(n_269), .B(n_374), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_270), .B(n_295), .Y(n_294) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_270), .A2(n_282), .B1(n_392), .B2(n_393), .Y(n_391) );
OR2x2_ASAP7_75t_L g422 ( .A(n_270), .B(n_290), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g399 ( .A(n_273), .Y(n_399) );
AND2x2_ASAP7_75t_L g424 ( .A(n_273), .B(n_367), .Y(n_424) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_SL g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g288 ( .A(n_278), .B(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_287), .B1(n_291), .B2(n_294), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g355 ( .A(n_283), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_283), .B(n_323), .Y(n_390) );
AOI322xp5_ASAP7_75t_L g314 ( .A1(n_285), .A2(n_315), .A3(n_317), .B1(n_318), .B2(n_320), .C1(n_321), .C2(n_325), .Y(n_314) );
INVxp67_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_288), .A2(n_293), .B1(n_310), .B2(n_312), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_289), .B(n_302), .Y(n_389) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_290), .B(n_328), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_290), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g386 ( .A(n_292), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND3xp33_ASAP7_75t_SL g297 ( .A(n_298), .B(n_314), .C(n_329), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_305), .B2(n_307), .C(n_309), .Y(n_298) );
AND2x2_ASAP7_75t_L g305 ( .A(n_301), .B(n_306), .Y(n_305) );
INVx3_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g315 ( .A(n_306), .B(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_308), .Y(n_387) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_313), .B(n_327), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_316), .B(n_374), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_317), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g392 ( .A(n_320), .Y(n_392) );
AND2x2_ASAP7_75t_L g407 ( .A(n_320), .B(n_384), .Y(n_407) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI211xp5_ASAP7_75t_L g401 ( .A1(n_331), .A2(n_402), .B(n_408), .C(n_416), .Y(n_401) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g370 ( .A(n_341), .B(n_371), .Y(n_370) );
NAND2x1_ASAP7_75t_SL g412 ( .A(n_342), .B(n_413), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g382 ( .A(n_345), .Y(n_382) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
AND2x2_ASAP7_75t_L g381 ( .A(n_351), .B(n_367), .Y(n_381) );
NOR5xp2_ASAP7_75t_L g352 ( .A(n_353), .B(n_368), .C(n_385), .D(n_391), .E(n_394), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_356), .B2(n_358), .C(n_360), .Y(n_353) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_357), .B(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g383 ( .A(n_367), .B(n_384), .Y(n_383) );
OAI221xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_372), .B1(n_373), .B2(n_375), .C(n_378), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_382), .B2(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
AOI211xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_397), .B(n_399), .C(n_400), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
CKINVDCx14_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g436 ( .A(n_430), .Y(n_436) );
INVx1_ASAP7_75t_SL g752 ( .A(n_430), .Y(n_752) );
BUFx2_ASAP7_75t_L g755 ( .A(n_430), .Y(n_755) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_431), .B(n_743), .Y(n_744) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g742 ( .A(n_432), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g750 ( .A(n_440), .B(n_442), .Y(n_750) );
OA21x2_ASAP7_75t_L g754 ( .A1(n_440), .A2(n_441), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g746 ( .A(n_460), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_664), .Y(n_460) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_462), .B(n_622), .Y(n_461) );
NOR4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_562), .C(n_598), .D(n_612), .Y(n_462) );
OAI221xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_510), .B1(n_540), .B2(n_549), .C(n_553), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_464), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_490), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_478), .Y(n_466) );
AND2x2_ASAP7_75t_L g559 ( .A(n_467), .B(n_479), .Y(n_559) );
INVx3_ASAP7_75t_L g567 ( .A(n_467), .Y(n_567) );
AND2x2_ASAP7_75t_L g621 ( .A(n_467), .B(n_493), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_467), .B(n_492), .Y(n_657) );
AND2x2_ASAP7_75t_L g715 ( .A(n_467), .B(n_577), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g486 ( .A(n_475), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_476), .A2(n_486), .B(n_500), .C(n_501), .Y(n_499) );
AND2x2_ASAP7_75t_L g550 ( .A(n_478), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g564 ( .A(n_478), .B(n_493), .Y(n_564) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_479), .B(n_493), .Y(n_579) );
AND2x2_ASAP7_75t_L g591 ( .A(n_479), .B(n_567), .Y(n_591) );
OR2x2_ASAP7_75t_L g593 ( .A(n_479), .B(n_551), .Y(n_593) );
AND2x2_ASAP7_75t_L g628 ( .A(n_479), .B(n_551), .Y(n_628) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_479), .Y(n_673) );
INVx1_ASAP7_75t_L g681 ( .A(n_479), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B(n_488), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_490), .A2(n_599), .B1(n_603), .B2(n_607), .C(n_608), .Y(n_598) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
INVx2_ASAP7_75t_L g557 ( .A(n_492), .Y(n_557) );
AND2x2_ASAP7_75t_L g610 ( .A(n_492), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g629 ( .A(n_492), .B(n_567), .Y(n_629) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g692 ( .A(n_493), .B(n_567), .Y(n_692) );
AND2x2_ASAP7_75t_L g614 ( .A(n_503), .B(n_559), .Y(n_614) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_503), .A2(n_638), .A3(n_683), .B1(n_685), .B2(n_688), .C1(n_690), .C2(n_694), .Y(n_682) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_504), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
AND2x2_ASAP7_75t_L g687 ( .A(n_504), .B(n_567), .Y(n_687) );
AND2x2_ASAP7_75t_L g719 ( .A(n_504), .B(n_591), .Y(n_719) );
OR2x2_ASAP7_75t_L g722 ( .A(n_504), .B(n_723), .Y(n_722) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g552 ( .A(n_505), .Y(n_552) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
INVx1_ASAP7_75t_L g735 ( .A(n_512), .Y(n_735) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g542 ( .A(n_513), .B(n_530), .Y(n_542) );
INVx2_ASAP7_75t_L g575 ( .A(n_513), .Y(n_575) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g597 ( .A(n_514), .Y(n_597) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_514), .Y(n_605) );
OR2x2_ASAP7_75t_L g729 ( .A(n_514), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g554 ( .A(n_523), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g594 ( .A(n_523), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g646 ( .A(n_523), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_530), .Y(n_523) );
AND2x2_ASAP7_75t_L g543 ( .A(n_524), .B(n_544), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g601 ( .A(n_524), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g655 ( .A(n_524), .B(n_545), .Y(n_655) );
OR2x2_ASAP7_75t_L g663 ( .A(n_524), .B(n_597), .Y(n_663) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g572 ( .A(n_525), .Y(n_572) );
AND2x2_ASAP7_75t_L g582 ( .A(n_525), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g606 ( .A(n_525), .B(n_530), .Y(n_606) );
AND2x2_ASAP7_75t_L g670 ( .A(n_525), .B(n_545), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_530), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_530), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
INVx1_ASAP7_75t_L g588 ( .A(n_530), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_530), .Y(n_678) );
INVx1_ASAP7_75t_L g730 ( .A(n_530), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x2_ASAP7_75t_L g707 ( .A(n_541), .B(n_616), .Y(n_707) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g634 ( .A(n_543), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g733 ( .A(n_543), .B(n_668), .Y(n_733) );
INVx1_ASAP7_75t_L g555 ( .A(n_544), .Y(n_555) );
AND2x2_ASAP7_75t_L g581 ( .A(n_544), .B(n_575), .Y(n_581) );
BUFx2_ASAP7_75t_L g640 ( .A(n_544), .Y(n_640) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_545), .Y(n_561) );
INVx1_ASAP7_75t_L g571 ( .A(n_545), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g709 ( .A(n_549), .B(n_556), .Y(n_709) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI32xp33_ASAP7_75t_L g553 ( .A1(n_550), .A2(n_554), .A3(n_556), .B1(n_558), .B2(n_560), .Y(n_553) );
AND2x2_ASAP7_75t_L g693 ( .A(n_550), .B(n_566), .Y(n_693) );
AND2x2_ASAP7_75t_L g731 ( .A(n_550), .B(n_629), .Y(n_731) );
INVx1_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_555), .B(n_617), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_556), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_556), .B(n_559), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_556), .B(n_628), .Y(n_710) );
OR2x2_ASAP7_75t_L g724 ( .A(n_556), .B(n_593), .Y(n_724) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g651 ( .A(n_557), .B(n_559), .Y(n_651) );
OR2x2_ASAP7_75t_L g660 ( .A(n_557), .B(n_647), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_559), .B(n_610), .Y(n_632) );
INVx2_ASAP7_75t_L g647 ( .A(n_561), .Y(n_647) );
OR2x2_ASAP7_75t_L g662 ( .A(n_561), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g677 ( .A(n_561), .B(n_678), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_561), .A2(n_654), .B(n_735), .C(n_736), .Y(n_734) );
OAI321xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_568), .A3(n_573), .B1(n_576), .B2(n_580), .C(n_584), .Y(n_562) );
INVx1_ASAP7_75t_L g675 ( .A(n_563), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g686 ( .A(n_564), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g638 ( .A(n_566), .Y(n_638) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_567), .B(n_681), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_568), .A2(n_706), .B1(n_708), .B2(n_710), .C(n_711), .Y(n_705) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g643 ( .A(n_570), .B(n_617), .Y(n_643) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_571), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g616 ( .A(n_572), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_573), .A2(n_614), .B(n_659), .C(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g625 ( .A(n_575), .B(n_582), .Y(n_625) );
BUFx2_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
INVx1_ASAP7_75t_L g650 ( .A(n_575), .Y(n_650) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OR2x2_ASAP7_75t_L g656 ( .A(n_578), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g739 ( .A(n_578), .Y(n_739) );
INVx1_ASAP7_75t_L g732 ( .A(n_579), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g585 ( .A(n_581), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g689 ( .A(n_581), .B(n_606), .Y(n_689) );
INVx1_ASAP7_75t_L g618 ( .A(n_582), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B1(n_592), .B2(n_594), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_586), .B(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g654 ( .A(n_587), .B(n_655), .Y(n_654) );
BUFx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_588), .B(n_597), .Y(n_617) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g609 ( .A(n_591), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g619 ( .A(n_593), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_596), .A2(n_714), .B1(n_716), .B2(n_717), .C(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g602 ( .A(n_597), .Y(n_602) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_597), .Y(n_668) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_600), .B(n_719), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_601), .A2(n_606), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_604), .B(n_614), .Y(n_711) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g680 ( .A(n_605), .Y(n_680) );
AND2x2_ASAP7_75t_L g639 ( .A(n_606), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g728 ( .A(n_606), .Y(n_728) );
INVx1_ASAP7_75t_L g644 ( .A(n_609), .Y(n_644) );
INVx1_ASAP7_75t_L g699 ( .A(n_610), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B1(n_618), .B2(n_619), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_616), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g684 ( .A(n_617), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_617), .B(n_655), .Y(n_721) );
OR2x2_ASAP7_75t_L g694 ( .A(n_618), .B(n_647), .Y(n_694) );
INVx1_ASAP7_75t_L g633 ( .A(n_619), .Y(n_633) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_621), .B(n_672), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_641), .C(n_652), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_630), .C(n_636), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_625), .A2(n_696), .B1(n_700), .B2(n_703), .C(n_705), .Y(n_695) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g637 ( .A(n_628), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g691 ( .A(n_628), .B(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_629), .A2(n_677), .B(n_679), .C(n_681), .Y(n_676) );
INVx2_ASAP7_75t_L g723 ( .A(n_629), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_633), .B(n_634), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g702 ( .A(n_635), .B(n_655), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_644), .B(n_645), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B(n_651), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_646), .B(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_651), .B(n_738), .Y(n_737) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B(n_658), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g679 ( .A(n_655), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND4x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_695), .C(n_712), .D(n_734), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_682), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_671), .B(n_674), .C(n_676), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_670), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_681), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g716 ( .A(n_691), .Y(n_716) );
INVx2_ASAP7_75t_SL g704 ( .A(n_692), .Y(n_704) );
OR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g717 ( .A(n_702), .Y(n_717) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_720), .Y(n_712) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
OAI221xp5_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_722), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g747 ( .A(n_741), .Y(n_747) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
NAND2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
endmodule