module fake_jpeg_6582_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_35),
.B1(n_23),
.B2(n_25),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_35),
.B1(n_23),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_56),
.B1(n_74),
.B2(n_23),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_35),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_69),
.B(n_26),
.C(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_35),
.B1(n_48),
.B2(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_92),
.B1(n_94),
.B2(n_100),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_17),
.Y(n_128)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_86),
.B1(n_99),
.B2(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_40),
.B1(n_39),
.B2(n_47),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_98),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_47),
.B1(n_41),
.B2(n_29),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_66),
.B1(n_62),
.B2(n_65),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_65),
.B1(n_64),
.B2(n_55),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_128),
.B(n_21),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_112),
.B1(n_76),
.B2(n_78),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_82),
.B1(n_68),
.B2(n_73),
.Y(n_130)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_58),
.B1(n_71),
.B2(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_116),
.B1(n_121),
.B2(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_119),
.Y(n_141)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_118),
.B(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_58),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_89),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_28),
.C(n_19),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_136),
.B1(n_143),
.B2(n_147),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_139),
.B1(n_150),
.B2(n_109),
.Y(n_161)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_106),
.B1(n_113),
.B2(n_116),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_98),
.C(n_19),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_149),
.C(n_125),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_67),
.B1(n_81),
.B2(n_90),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_55),
.B1(n_81),
.B2(n_17),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_49),
.B1(n_96),
.B2(n_90),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_19),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_19),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_153),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_96),
.B1(n_87),
.B2(n_41),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_19),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_30),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_120),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_105),
.B(n_108),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_87),
.B1(n_84),
.B2(n_18),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_102),
.A2(n_84),
.B1(n_18),
.B2(n_22),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_154),
.B1(n_121),
.B2(n_122),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_97),
.C(n_77),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_22),
.B1(n_77),
.B2(n_21),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_156),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_128),
.B(n_126),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_163),
.B(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_162),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_165),
.B1(n_31),
.B2(n_29),
.Y(n_206)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_106),
.B1(n_111),
.B2(n_108),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_185),
.C(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_139),
.B1(n_137),
.B2(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_19),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_19),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_115),
.B(n_110),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_181),
.B(n_31),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

OAI21x1_ASAP7_75t_R g205 ( 
.A1(n_180),
.A2(n_151),
.B(n_31),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_30),
.B(n_24),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_182),
.B(n_145),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_0),
.Y(n_183)
);

AO22x1_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_30),
.B1(n_24),
.B2(n_29),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_143),
.B1(n_130),
.B2(n_136),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_115),
.C(n_30),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_188),
.B(n_197),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_134),
.B(n_152),
.C(n_146),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_173),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_134),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_204),
.C(n_185),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_153),
.B1(n_146),
.B2(n_133),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_170),
.A2(n_151),
.B1(n_24),
.B2(n_29),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_151),
.C(n_24),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_206),
.B1(n_164),
.B2(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_31),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_211),
.B1(n_161),
.B2(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_177),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_184),
.B(n_176),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_15),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_191),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_196),
.B(n_194),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_166),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_163),
.B(n_181),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_210),
.B(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_182),
.B1(n_179),
.B2(n_158),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_235),
.B1(n_200),
.B2(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_227),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_232),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_234),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_175),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_237),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_166),
.C(n_186),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_240),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_167),
.B1(n_172),
.B2(n_4),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_0),
.C(n_3),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_15),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_247),
.B1(n_218),
.B2(n_226),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_259),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_208),
.B1(n_193),
.B2(n_196),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_202),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_202),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_265),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_190),
.C(n_212),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_232),
.C(n_229),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_189),
.B(n_211),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_235),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_189),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_239),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_250),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_221),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_280),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_278),
.B1(n_264),
.B2(n_258),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_244),
.C(n_238),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.C(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_226),
.B1(n_236),
.B2(n_225),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_231),
.C(n_237),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_241),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_228),
.C(n_240),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_263),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_14),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.C(n_265),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_3),
.C(n_4),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_245),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_298),
.B(n_299),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_242),
.B1(n_261),
.B2(n_251),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_249),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_295),
.C(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_260),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_262),
.C(n_247),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_285),
.A2(n_279),
.B1(n_287),
.B2(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_313),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_257),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_305),
.B(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_267),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_271),
.A3(n_281),
.B1(n_267),
.B2(n_280),
.C(n_14),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_5),
.B(n_7),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_289),
.C(n_293),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_12),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_12),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_302),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_289),
.C(n_293),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_324),
.B(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

AOI21x1_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_4),
.B(n_5),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_7),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_314),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_5),
.C(n_7),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_327),
.B(n_329),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_306),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_331),
.B(n_332),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_304),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_315),
.B(n_320),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_333),
.A2(n_336),
.B(n_328),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_316),
.B(n_9),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_339),
.B(n_337),
.Y(n_340)
);

A2O1A1O1Ixp25_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_8),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_335),
.C(n_10),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_11),
.Y(n_342)
);

OAI321xp33_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_334),
.C(n_337),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.Y(n_344)
);


endmodule