module fake_jpeg_2576_n_681 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_681);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_681;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_59),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_60),
.Y(n_197)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g156 ( 
.A(n_61),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_21),
.B(n_9),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_62),
.B(n_72),
.Y(n_141)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_64),
.B(n_66),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_61),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_67),
.B(n_70),
.Y(n_158)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_9),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_21),
.B(n_9),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_74),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_82),
.Y(n_179)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_85),
.B(n_95),
.Y(n_187)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_88),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx16f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_101),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_97),
.Y(n_216)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_7),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_32),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_102),
.B(n_107),
.Y(n_172)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_7),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_104),
.B(n_127),
.Y(n_217)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_26),
.B(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_110),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_32),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_46),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_122),
.B(n_131),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_43),
.Y(n_126)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

HAxp5_ASAP7_75t_SL g127 ( 
.A(n_48),
.B(n_0),
.CON(n_127),
.SN(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_26),
.B(n_10),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_142),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_59),
.A2(n_44),
.B1(n_31),
.B2(n_55),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_144),
.A2(n_159),
.B1(n_165),
.B2(n_167),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_55),
.B1(n_44),
.B2(n_31),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_147),
.A2(n_168),
.B1(n_175),
.B2(n_176),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_70),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_154),
.A2(n_182),
.B1(n_209),
.B2(n_230),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_61),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_157),
.B(n_173),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_59),
.A2(n_44),
.B1(n_31),
.B2(n_55),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_67),
.A2(n_55),
.B1(n_30),
.B2(n_33),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_104),
.A2(n_33),
.B1(n_35),
.B2(n_52),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_99),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_25),
.B1(n_27),
.B2(n_38),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_174),
.A2(n_185),
.B1(n_196),
.B2(n_204),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_69),
.A2(n_35),
.B1(n_36),
.B2(n_52),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_93),
.A2(n_36),
.B1(n_41),
.B2(n_25),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_68),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_130),
.A2(n_27),
.B1(n_39),
.B2(n_45),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_214),
.B1(n_227),
.B2(n_231),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_77),
.A2(n_53),
.B1(n_29),
.B2(n_48),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_90),
.B(n_29),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_83),
.B(n_29),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_79),
.A2(n_53),
.B1(n_48),
.B2(n_58),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_71),
.A2(n_53),
.B1(n_48),
.B2(n_56),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_207),
.A2(n_213),
.B1(n_220),
.B2(n_223),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_73),
.A2(n_75),
.B1(n_128),
.B2(n_124),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_86),
.B(n_10),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_74),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_87),
.A2(n_56),
.B1(n_11),
.B2(n_12),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_78),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_218),
.B(n_229),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_91),
.A2(n_6),
.B1(n_17),
.B2(n_16),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_127),
.A2(n_18),
.B1(n_16),
.B2(n_13),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_18),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_0),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_96),
.A2(n_6),
.B1(n_16),
.B2(n_13),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_80),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_98),
.A2(n_18),
.B1(n_11),
.B2(n_6),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_111),
.Y(n_232)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_233),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_142),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_237),
.B(n_277),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_238),
.A2(n_248),
.B1(n_286),
.B2(n_305),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_239),
.B(n_254),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_89),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_240),
.Y(n_320)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_242),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_141),
.B(n_89),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_244),
.B(n_256),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_147),
.A2(n_123),
.B1(n_119),
.B2(n_114),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_247),
.A2(n_316),
.B1(n_318),
.B2(n_143),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_112),
.B1(n_97),
.B2(n_82),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_249),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_135),
.Y(n_250)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_250),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_251),
.Y(n_321)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_252),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_197),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_253),
.B(n_265),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_151),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_121),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_255),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_141),
.B(n_121),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_133),
.B(n_92),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_257),
.B(n_276),
.Y(n_348)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_258),
.Y(n_371)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_164),
.Y(n_261)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_76),
.B(n_118),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_263),
.A2(n_220),
.B(n_196),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_152),
.Y(n_264)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_264),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_158),
.A2(n_88),
.B(n_113),
.C(n_103),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_150),
.Y(n_266)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_267),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_268),
.Y(n_353)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_269),
.Y(n_356)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_270),
.Y(n_340)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_156),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_274),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_140),
.Y(n_275)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_200),
.B(n_6),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_137),
.B(n_81),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_174),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_283),
.Y(n_326)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_140),
.Y(n_280)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_280),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_149),
.A2(n_88),
.B1(n_11),
.B2(n_4),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_281),
.A2(n_295),
.B1(n_296),
.B2(n_237),
.Y(n_377)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_156),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_172),
.B(n_11),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_284),
.B(n_288),
.Y(n_351)
);

INVx2_ASAP7_75t_R g285 ( 
.A(n_149),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_309),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_231),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_138),
.Y(n_287)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_145),
.B(n_1),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_153),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_289),
.B(n_290),
.Y(n_370)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_226),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_169),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_291),
.B(n_303),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_202),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_171),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_209),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_222),
.A2(n_5),
.B1(n_186),
.B2(n_136),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_162),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_298),
.Y(n_333)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_170),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_300),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_191),
.B(n_155),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_202),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_304),
.Y(n_354)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_181),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_178),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_167),
.A2(n_193),
.B1(n_204),
.B2(n_144),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_225),
.B(n_215),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_306),
.B(n_185),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_307),
.B(n_308),
.Y(n_361)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_148),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_139),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_180),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_311),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_161),
.B(n_205),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_160),
.C(n_192),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_162),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_314),
.Y(n_360)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_184),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_178),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_315),
.A2(n_186),
.B1(n_139),
.B2(n_180),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_159),
.A2(n_207),
.B1(n_225),
.B2(n_188),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_214),
.B1(n_222),
.B2(n_213),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_198),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_327),
.A2(n_350),
.B1(n_352),
.B2(n_366),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_334),
.B(n_304),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_336),
.A2(n_357),
.B(n_245),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_345),
.B(n_369),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_346),
.A2(n_365),
.B1(n_377),
.B2(n_332),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_306),
.A2(n_143),
.B1(n_219),
.B2(n_189),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_277),
.B1(n_312),
.B2(n_303),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_235),
.A2(n_195),
.B1(n_163),
.B2(n_216),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_235),
.A2(n_195),
.B1(n_163),
.B2(n_216),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_272),
.A2(n_177),
.B1(n_192),
.B2(n_179),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_355),
.A2(n_363),
.B1(n_332),
.B2(n_379),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_263),
.A2(n_202),
.B(n_226),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_236),
.B(n_241),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_364),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_248),
.B(n_177),
.CI(n_226),
.CON(n_363),
.SN(n_363)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_363),
.B(n_242),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_240),
.B(n_160),
.C(n_179),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_294),
.A2(n_189),
.B1(n_219),
.B2(n_228),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_317),
.A2(n_305),
.B1(n_279),
.B2(n_238),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_240),
.B(n_255),
.Y(n_369)
);

AOI32xp33_ASAP7_75t_L g372 ( 
.A1(n_278),
.A2(n_265),
.A3(n_255),
.B1(n_243),
.B2(n_294),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_271),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_279),
.A2(n_238),
.B1(n_286),
.B2(n_277),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_375),
.A2(n_364),
.B1(n_334),
.B2(n_333),
.Y(n_428)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_382),
.A2(n_387),
.B(n_388),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_357),
.A2(n_259),
.B(n_285),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_383),
.A2(n_380),
.B(n_379),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_401),
.B1(n_407),
.B2(n_415),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_301),
.B(n_312),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_386),
.B(n_392),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_378),
.A2(n_239),
.B(n_254),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_282),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_393),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_391),
.B(n_328),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_337),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_234),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_314),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_396),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_330),
.B(n_252),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_280),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_397),
.A2(n_402),
.B(n_420),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_366),
.A2(n_262),
.B1(n_246),
.B2(n_289),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_398),
.A2(n_413),
.B1(n_424),
.B2(n_370),
.Y(n_441)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_324),
.A2(n_233),
.B1(n_297),
.B2(n_250),
.Y(n_401)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_337),
.A2(n_261),
.B(n_267),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_330),
.B(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_348),
.B(n_269),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_406),
.B(n_416),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_324),
.A2(n_264),
.B1(n_268),
.B2(n_313),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_408),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_319),
.B(n_246),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_273),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_410),
.B(n_412),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_374),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_291),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_375),
.A2(n_315),
.B1(n_275),
.B2(n_309),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_326),
.A2(n_347),
.B1(n_350),
.B2(n_352),
.Y(n_414)
);

OA22x2_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_353),
.B1(n_335),
.B2(n_349),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_327),
.A2(n_311),
.B1(n_308),
.B2(n_283),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_308),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_368),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_421),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_351),
.B(n_274),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_418),
.B(n_419),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_351),
.B(n_283),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_320),
.A2(n_290),
.B(n_332),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_SL g423 ( 
.A(n_363),
.B(n_369),
.C(n_354),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_370),
.Y(n_454)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_426),
.A2(n_428),
.B1(n_430),
.B2(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_362),
.Y(n_427)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_429),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_338),
.A2(n_321),
.B1(n_340),
.B2(n_353),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_338),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_438),
.C(n_448),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_395),
.B(n_322),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_439),
.Y(n_504)
);

AOI322xp5_ASAP7_75t_L g440 ( 
.A1(n_387),
.A2(n_329),
.A3(n_361),
.B1(n_321),
.B2(n_374),
.C1(n_370),
.C2(n_340),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_440),
.B(n_388),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_399),
.B1(n_383),
.B2(n_386),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_413),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_395),
.B(n_343),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_389),
.B(n_341),
.C(n_343),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_458),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_409),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_451),
.B(n_454),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_397),
.A2(n_335),
.B1(n_376),
.B2(n_349),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_460),
.B1(n_399),
.B2(n_426),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_325),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_456),
.B(n_420),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_390),
.B(n_325),
.C(n_367),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_459),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_397),
.A2(n_380),
.B(n_373),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_462),
.A2(n_420),
.B(n_391),
.Y(n_495)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_419),
.B(n_331),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_467),
.B(n_468),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_406),
.B(n_331),
.Y(n_468)
);

XOR2x2_ASAP7_75t_L g470 ( 
.A(n_412),
.B(n_428),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_470),
.Y(n_473)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_474),
.A2(n_479),
.B1(n_485),
.B2(n_490),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_475),
.B(n_493),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_400),
.Y(n_476)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_476),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_443),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_480),
.Y(n_531)
);

A2O1A1O1Ixp25_ASAP7_75t_L g481 ( 
.A1(n_470),
.A2(n_404),
.B(n_386),
.C(n_423),
.D(n_396),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_481),
.A2(n_495),
.B(n_459),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_381),
.Y(n_486)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_486),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_435),
.Y(n_487)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_422),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_488),
.B(n_499),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_436),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_489),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_460),
.A2(n_424),
.B1(n_414),
.B2(n_398),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_466),
.A2(n_392),
.B1(n_402),
.B2(n_421),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_491),
.A2(n_498),
.B1(n_505),
.B2(n_459),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_433),
.A2(n_398),
.B1(n_413),
.B2(n_382),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_492),
.A2(n_497),
.B1(n_416),
.B2(n_446),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_418),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_457),
.B(n_393),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_494),
.B(n_502),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_433),
.A2(n_384),
.B1(n_401),
.B2(n_411),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_437),
.A2(n_384),
.B1(n_411),
.B2(n_401),
.Y(n_498)
);

AO22x1_ASAP7_75t_L g499 ( 
.A1(n_453),
.A2(n_415),
.B1(n_407),
.B2(n_423),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_432),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_500),
.B(n_471),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_501),
.B(n_469),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_442),
.B(n_394),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_503),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_437),
.A2(n_441),
.B1(n_462),
.B2(n_431),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_438),
.B(n_411),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_510),
.Y(n_518)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_509),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_434),
.B(n_410),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_442),
.B(n_417),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_457),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_448),
.C(n_470),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_513),
.B(n_515),
.C(n_529),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_456),
.C(n_450),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_516),
.B(n_522),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_505),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_550),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_483),
.B(n_506),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_483),
.B(n_469),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_528),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_512),
.Y(n_524)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_524),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_487),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_525),
.B(n_536),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_449),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_439),
.C(n_458),
.Y(n_529)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_478),
.A2(n_449),
.B(n_431),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_461),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_534),
.B(n_535),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_461),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_512),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_476),
.B(n_447),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_537),
.B(n_499),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_473),
.B(n_447),
.C(n_472),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_539),
.B(n_549),
.C(n_518),
.Y(n_568)
);

XOR2x1_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_495),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_541),
.A2(n_490),
.B1(n_479),
.B2(n_492),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_488),
.Y(n_543)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_543),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_478),
.A2(n_446),
.B(n_444),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_545),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_546),
.A2(n_474),
.B1(n_496),
.B2(n_503),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_480),
.Y(n_547)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_547),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_473),
.B(n_444),
.C(n_443),
.Y(n_549)
);

XNOR2x1_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_533),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_545),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_556),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_550),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_557),
.A2(n_560),
.B1(n_562),
.B2(n_574),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_521),
.A2(n_497),
.B1(n_482),
.B2(n_498),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_514),
.A2(n_482),
.B1(n_477),
.B2(n_499),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_537),
.B(n_486),
.Y(n_564)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_564),
.Y(n_592)
);

FAx1_ASAP7_75t_SL g567 ( 
.A(n_540),
.B(n_481),
.CI(n_484),
.CON(n_567),
.SN(n_567)
);

AOI322xp5_ASAP7_75t_L g597 ( 
.A1(n_567),
.A2(n_527),
.A3(n_526),
.B1(n_532),
.B2(n_544),
.C1(n_538),
.C2(n_531),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_568),
.A2(n_570),
.B(n_559),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_517),
.B(n_500),
.Y(n_569)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_489),
.C(n_480),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_572),
.B(n_573),
.C(n_578),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_515),
.B(n_509),
.C(n_508),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_519),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_575),
.B(n_577),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_520),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_513),
.B(n_496),
.C(n_484),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_531),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_579),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_580),
.B(n_528),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_549),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_523),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_583),
.B(n_587),
.Y(n_621)
);

MAJx2_ASAP7_75t_L g584 ( 
.A(n_555),
.B(n_535),
.C(n_534),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_584),
.B(n_586),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_572),
.B(n_529),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_578),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_588),
.B(n_589),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_518),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_552),
.A2(n_565),
.B1(n_561),
.B2(n_574),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_590),
.A2(n_606),
.B1(n_557),
.B2(n_601),
.Y(n_624)
);

CKINVDCx14_ASAP7_75t_R g625 ( 
.A(n_591),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_555),
.B(n_539),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_564),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_573),
.B(n_516),
.C(n_548),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_598),
.C(n_558),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_566),
.B(n_546),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_595),
.B(n_600),
.Y(n_608)
);

OA22x2_ASAP7_75t_L g596 ( 
.A1(n_562),
.A2(n_526),
.B1(n_548),
.B2(n_544),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_596),
.B(n_571),
.Y(n_615)
);

AOI31xp33_ASAP7_75t_L g617 ( 
.A1(n_597),
.A2(n_599),
.A3(n_605),
.B(n_569),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_559),
.B(n_547),
.C(n_532),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_551),
.B(n_542),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_563),
.B(n_429),
.Y(n_604)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_604),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_554),
.B(n_429),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_590),
.A2(n_561),
.B(n_552),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_607),
.A2(n_609),
.B(n_600),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_585),
.A2(n_565),
.B(n_576),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_610),
.B(n_614),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_570),
.C(n_580),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_611),
.B(n_612),
.Y(n_641)
);

BUFx24_ASAP7_75t_SL g612 ( 
.A(n_588),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_579),
.C(n_571),
.Y(n_614)
);

NOR2x1_ASAP7_75t_SL g645 ( 
.A(n_615),
.B(n_620),
.Y(n_645)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_617),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_595),
.B(n_558),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_619),
.B(n_622),
.Y(n_638)
);

FAx1_ASAP7_75t_L g620 ( 
.A(n_586),
.B(n_567),
.CI(n_560),
.CON(n_620),
.SN(n_620)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_594),
.B(n_577),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_623),
.B(n_445),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_624),
.A2(n_602),
.B1(n_592),
.B2(n_596),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_602),
.A2(n_575),
.B1(n_567),
.B2(n_445),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_626),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_587),
.B(n_465),
.C(n_464),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_627),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_627),
.B(n_589),
.C(n_593),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_629),
.B(n_633),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_630),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_620),
.A2(n_609),
.B1(n_607),
.B2(n_615),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_618),
.B(n_598),
.C(n_584),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_634),
.B(n_639),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_635),
.A2(n_637),
.B1(n_608),
.B2(n_611),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_614),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_636),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_624),
.A2(n_603),
.B1(n_596),
.B2(n_583),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_620),
.A2(n_615),
.B1(n_625),
.B2(n_616),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_642),
.B(n_643),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_610),
.B(n_465),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_613),
.A2(n_445),
.B(n_427),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_644),
.B(n_613),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_648),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_630),
.B(n_622),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_649),
.B(n_658),
.Y(n_659)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_650),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_628),
.B(n_621),
.C(n_376),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_652),
.B(n_654),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_641),
.B(n_621),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_643),
.B(n_408),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_655),
.B(n_656),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_631),
.B(n_629),
.C(n_634),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_632),
.B(n_403),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_656),
.B(n_639),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_661),
.A2(n_662),
.B(n_663),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_653),
.B(n_638),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_647),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_646),
.B(n_637),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_667),
.B(n_651),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_668),
.B(n_669),
.C(n_671),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_666),
.Y(n_669)
);

AOI21xp33_ASAP7_75t_L g671 ( 
.A1(n_664),
.A2(n_647),
.B(n_657),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_SL g672 ( 
.A1(n_660),
.A2(n_645),
.B(n_633),
.C(n_640),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_672),
.B(n_673),
.C(n_642),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_665),
.B(n_650),
.C(n_652),
.Y(n_673)
);

OAI311xp33_ASAP7_75t_L g674 ( 
.A1(n_670),
.A2(n_645),
.A3(n_640),
.B1(n_659),
.C1(n_660),
.Y(n_674)
);

OAI321xp33_ASAP7_75t_L g678 ( 
.A1(n_674),
.A2(n_644),
.A3(n_405),
.B1(n_328),
.B2(n_342),
.C(n_373),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_675),
.B(n_649),
.C(n_635),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_677),
.A2(n_678),
.B(n_676),
.Y(n_679)
);

MAJx2_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_367),
.C(n_385),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_342),
.Y(n_681)
);


endmodule