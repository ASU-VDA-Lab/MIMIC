module fake_jpeg_21235_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_17),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_8),
.C(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_21),
.B1(n_0),
.B2(n_3),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_64),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_28),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_21),
.B1(n_18),
.B2(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_58),
.B1(n_74),
.B2(n_51),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_30),
.B1(n_22),
.B2(n_31),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_23),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_24),
.B1(n_16),
.B2(n_18),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_32),
.C(n_20),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_23),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_27),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_69),
.B1(n_73),
.B2(n_54),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_26),
.B1(n_32),
.B2(n_20),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_79),
.B1(n_88),
.B2(n_90),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_64),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_27),
.B(n_25),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_102),
.B(n_71),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_98),
.B1(n_49),
.B2(n_55),
.Y(n_118)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_91),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_95),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_19),
.B1(n_0),
.B2(n_5),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_73),
.B1(n_54),
.B2(n_48),
.Y(n_115)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_103),
.B1(n_10),
.B2(n_12),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_4),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_75),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_9),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_72),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_109),
.C(n_94),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_118),
.B1(n_88),
.B2(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_113),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_48),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_123),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_77),
.B(n_13),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_86),
.B1(n_94),
.B2(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_65),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_139),
.Y(n_156)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_107),
.B1(n_123),
.B2(n_127),
.Y(n_165)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_81),
.B1(n_102),
.B2(n_84),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_150),
.B1(n_91),
.B2(n_104),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_102),
.B1(n_76),
.B2(n_77),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_153),
.B1(n_118),
.B2(n_113),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_81),
.B1(n_94),
.B2(n_101),
.Y(n_150)
);

AO21x2_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_94),
.B(n_85),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_87),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_159),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_106),
.C(n_121),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_160),
.C(n_164),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_114),
.A3(n_117),
.B1(n_116),
.B2(n_130),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_129),
.C(n_109),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_151),
.A3(n_149),
.B1(n_150),
.B2(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_122),
.B(n_113),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_167),
.B(n_135),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_112),
.C(n_105),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_151),
.B1(n_153),
.B2(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_99),
.C(n_65),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_170),
.C(n_141),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_126),
.B(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_92),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_140),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_177),
.C(n_174),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_182),
.B(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_141),
.C(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_137),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_181),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_147),
.B(n_134),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_151),
.B1(n_148),
.B2(n_133),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_186),
.B1(n_155),
.B2(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_151),
.B1(n_146),
.B2(n_134),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_174),
.C(n_160),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_169),
.C(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_192),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_193),
.B1(n_196),
.B2(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_194),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_169),
.B1(n_158),
.B2(n_156),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_157),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_205),
.C(n_197),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_177),
.C(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_171),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_192),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_191),
.B(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_181),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_164),
.C(n_189),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_205),
.B(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.C(n_212),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_207),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_209),
.B(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_184),
.B1(n_139),
.B2(n_144),
.Y(n_223)
);


endmodule