module fake_ibex_1660_n_21 (n_1, n_4, n_3, n_6, n_5, n_2, n_0, n_21);

input n_1;
input n_4;
input n_3;
input n_6;
input n_5;
input n_2;
input n_0;

output n_21;


SDFHx1_ASAP7_75t_R g7 ( 
.CLK(n_4),
.D(n_3),
.SE(n_0),
.SI(n_1),
.QN(n_7)
);


endmodule