module fake_jpeg_7397_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_23),
.B1(n_19),
.B2(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_59),
.B1(n_30),
.B2(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_16),
.B(n_31),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_0),
.C(n_1),
.Y(n_80)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_18),
.B1(n_20),
.B2(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_30),
.B1(n_32),
.B2(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_77),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_56),
.B1(n_20),
.B2(n_17),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_91),
.B1(n_60),
.B2(n_27),
.Y(n_99)
);

AOI22x1_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_40),
.B1(n_16),
.B2(n_39),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_80),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_71),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_40),
.B1(n_36),
.B2(n_31),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_40),
.B(n_50),
.C(n_36),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_81),
.B1(n_24),
.B2(n_3),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_18),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_36),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_82),
.B1(n_90),
.B2(n_16),
.Y(n_109)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_40),
.B1(n_36),
.B2(n_22),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_35),
.B1(n_34),
.B2(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_22),
.B1(n_16),
.B2(n_24),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_40),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_50),
.C(n_36),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_34),
.B1(n_27),
.B2(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_117),
.CON(n_134),
.SN(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_110),
.B1(n_81),
.B2(n_88),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_88),
.B1(n_83),
.B2(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_67),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_24),
.A3(n_8),
.B1(n_9),
.B2(n_15),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_1),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_66),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_76),
.B1(n_64),
.B2(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_75),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_121),
.A2(n_103),
.B(n_92),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g180 ( 
.A1(n_125),
.A2(n_113),
.B1(n_8),
.B2(n_11),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_131),
.B(n_102),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_68),
.B1(n_81),
.B2(n_73),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_130),
.B1(n_132),
.B2(n_146),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_81),
.B1(n_73),
.B2(n_88),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_78),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_85),
.B1(n_84),
.B2(n_71),
.Y(n_132)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_139),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_79),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_142),
.C(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_141),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_64),
.C(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_76),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_148),
.B(n_99),
.C(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_89),
.B1(n_76),
.B2(n_24),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_89),
.B1(n_24),
.B2(n_10),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_150),
.A2(n_156),
.B(n_158),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_93),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_168),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_96),
.B(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_120),
.B(n_101),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_161),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_129),
.B(n_134),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_165),
.B(n_130),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_164),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_93),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_104),
.B(n_114),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_179),
.B1(n_180),
.B2(n_148),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_101),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_100),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_97),
.C(n_92),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_124),
.B1(n_140),
.B2(n_147),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_188),
.B1(n_190),
.B2(n_164),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_198),
.B(n_201),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_194),
.B1(n_206),
.B2(n_171),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_149),
.B1(n_135),
.B2(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_196),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_204),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_135),
.B1(n_136),
.B2(n_145),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_158),
.B1(n_153),
.B2(n_165),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_123),
.B1(n_3),
.B2(n_4),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_2),
.B(n_4),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_4),
.B(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_207),
.Y(n_217)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_211),
.B1(n_228),
.B2(n_231),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_160),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_216),
.C(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_162),
.B1(n_170),
.B2(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_224),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_192),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_195),
.C(n_163),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_152),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_220),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_168),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_155),
.B(n_151),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_223),
.B1(n_208),
.B2(n_189),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_208),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_183),
.C(n_199),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_182),
.C(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_218),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_215),
.B1(n_211),
.B2(n_209),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_237),
.C(n_238),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_198),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_229),
.B(n_186),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_200),
.B(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_246),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_233),
.B1(n_239),
.B2(n_201),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_234),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_268),
.B(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_269),
.C(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_244),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_248),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_254),
.B(n_182),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_250),
.B1(n_260),
.B2(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_255),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_279),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_263),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_237),
.B(n_252),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_274),
.B1(n_188),
.B2(n_271),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_277),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_247),
.B1(n_265),
.B2(n_269),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_291),
.B1(n_276),
.B2(n_283),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_292),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_283),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_293),
.C(n_285),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_296),
.B(n_295),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_288),
.B(n_291),
.C(n_289),
.Y(n_300)
);

AOI32xp33_ASAP7_75t_SL g301 ( 
.A1(n_300),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_14),
.Y(n_302)
);


endmodule