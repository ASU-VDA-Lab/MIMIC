module fake_jpeg_18501_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_17),
.Y(n_51)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_27),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_55),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_32),
.B(n_16),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_59),
.B(n_75),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_19),
.B1(n_21),
.B2(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_24),
.B1(n_33),
.B2(n_30),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_16),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_35),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_17),
.B1(n_19),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_18),
.B1(n_33),
.B2(n_30),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

OR2x4_ASAP7_75t_SL g75 ( 
.A(n_41),
.B(n_31),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_19),
.B(n_21),
.C(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_79),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_45),
.B1(n_38),
.B2(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_64),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_53),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_18),
.B1(n_23),
.B2(n_31),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_23),
.B1(n_31),
.B2(n_3),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_31),
.C(n_23),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_74),
.C(n_57),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_69),
.B1(n_50),
.B2(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_60),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_103),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_50),
.B1(n_60),
.B2(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_59),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_111),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_128),
.B1(n_99),
.B2(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_14),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_120),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_49),
.B(n_13),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_116),
.C(n_129),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_71),
.C(n_13),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_71),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_100),
.B1(n_99),
.B2(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_57),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_4),
.Y(n_127)
);

NOR2x1_ASAP7_75t_R g129 ( 
.A(n_91),
.B(n_4),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_5),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_84),
.B1(n_83),
.B2(n_79),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_139),
.B1(n_152),
.B2(n_10),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

AO221x1_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_153),
.B1(n_102),
.B2(n_6),
.C(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_95),
.C(n_90),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_131),
.B(n_110),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_100),
.B1(n_90),
.B2(n_104),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_106),
.B(n_109),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_158),
.B(n_159),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_165),
.B1(n_133),
.B2(n_162),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_123),
.B(n_117),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_123),
.B(n_117),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_172),
.B1(n_146),
.B2(n_144),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_124),
.C(n_130),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.C(n_156),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_115),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_154),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_164),
.B(n_143),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_115),
.B1(n_98),
.B2(n_102),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_15),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_12),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_176),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_181),
.C(n_178),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_172),
.A3(n_155),
.B1(n_167),
.B2(n_145),
.C1(n_166),
.C2(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_183),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_159),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_165),
.B1(n_138),
.B2(n_134),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_132),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_190),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_149),
.B1(n_158),
.B2(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_147),
.B1(n_171),
.B2(n_137),
.Y(n_197)
);

NAND4xp25_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_182),
.C(n_180),
.D(n_179),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_187),
.B(n_195),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_180),
.B(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_205),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_179),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_181),
.B(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_189),
.Y(n_210)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_211),
.B1(n_203),
.B2(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_190),
.C(n_102),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_193),
.C(n_11),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

OAI221xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_205),
.B1(n_199),
.B2(n_201),
.C(n_198),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_214),
.A2(n_208),
.B(n_209),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_12),
.C(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_212),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_218),
.B(n_10),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);


endmodule