module real_jpeg_16603_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AND2x2_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_3),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_3),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_4),
.B(n_44),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_4),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_4),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_5),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_5),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_56),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_9),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_10),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_10),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_10),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_10),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_10),
.B(n_156),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_116),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_114),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_17),
.B(n_73),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.C(n_57),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_18),
.B(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_20),
.B(n_26),
.C(n_34),
.Y(n_113)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_32),
.Y(n_112)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_30),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_35),
.B(n_39),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_37),
.Y(n_94)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_37),
.Y(n_129)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_37),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_41),
.B(n_57),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.C(n_53),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_42),
.B(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_47),
.B(n_53),
.Y(n_122)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_56),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_63),
.C(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_98),
.B2(n_99),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_86),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_84),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_113),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_112),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_134),
.B(n_179),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_132),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_119),
.B(n_132),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_130),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_121),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_130),
.B1(n_131),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_147),
.B(n_178),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_143),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_140),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_144),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_162),
.B(n_177),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_159),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_155),
.Y(n_167)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_168),
.B(n_176),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);


endmodule