module fake_jpeg_6897_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_0),
.B(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_4),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_12),
.B(n_1),
.Y(n_14)
);

NAND3xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_17),
.C(n_22),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_17),
.Y(n_28)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_25)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_14),
.A3(n_15),
.B1(n_18),
.B2(n_27),
.C1(n_24),
.C2(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_21),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_14),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_34),
.C(n_25),
.Y(n_39)
);

OAI21x1_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_32),
.B(n_38),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_15),
.Y(n_41)
);


endmodule