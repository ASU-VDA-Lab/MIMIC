module real_aes_2989_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_0), .B(n_141), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_1), .A2(n_135), .B(n_183), .Y(n_182) );
INVxp33_ASAP7_75t_L g751 ( .A(n_2), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_3), .B(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_4), .B(n_141), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_5), .B(n_152), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_6), .B(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g140 ( .A(n_7), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_8), .B(n_152), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_9), .Y(n_105) );
NAND2xp33_ASAP7_75t_L g203 ( .A(n_10), .B(n_150), .Y(n_203) );
AND2x2_ASAP7_75t_L g454 ( .A(n_11), .B(n_197), .Y(n_454) );
AND2x2_ASAP7_75t_L g462 ( .A(n_12), .B(n_164), .Y(n_462) );
INVx2_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
AOI221x1_ASAP7_75t_L g134 ( .A1(n_14), .A2(n_26), .B1(n_135), .B2(n_141), .C(n_148), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_15), .B(n_152), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_16), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_17), .Y(n_111) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_18), .A2(n_197), .B(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_19), .B(n_141), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_20), .B(n_130), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_21), .B(n_152), .Y(n_211) );
AO21x1_ASAP7_75t_L g222 ( .A1(n_22), .A2(n_141), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_23), .B(n_141), .Y(n_493) );
NOR2xp33_ASAP7_75t_SL g101 ( .A(n_24), .B(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g117 ( .A(n_24), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_25), .A2(n_88), .B1(n_141), .B2(n_523), .Y(n_522) );
NAND2x1_ASAP7_75t_L g160 ( .A(n_27), .B(n_152), .Y(n_160) );
NAND2x1_ASAP7_75t_L g190 ( .A(n_28), .B(n_150), .Y(n_190) );
OR2x2_ASAP7_75t_L g133 ( .A(n_29), .B(n_85), .Y(n_133) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_29), .A2(n_85), .B(n_132), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_30), .B(n_150), .Y(n_185) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_31), .A2(n_119), .B1(n_732), .B2(n_735), .C(n_736), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_31), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_32), .B(n_152), .Y(n_202) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_33), .A2(n_164), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_34), .B(n_150), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_35), .A2(n_135), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_36), .B(n_152), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_37), .A2(n_135), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g136 ( .A(n_38), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g147 ( .A(n_38), .B(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g531 ( .A(n_38), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g103 ( .A(n_39), .B(n_104), .C(n_106), .Y(n_103) );
OR2x6_ASAP7_75t_L g115 ( .A(n_39), .B(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_40), .B(n_141), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_41), .B(n_141), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_42), .B(n_152), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_43), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_44), .B(n_150), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_45), .B(n_141), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_46), .A2(n_135), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_47), .A2(n_135), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_48), .B(n_150), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_49), .B(n_150), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_50), .B(n_141), .Y(n_467) );
INVx1_ASAP7_75t_L g139 ( .A(n_51), .Y(n_139) );
INVx1_ASAP7_75t_L g144 ( .A(n_51), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_52), .B(n_152), .Y(n_460) );
OAI22xp33_ASAP7_75t_SL g747 ( .A1(n_53), .A2(n_430), .B1(n_431), .B2(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_53), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_54), .Y(n_737) );
AND2x2_ASAP7_75t_L g484 ( .A(n_55), .B(n_130), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_56), .B(n_150), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_57), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_58), .B(n_150), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_59), .A2(n_135), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_60), .B(n_141), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_61), .B(n_141), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_62), .A2(n_135), .B(n_475), .Y(n_474) );
AO21x1_ASAP7_75t_L g224 ( .A1(n_63), .A2(n_135), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g499 ( .A(n_64), .B(n_131), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_65), .B(n_141), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_66), .B(n_150), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_67), .B(n_141), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_68), .B(n_150), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_69), .A2(n_93), .B1(n_135), .B2(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g175 ( .A(n_70), .B(n_131), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_71), .B(n_152), .Y(n_496) );
INVx1_ASAP7_75t_L g137 ( .A(n_72), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_72), .Y(n_146) );
AND2x2_ASAP7_75t_L g194 ( .A(n_73), .B(n_164), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_74), .B(n_150), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_75), .A2(n_135), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_76), .A2(n_135), .B(n_441), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_77), .A2(n_135), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g479 ( .A(n_78), .B(n_131), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_79), .B(n_130), .Y(n_520) );
INVx1_ASAP7_75t_L g102 ( .A(n_80), .Y(n_102) );
AND2x2_ASAP7_75t_L g179 ( .A(n_81), .B(n_164), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_82), .B(n_141), .Y(n_213) );
AND2x2_ASAP7_75t_L g444 ( .A(n_83), .B(n_197), .Y(n_444) );
AND2x2_ASAP7_75t_L g223 ( .A(n_84), .B(n_204), .Y(n_223) );
AND2x2_ASAP7_75t_L g167 ( .A(n_86), .B(n_164), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_87), .B(n_150), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_89), .B(n_152), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_90), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_91), .A2(n_135), .B(n_210), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_92), .A2(n_135), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_94), .B(n_152), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_95), .B(n_152), .Y(n_184) );
BUFx2_ASAP7_75t_L g498 ( .A(n_96), .Y(n_498) );
BUFx2_ASAP7_75t_L g743 ( .A(n_97), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_98), .A2(n_135), .B(n_201), .Y(n_200) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_107), .B(n_750), .Y(n_99) );
INVx2_ASAP7_75t_L g753 ( .A(n_100), .Y(n_753) );
AND2x2_ASAP7_75t_SL g100 ( .A(n_101), .B(n_103), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_102), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_106), .B(n_114), .Y(n_113) );
OR2x6_ASAP7_75t_SL g429 ( .A(n_106), .B(n_114), .Y(n_429) );
AND2x6_ASAP7_75t_SL g731 ( .A(n_106), .B(n_115), .Y(n_731) );
OR2x2_ASAP7_75t_L g738 ( .A(n_106), .B(n_115), .Y(n_738) );
AO21x2_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_739), .B(n_744), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_118), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_SL g746 ( .A1(n_110), .A2(n_747), .B(n_749), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g749 ( .A(n_113), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_427), .B1(n_430), .B2(n_730), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_121), .A2(n_429), .B1(n_431), .B2(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_339), .Y(n_121) );
AND4x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_251), .C(n_278), .D(n_313), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_176), .B1(n_216), .B2(n_231), .C(n_235), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_155), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_126), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g292 ( .A(n_127), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g347 ( .A(n_127), .B(n_302), .Y(n_347) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g250 ( .A(n_128), .B(n_168), .Y(n_250) );
AND2x4_ASAP7_75t_L g286 ( .A(n_128), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g300 ( .A(n_128), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g217 ( .A(n_129), .Y(n_217) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_129), .Y(n_389) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_130), .A2(n_181), .B(n_182), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_130), .Y(n_193) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_130), .A2(n_439), .B(n_440), .Y(n_438) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_130), .A2(n_522), .B(n_528), .Y(n_521) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x4_ASAP7_75t_L g204 ( .A(n_132), .B(n_133), .Y(n_204) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
BUFx3_ASAP7_75t_L g527 ( .A(n_136), .Y(n_527) );
AND2x6_ASAP7_75t_L g150 ( .A(n_137), .B(n_143), .Y(n_150) );
INVx2_ASAP7_75t_L g533 ( .A(n_137), .Y(n_533) );
AND2x4_ASAP7_75t_L g529 ( .A(n_138), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g152 ( .A(n_139), .B(n_145), .Y(n_152) );
INVx2_ASAP7_75t_L g525 ( .A(n_139), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_140), .Y(n_526) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx5_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B(n_153), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_150), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_153), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_153), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_153), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_153), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_153), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_153), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_153), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_153), .A2(n_442), .B(n_443), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_153), .A2(n_451), .B(n_452), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_153), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_153), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_153), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_153), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_153), .A2(n_496), .B(n_497), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_SL g244 ( .A1(n_155), .A2(n_217), .B(n_245), .C(n_249), .Y(n_244) );
AND2x2_ASAP7_75t_L g265 ( .A(n_155), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_155), .B(n_217), .Y(n_405) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_168), .Y(n_155) );
INVx2_ASAP7_75t_L g285 ( .A(n_156), .Y(n_285) );
BUFx3_ASAP7_75t_L g301 ( .A(n_156), .Y(n_301) );
INVxp67_ASAP7_75t_L g305 ( .A(n_156), .Y(n_305) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_163), .B(n_167), .Y(n_156) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_157), .A2(n_163), .B(n_167), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_163), .A2(n_169), .B(n_175), .Y(n_168) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_163), .A2(n_169), .B(n_175), .Y(n_230) );
AO21x1_ASAP7_75t_SL g472 ( .A1(n_163), .A2(n_473), .B(n_479), .Y(n_472) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_163), .A2(n_473), .B(n_479), .Y(n_506) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_165), .A2(n_456), .B(n_462), .Y(n_455) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
INVx2_ASAP7_75t_L g284 ( .A(n_168), .Y(n_284) );
AND2x2_ASAP7_75t_L g290 ( .A(n_168), .B(n_263), .Y(n_290) );
AND2x2_ASAP7_75t_L g316 ( .A(n_168), .B(n_285), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AOI211xp5_ASAP7_75t_L g313 ( .A1(n_176), .A2(n_314), .B(n_317), .C(n_327), .Y(n_313) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_177), .B(n_195), .Y(n_176) );
OAI321xp33_ASAP7_75t_L g288 ( .A1(n_177), .A2(n_236), .A3(n_289), .B1(n_291), .B2(n_292), .C(n_294), .Y(n_288) );
AND2x2_ASAP7_75t_L g409 ( .A(n_177), .B(n_384), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_177), .Y(n_412) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_186), .Y(n_177) );
INVx5_ASAP7_75t_L g234 ( .A(n_178), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_178), .B(n_248), .Y(n_247) );
NOR2x1_ASAP7_75t_SL g279 ( .A(n_178), .B(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g324 ( .A(n_178), .Y(n_324) );
AND2x2_ASAP7_75t_L g426 ( .A(n_178), .B(n_196), .Y(n_426) );
OR2x6_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AND2x2_ASAP7_75t_L g233 ( .A(n_186), .B(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_186), .Y(n_243) );
INVx4_ASAP7_75t_L g248 ( .A(n_186), .Y(n_248) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_193), .B(n_194), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_192), .Y(n_187) );
AOI21x1_ASAP7_75t_L g447 ( .A1(n_193), .A2(n_448), .B(n_454), .Y(n_447) );
INVx1_ASAP7_75t_L g291 ( .A(n_195), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_R g394 ( .A1(n_195), .A2(n_233), .B(n_265), .C(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g414 ( .A(n_195), .B(n_239), .Y(n_414) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
INVx1_ASAP7_75t_L g232 ( .A(n_196), .Y(n_232) );
INVx2_ASAP7_75t_L g238 ( .A(n_196), .Y(n_238) );
OR2x2_ASAP7_75t_L g257 ( .A(n_196), .B(n_248), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_196), .B(n_280), .Y(n_326) );
BUFx3_ASAP7_75t_L g333 ( .A(n_196), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_197), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_204), .Y(n_198) );
INVx1_ASAP7_75t_SL g207 ( .A(n_204), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_204), .B(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_204), .A2(n_467), .B(n_468), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_204), .A2(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g296 ( .A(n_205), .Y(n_296) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_205), .Y(n_309) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g242 ( .A(n_206), .Y(n_242) );
INVx1_ASAP7_75t_L g351 ( .A(n_206), .Y(n_351) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_214), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_207), .B(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_207), .A2(n_208), .B(n_214), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_213), .Y(n_208) );
AND2x2_ASAP7_75t_L g252 ( .A(n_216), .B(n_253), .Y(n_252) );
OAI31xp33_ASAP7_75t_L g403 ( .A1(n_216), .A2(n_404), .A3(n_406), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_SL g421 ( .A(n_216), .Y(n_421) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
AOI21xp33_ASAP7_75t_L g235 ( .A1(n_217), .A2(n_236), .B(n_244), .Y(n_235) );
NAND2x1_ASAP7_75t_L g315 ( .A(n_217), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g344 ( .A(n_217), .Y(n_344) );
INVx2_ASAP7_75t_L g293 ( .A(n_218), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_218), .B(n_276), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_218), .B(n_275), .Y(n_385) );
NOR2xp33_ASAP7_75t_SL g393 ( .A(n_218), .B(n_344), .Y(n_393) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_230), .Y(n_218) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_219), .B(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g273 ( .A(n_219), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g302 ( .A(n_219), .B(n_284), .Y(n_302) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx2_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
OAI21x1_ASAP7_75t_SL g221 ( .A1(n_222), .A2(n_224), .B(n_228), .Y(n_221) );
INVx1_ASAP7_75t_L g229 ( .A(n_223), .Y(n_229) );
INVx2_ASAP7_75t_L g274 ( .A(n_230), .Y(n_274) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_230), .Y(n_334) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx1_ASAP7_75t_L g270 ( .A(n_232), .Y(n_270) );
AND2x2_ASAP7_75t_L g349 ( .A(n_232), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g260 ( .A(n_233), .B(n_254), .Y(n_260) );
INVx2_ASAP7_75t_SL g308 ( .A(n_233), .Y(n_308) );
INVx4_ASAP7_75t_L g239 ( .A(n_234), .Y(n_239) );
AND2x2_ASAP7_75t_L g337 ( .A(n_234), .B(n_280), .Y(n_337) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_234), .B(n_350), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_234), .B(n_248), .Y(n_372) );
INVx1_ASAP7_75t_L g378 ( .A(n_236), .Y(n_378) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g297 ( .A(n_237), .Y(n_297) );
OR2x2_ASAP7_75t_L g310 ( .A(n_237), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
OR2x2_ASAP7_75t_L g362 ( .A(n_238), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g392 ( .A(n_238), .B(n_280), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_239), .B(n_242), .Y(n_268) );
AND2x2_ASAP7_75t_L g360 ( .A(n_239), .B(n_350), .Y(n_360) );
AND2x4_ASAP7_75t_L g422 ( .A(n_239), .B(n_301), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
INVx2_ASAP7_75t_L g246 ( .A(n_241), .Y(n_246) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp67_ASAP7_75t_SL g245 ( .A(n_246), .B(n_247), .Y(n_245) );
OAI322xp33_ASAP7_75t_SL g258 ( .A1(n_246), .A2(n_259), .A3(n_261), .B1(n_264), .B2(n_267), .C1(n_269), .C2(n_271), .Y(n_258) );
INVx1_ASAP7_75t_L g416 ( .A(n_246), .Y(n_416) );
OR2x2_ASAP7_75t_L g269 ( .A(n_247), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g295 ( .A(n_248), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_248), .B(n_296), .Y(n_311) );
INVx2_ASAP7_75t_L g338 ( .A(n_248), .Y(n_338) );
AND2x4_ASAP7_75t_L g350 ( .A(n_248), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_SL g353 ( .A(n_250), .B(n_266), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_256), .B(n_258), .Y(n_251) );
AND2x2_ASAP7_75t_L g319 ( .A(n_253), .B(n_286), .Y(n_319) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_254), .B(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g277 ( .A(n_255), .Y(n_277) );
AND2x4_ASAP7_75t_SL g359 ( .A(n_255), .B(n_274), .Y(n_359) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g267 ( .A(n_257), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_260), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g395 ( .A(n_262), .B(n_359), .Y(n_395) );
NOR4xp25_ASAP7_75t_L g399 ( .A(n_262), .B(n_276), .C(n_316), .D(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g276 ( .A(n_263), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g312 ( .A(n_263), .B(n_287), .Y(n_312) );
AND2x4_ASAP7_75t_L g376 ( .A(n_263), .B(n_287), .Y(n_376) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_266), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
OR2x2_ASAP7_75t_L g365 ( .A(n_273), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g419 ( .A(n_273), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_274), .B(n_286), .Y(n_320) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AOI211xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_281), .B(n_288), .C(n_303), .Y(n_278) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_284), .B(n_287), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_285), .B(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g367 ( .A(n_285), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_286), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g382 ( .A(n_286), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_298), .Y(n_294) );
AND2x4_ASAP7_75t_L g331 ( .A(n_295), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g425 ( .A(n_295), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_SL g329 ( .A(n_301), .Y(n_329) );
AND2x2_ASAP7_75t_L g388 ( .A(n_302), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_306), .B(n_310), .C(n_312), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_304), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g380 ( .A(n_305), .B(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g401 ( .A(n_305), .B(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
OR2x2_ASAP7_75t_L g390 ( .A(n_308), .B(n_332), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_311), .A2(n_318), .B1(n_320), .B2(n_321), .Y(n_317) );
INVx1_ASAP7_75t_SL g408 ( .A(n_312), .Y(n_408) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_323), .B(n_332), .Y(n_374) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_326), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_334), .B2(n_335), .Y(n_327) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI21xp5_ASAP7_75t_SL g341 ( .A1(n_332), .A2(n_342), .B(n_345), .Y(n_341) );
AND2x2_ASAP7_75t_L g370 ( .A(n_332), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND3x2_ASAP7_75t_L g336 ( .A(n_333), .B(n_337), .C(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g398 ( .A(n_333), .B(n_355), .Y(n_398) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g383 ( .A(n_338), .B(n_384), .Y(n_383) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_340), .B(n_396), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_341), .B(n_356), .C(n_377), .D(n_394), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B1(n_352), .B2(n_354), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_348), .A2(n_362), .B1(n_382), .B2(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g363 ( .A(n_350), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_352), .A2(n_375), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx3_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B1(n_361), .B2(n_364), .C(n_368), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B1(n_374), .B2(n_375), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_371), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_371), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B1(n_383), .B2(n_385), .C(n_386), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B1(n_391), .B2(n_393), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_392), .A2(n_412), .B(n_413), .C(n_415), .Y(n_411) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_403), .C(n_410), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_417), .B1(n_420), .B2(n_422), .C(n_423), .Y(n_410) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
CKINVDCx11_ASAP7_75t_R g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_638), .Y(n_431) );
NOR3xp33_ASAP7_75t_SL g432 ( .A(n_433), .B(n_561), .C(n_596), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_463), .B(n_513), .C(n_551), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_445), .Y(n_435) );
AND2x2_ASAP7_75t_L g544 ( .A(n_436), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_436), .B(n_550), .Y(n_584) );
AND2x2_ASAP7_75t_L g609 ( .A(n_436), .B(n_564), .Y(n_609) );
INVx4_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
OR2x2_ASAP7_75t_L g547 ( .A(n_437), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g555 ( .A(n_437), .B(n_455), .Y(n_555) );
AND2x2_ASAP7_75t_L g563 ( .A(n_437), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g590 ( .A(n_437), .B(n_591), .Y(n_590) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_437), .B(n_593), .Y(n_601) );
AND2x4_ASAP7_75t_L g618 ( .A(n_437), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g656 ( .A(n_437), .Y(n_656) );
AND2x4_ASAP7_75t_SL g661 ( .A(n_437), .B(n_446), .Y(n_661) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_444), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_445), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_445), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_455), .Y(n_445) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_446), .Y(n_556) );
INVx2_ASAP7_75t_L g592 ( .A(n_446), .Y(n_592) );
INVx1_ASAP7_75t_L g619 ( .A(n_446), .Y(n_619) );
AND2x2_ASAP7_75t_L g718 ( .A(n_446), .B(n_628), .Y(n_718) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_447), .Y(n_550) );
AND2x2_ASAP7_75t_L g564 ( .A(n_447), .B(n_455), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_453), .Y(n_448) );
INVx2_ASAP7_75t_L g593 ( .A(n_455), .Y(n_593) );
INVx2_ASAP7_75t_L g628 ( .A(n_455), .Y(n_628) );
OR2x2_ASAP7_75t_L g713 ( .A(n_455), .B(n_545), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_480), .B(n_500), .C(n_507), .Y(n_463) );
INVx2_ASAP7_75t_SL g602 ( .A(n_464), .Y(n_602) );
AND2x2_ASAP7_75t_L g608 ( .A(n_464), .B(n_481), .Y(n_608) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_472), .Y(n_464) );
INVx1_ASAP7_75t_L g504 ( .A(n_465), .Y(n_504) );
INVx1_ASAP7_75t_L g510 ( .A(n_465), .Y(n_510) );
INVx2_ASAP7_75t_L g535 ( .A(n_465), .Y(n_535) );
AND2x2_ASAP7_75t_L g559 ( .A(n_465), .B(n_483), .Y(n_559) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_465), .Y(n_588) );
OR2x2_ASAP7_75t_L g668 ( .A(n_465), .B(n_491), .Y(n_668) );
AND2x2_ASAP7_75t_L g534 ( .A(n_472), .B(n_535), .Y(n_534) );
NOR2x1_ASAP7_75t_SL g566 ( .A(n_472), .B(n_491), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g580 ( .A(n_481), .B(n_503), .Y(n_580) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_491), .Y(n_481) );
OR2x2_ASAP7_75t_L g512 ( .A(n_482), .B(n_491), .Y(n_512) );
BUFx2_ASAP7_75t_L g536 ( .A(n_482), .Y(n_536) );
NOR2xp67_ASAP7_75t_L g587 ( .A(n_482), .B(n_588), .Y(n_587) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_483), .Y(n_539) );
AND2x2_ASAP7_75t_L g565 ( .A(n_483), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g575 ( .A(n_483), .Y(n_575) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_483), .B(n_491), .Y(n_613) );
OR2x2_ASAP7_75t_L g688 ( .A(n_483), .B(n_505), .Y(n_688) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_SL g501 ( .A(n_491), .Y(n_501) );
AND2x2_ASAP7_75t_L g560 ( .A(n_491), .B(n_505), .Y(n_560) );
AND2x2_ASAP7_75t_L g631 ( .A(n_491), .B(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g652 ( .A(n_491), .Y(n_652) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_499), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g574 ( .A(n_503), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
BUFx2_ASAP7_75t_L g569 ( .A(n_504), .Y(n_569) );
AND2x2_ASAP7_75t_L g541 ( .A(n_505), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g632 ( .A(n_505), .Y(n_632) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
OR2x2_ASAP7_75t_L g578 ( .A(n_509), .B(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_SL g620 ( .A(n_509), .B(n_621), .Y(n_620) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_509), .A2(n_536), .A3(n_658), .B1(n_660), .B2(n_663), .C1(n_665), .C2(n_667), .Y(n_657) );
AND2x2_ASAP7_75t_L g722 ( .A(n_509), .B(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_510), .B(n_536), .Y(n_546) );
AOI322xp5_ASAP7_75t_L g597 ( .A1(n_511), .A2(n_598), .A3(n_602), .B1(n_603), .B2(n_606), .C1(n_608), .C2(n_609), .Y(n_597) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g649 ( .A(n_512), .B(n_602), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_512), .A2(n_709), .B1(n_711), .B2(n_714), .Y(n_708) );
OR2x2_ASAP7_75t_L g726 ( .A(n_512), .B(n_675), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_536), .B(n_537), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
AOI221xp5_ASAP7_75t_SL g576 ( .A1(n_515), .A2(n_552), .B1(n_577), .B2(n_580), .C(n_581), .Y(n_576) );
AND2x2_ASAP7_75t_L g603 ( .A(n_515), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_516), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g645 ( .A(n_516), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g674 ( .A(n_517), .Y(n_674) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_534), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_518), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g616 ( .A(n_518), .Y(n_616) );
OR2x2_ASAP7_75t_L g623 ( .A(n_518), .B(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g666 ( .A(n_519), .B(n_628), .Y(n_666) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x4_ASAP7_75t_L g545 ( .A(n_520), .B(n_521), .Y(n_545) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
NOR2x1p5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_534), .B(n_595), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_534), .B(n_575), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_534), .Y(n_675) );
INVx1_ASAP7_75t_L g542 ( .A(n_535), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_543), .B1(n_546), .B2(n_547), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_SL g653 ( .A(n_541), .Y(n_653) );
AND2x2_ASAP7_75t_L g710 ( .A(n_542), .B(n_566), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_544), .B(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_SL g582 ( .A(n_544), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_544), .B(n_703), .Y(n_702) );
BUFx3_ASAP7_75t_L g570 ( .A(n_545), .Y(n_570) );
INVx2_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
AND2x2_ASAP7_75t_L g643 ( .A(n_545), .B(n_627), .Y(n_643) );
INVx1_ASAP7_75t_L g557 ( .A(n_547), .Y(n_557) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_557), .B(n_558), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g636 ( .A(n_555), .Y(n_636) );
INVx2_ASAP7_75t_L g624 ( .A(n_556), .Y(n_624) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g621 ( .A(n_560), .B(n_575), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_560), .A2(n_658), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_562), .B(n_576), .Y(n_561) );
AOI32xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .A3(n_567), .B1(n_571), .B2(n_574), .Y(n_562) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_563), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_563), .A2(n_652), .B1(n_670), .B2(n_672), .C(n_678), .Y(n_669) );
AND2x2_ASAP7_75t_L g689 ( .A(n_563), .B(n_570), .Y(n_689) );
BUFx2_ASAP7_75t_L g573 ( .A(n_564), .Y(n_573) );
INVx1_ASAP7_75t_L g698 ( .A(n_564), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_564), .Y(n_703) );
INVx1_ASAP7_75t_SL g696 ( .A(n_565), .Y(n_696) );
INVx2_ASAP7_75t_L g579 ( .A(n_566), .Y(n_579) );
AND2x2_ASAP7_75t_L g691 ( .A(n_567), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g663 ( .A(n_569), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g635 ( .A(n_570), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_570), .B(n_661), .Y(n_683) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g595 ( .A(n_575), .Y(n_595) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g585 ( .A(n_579), .B(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g594 ( .A(n_579), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g699 ( .A(n_580), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B1(n_589), .B2(n_594), .Y(n_581) );
INVx2_ASAP7_75t_SL g673 ( .A(n_583), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_583), .B(n_712), .Y(n_714) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_585), .A2(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g630 ( .A(n_587), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g658 ( .A(n_590), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g605 ( .A(n_591), .Y(n_605) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g647 ( .A(n_593), .Y(n_647) );
INVx1_ASAP7_75t_L g692 ( .A(n_594), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_610), .C(n_633), .Y(n_596) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx2_ASAP7_75t_L g659 ( .A(n_599), .Y(n_659) );
AND2x2_ASAP7_75t_L g677 ( .A(n_599), .B(n_618), .Y(n_677) );
OR2x2_ASAP7_75t_L g716 ( .A(n_599), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_600), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g612 ( .A(n_602), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g679 ( .A(n_605), .B(n_616), .Y(n_679) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_608), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g720 ( .A(n_608), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_614), .B1(n_618), .B2(n_620), .C(n_622), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_611), .A2(n_634), .B(n_637), .Y(n_633) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g664 ( .A(n_613), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_613), .B(n_707), .Y(n_706) );
INVxp33_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g625 ( .A(n_621), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B1(n_626), .B2(n_629), .Y(n_622) );
INVx2_ASAP7_75t_L g728 ( .A(n_624), .Y(n_728) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVxp67_ASAP7_75t_L g707 ( .A(n_632), .Y(n_707) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_684), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_657), .C(n_669), .D(n_681), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B(n_648), .C(n_650), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g680 ( .A(n_643), .Y(n_680) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_645), .A2(n_651), .B(n_654), .Y(n_650) );
INVx2_ASAP7_75t_L g729 ( .A(n_646), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_647), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g662 ( .A(n_647), .Y(n_662) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
OR2x2_ASAP7_75t_L g724 ( .A(n_652), .B(n_688), .Y(n_724) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_659), .Y(n_695) );
AND2x2_ASAP7_75t_SL g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g665 ( .A(n_661), .B(n_666), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_661), .A2(n_691), .B(n_693), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_661), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_SL g719 ( .A(n_661), .Y(n_719) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_685), .B(n_690), .C(n_700), .D(n_721), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_697), .B2(n_699), .Y(n_693) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI211xp5_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_704), .B(n_708), .C(n_715), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B(n_720), .Y(n_715) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_725), .B(n_727), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx3_ASAP7_75t_SL g734 ( .A(n_730), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
CKINVDCx6p67_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
BUFx3_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_741), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
endmodule