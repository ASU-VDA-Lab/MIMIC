module fake_jpeg_20030_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_46),
.B1(n_43),
.B2(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_78),
.B1(n_49),
.B2(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_1),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_46),
.B1(n_57),
.B2(n_55),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_59),
.B1(n_52),
.B2(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_85),
.B1(n_16),
.B2(n_32),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_50),
.B1(n_45),
.B2(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_1),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_21),
.C(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_90),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_24),
.B1(n_37),
.B2(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_91),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_17),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_14),
.Y(n_95)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_20),
.B1(n_35),
.B2(n_33),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_76),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_4),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_2),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_94),
.C(n_93),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_102),
.B(n_5),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_100),
.B(n_5),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_92),
.B1(n_100),
.B2(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_112),
.C(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_109),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_107),
.A3(n_105),
.B1(n_11),
.B2(n_12),
.C1(n_27),
.C2(n_8),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_118),
.B(n_39),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_9),
.Y(n_120)
);


endmodule