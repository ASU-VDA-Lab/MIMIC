module fake_jpeg_1851_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_60),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_5),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_49),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_11),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_68),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_14),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_3),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_4),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_37),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_32),
.B1(n_73),
.B2(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_86),
.B1(n_90),
.B2(n_108),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_84),
.B(n_93),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_41),
.B1(n_35),
.B2(n_40),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_92),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_32),
.B1(n_35),
.B2(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_43),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_94),
.B(n_102),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_118),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_23),
.B1(n_27),
.B2(n_7),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_50),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_5),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_27),
.B1(n_7),
.B2(n_8),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_106),
.A2(n_96),
.B(n_100),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_42),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_6),
.B1(n_45),
.B2(n_65),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_78),
.B1(n_85),
.B2(n_116),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_101),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_76),
.C(n_51),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_103),
.C(n_80),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_71),
.B1(n_62),
.B2(n_57),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_96),
.B1(n_118),
.B2(n_91),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_62),
.B(n_59),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_152),
.B(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_138),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_132),
.B(n_141),
.Y(n_163)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_55),
.B1(n_106),
.B2(n_81),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_140),
.B1(n_78),
.B2(n_85),
.Y(n_168)
);

AND2x4_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_144),
.Y(n_161)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_120),
.B1(n_113),
.B2(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_104),
.C(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_82),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_110),
.B1(n_116),
.B2(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_110),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_139),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_129),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_171),
.B1(n_179),
.B2(n_128),
.Y(n_185)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_178),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_128),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_144),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_128),
.B1(n_125),
.B2(n_130),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_126),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_182),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_145),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_183),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_124),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_153),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_179),
.B1(n_171),
.B2(n_175),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_166),
.A2(n_122),
.B(n_152),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_189),
.B(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_197),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_201),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_132),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_135),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_202),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_159),
.CI(n_161),
.CON(n_200),
.SN(n_200)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_158),
.C(n_163),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_157),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_204),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_158),
.B(n_162),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_173),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_215),
.B1(n_222),
.B2(n_195),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_212),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_200),
.Y(n_214)
);

OAI322xp33_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_220),
.A3(n_205),
.B1(n_202),
.B2(n_188),
.C1(n_200),
.C2(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_163),
.B1(n_183),
.B2(n_164),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_183),
.B(n_176),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_192),
.B(n_194),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_181),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_224),
.B(n_197),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_169),
.B1(n_170),
.B2(n_173),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_214),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_233),
.C(n_234),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_230),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

AO221x1_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_210),
.B1(n_215),
.B2(n_217),
.C(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_199),
.B1(n_195),
.B2(n_193),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_228),
.B1(n_231),
.B2(n_191),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_212),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_245),
.C(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_220),
.C(n_208),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_219),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_246),
.A2(n_232),
.B(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_247),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_160),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_237),
.B1(n_233),
.B2(n_228),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_241),
.B1(n_191),
.B2(n_245),
.Y(n_261)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_256),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_250),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_254),
.C(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_257),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_259),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_267),
.A2(n_260),
.B1(n_268),
.B2(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_244),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_271),
.B(n_266),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_169),
.Y(n_274)
);


endmodule