module fake_jpeg_12447_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_182;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_241;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_47),
.Y(n_98)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_15),
.B(n_1),
.CON(n_56),
.SN(n_56)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_31),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_3),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_3),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_63),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_72),
.B(n_76),
.Y(n_131)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_20),
.B1(n_35),
.B2(n_21),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_75),
.A2(n_25),
.B(n_19),
.Y(n_142)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_30),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_91),
.Y(n_115)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_84),
.Y(n_129)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_21),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_23),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_20),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_38),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_36),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_32),
.B1(n_23),
.B2(n_17),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_125),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_121),
.C(n_111),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_28),
.B(n_25),
.C(n_7),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_94),
.B(n_6),
.Y(n_157)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_17),
.Y(n_125)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_72),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_65),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_159),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_95),
.B1(n_70),
.B2(n_66),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_167),
.B1(n_168),
.B2(n_129),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_64),
.B1(n_67),
.B2(n_66),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_88),
.B1(n_128),
.B2(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_157),
.B(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_69),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_73),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_161),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_86),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_70),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_63),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_171),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_92),
.B1(n_89),
.B2(n_79),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_92),
.B1(n_89),
.B2(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_62),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_105),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_4),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_4),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_157),
.B(n_144),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_186),
.B1(n_189),
.B2(n_173),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_127),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_194),
.C(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_142),
.B(n_139),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_153),
.B(n_155),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_130),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_192),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_197),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_110),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_199),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_137),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_143),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_149),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_147),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_129),
.B1(n_137),
.B2(n_135),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_150),
.B(n_144),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_214),
.B(n_196),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_147),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_208),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_199),
.B(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_149),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_215),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_134),
.B(n_140),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_164),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_163),
.B(n_134),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_176),
.B1(n_138),
.B2(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_225),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_232),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_234),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_185),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_194),
.C(n_177),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_212),
.C(n_204),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_176),
.B(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_245),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_203),
.C(n_219),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_207),
.C(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_202),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_211),
.B1(n_206),
.B2(n_230),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_241),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_239),
.A2(n_230),
.B1(n_232),
.B2(n_222),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_201),
.B1(n_220),
.B2(n_228),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_238),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_254),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_241),
.A2(n_227),
.B1(n_201),
.B2(n_229),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_238),
.C(n_234),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_202),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_182),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_215),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_250),
.A3(n_254),
.B1(n_235),
.B2(n_225),
.C1(n_248),
.C2(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_265),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_264),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_213),
.A3(n_205),
.B1(n_198),
.B2(n_175),
.C1(n_158),
.C2(n_169),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_145),
.B1(n_156),
.B2(n_162),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_140),
.B(n_8),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_257),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_135),
.C(n_138),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_268),
.B1(n_145),
.B2(n_158),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_269),
.A3(n_272),
.B1(n_19),
.B2(n_10),
.C1(n_4),
.C2(n_9),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

XNOR2x2_ASAP7_75t_SL g279 ( 
.A(n_278),
.B(n_277),
.Y(n_279)
);


endmodule