module fake_jpeg_21473_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_240;
wire n_131;
wire n_56;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_59),
.B1(n_38),
.B2(n_39),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_59),
.B1(n_38),
.B2(n_40),
.Y(n_78)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_65),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_18),
.B1(n_16),
.B2(n_39),
.Y(n_73)
);

OAI211xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_44),
.B(n_45),
.C(n_57),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_30),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_81),
.Y(n_104)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_72),
.B1(n_47),
.B2(n_40),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_86),
.B(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_89),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_35),
.B(n_34),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_111),
.B1(n_58),
.B2(n_37),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_60),
.B(n_38),
.C(n_35),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_38),
.B1(n_40),
.B2(n_37),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_106),
.B1(n_58),
.B2(n_37),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_24),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_66),
.B(n_22),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_37),
.B1(n_40),
.B2(n_53),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_117),
.Y(n_150)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_21),
.B(n_66),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_129),
.B(n_136),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_119),
.Y(n_146)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_130),
.B1(n_99),
.B2(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_31),
.B1(n_40),
.B2(n_37),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_85),
.B1(n_80),
.B2(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_99),
.B1(n_95),
.B2(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_34),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_138),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_155),
.B1(n_129),
.B2(n_113),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_144),
.B1(n_128),
.B2(n_133),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_123),
.B1(n_134),
.B2(n_135),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_90),
.B(n_93),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_10),
.C(n_15),
.Y(n_186)
);

OAI211xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_87),
.B(n_97),
.C(n_104),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_53),
.A3(n_70),
.B1(n_61),
.B2(n_34),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_88),
.B1(n_104),
.B2(n_110),
.Y(n_148)
);

OAI22x1_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_151),
.B1(n_158),
.B2(n_147),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_110),
.B1(n_82),
.B2(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_89),
.B1(n_111),
.B2(n_98),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_111),
.B(n_107),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_62),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_162),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_111),
.B1(n_75),
.B2(n_58),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_166),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_62),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_35),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_56),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_34),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_20),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_131),
.C(n_132),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_177),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_127),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_146),
.B1(n_161),
.B2(n_139),
.Y(n_198)
);

OAI221xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_127),
.B1(n_29),
.B2(n_22),
.C(n_113),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_183),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_120),
.B1(n_101),
.B2(n_71),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_159),
.A2(n_101),
.B1(n_25),
.B2(n_34),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_186),
.B(n_154),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_159),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_51),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_149),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_195),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_164),
.C(n_168),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_163),
.C(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_25),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_216),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_146),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_163),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_25),
.B(n_23),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_141),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_23),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_25),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_180),
.B1(n_184),
.B2(n_183),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_84),
.B1(n_55),
.B2(n_2),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_84),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_218),
.B1(n_173),
.B2(n_8),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_171),
.B1(n_181),
.B2(n_175),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_195),
.C(n_175),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_207),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_193),
.C(n_176),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_230),
.C(n_205),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_228),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_231),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_176),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_197),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_23),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_12),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_215),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_245),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_209),
.B1(n_210),
.B2(n_214),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_247),
.B1(n_251),
.B2(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_209),
.C(n_215),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.C(n_224),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_200),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_210),
.B1(n_198),
.B2(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_248),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_235),
.A2(n_216),
.B1(n_196),
.B2(n_212),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_221),
.B1(n_196),
.B2(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_231),
.C(n_232),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_204),
.C(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_229),
.C(n_217),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_263),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_13),
.C(n_12),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_12),
.C(n_11),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_242),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_250),
.B1(n_249),
.B2(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_275),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_254),
.B(n_9),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_248),
.B(n_11),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_0),
.Y(n_279)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_11),
.A3(n_10),
.B1(n_9),
.B2(n_7),
.C(n_4),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_0),
.B(n_1),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_266),
.A2(n_253),
.B(n_254),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_272),
.B(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_282),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_7),
.B(n_1),
.C(n_3),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_0),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_3),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_275),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

OA21x2_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_270),
.B(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_5),
.B1(n_6),
.B2(n_287),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_289),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_286),
.B(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_291),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_292),
.C(n_284),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_5),
.B(n_6),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_5),
.Y(n_298)
);


endmodule