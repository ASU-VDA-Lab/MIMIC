module real_jpeg_18377_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_531),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_0),
.B(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_1),
.A2(n_13),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_1),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_1),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_1),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_1),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_2),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_2),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_3),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_3),
.B(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_4),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_4),
.Y(n_461)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_5),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_6),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_6),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_6),
.B(n_38),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_6),
.B(n_153),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_6),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_6),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_6),
.B(n_323),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_7),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_7),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_7),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_7),
.B(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_7),
.B(n_490),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_7),
.B(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_7),
.B(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_8),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_8),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_8),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_8),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_8),
.B(n_322),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_9),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_9),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_10),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_12),
.B(n_72),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_12),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_12),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_12),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_12),
.B(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_12),
.B(n_103),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_12),
.B(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_12),
.B(n_503),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_13),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_13),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_13),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_15),
.Y(n_532)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_16),
.Y(n_143)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_16),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_16),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_17),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_73),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_23),
.B(n_73),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_53),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.C(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_26),
.A2(n_27),
.B1(n_63),
.B2(n_64),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_26),
.B(n_166),
.C(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_26),
.A2(n_27),
.B1(n_236),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_63),
.C(n_67),
.Y(n_62)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_32),
.B(n_128),
.C(n_134),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_32),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_35),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_46),
.B2(n_50),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_36),
.B(n_249),
.C(n_259),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_36),
.A2(n_37),
.B1(n_259),
.B2(n_260),
.Y(n_307)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_38),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_39),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_80),
.C(n_86),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_41),
.A2(n_51),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_46),
.B(n_140),
.C(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_46),
.B(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.C(n_62),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_60),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_61),
.Y(n_217)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_63),
.A2(n_64),
.B1(n_101),
.B2(n_102),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_63),
.A2(n_64),
.B1(n_159),
.B2(n_160),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_101),
.C(n_106),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_64),
.B(n_160),
.C(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.C(n_97),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_90),
.C(n_94),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_83),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_84),
.Y(n_278)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_85),
.Y(n_372)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_86),
.B(n_210),
.C(n_213),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_86),
.B(n_213),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_88),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_89),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_93),
.Y(n_365)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_94),
.B(n_209),
.C(n_215),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_94),
.A2(n_95),
.B1(n_215),
.B2(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_172),
.C(n_177),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_95),
.B(n_178),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.C(n_109),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_101),
.A2(n_102),
.B1(n_139),
.B2(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_101),
.A2(n_102),
.B1(n_325),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_139),
.C(n_144),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_102),
.B(n_325),
.C(n_328),
.Y(n_324)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_126),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_110),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21x1_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_180),
.B(n_529),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_117),
.B(n_120),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_146),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_138),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_138),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_129),
.B1(n_134),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_134),
.A2(n_166),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_137),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_139),
.A2(n_140),
.B1(n_174),
.B2(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_140),
.B(n_256),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_140),
.B(n_272),
.Y(n_429)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_144),
.B(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_167),
.C(n_171),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_164),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_148),
.B(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_150),
.B(n_164),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_158),
.Y(n_457)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_173),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_198),
.C(n_201),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_174),
.A2(n_175),
.B1(n_201),
.B2(n_202),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_174),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_175),
.B(n_437),
.Y(n_481)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_176),
.Y(n_504)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_262),
.B(n_526),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_221),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_184),
.A2(n_527),
.B(n_528),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_185),
.B(n_187),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_192),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_190),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_208),
.C(n_218),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_194),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_206),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_195),
.B(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_197),
.B(n_206),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_199),
.B(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_199),
.B(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_201),
.A2(n_202),
.B1(n_320),
.B2(n_321),
.Y(n_387)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_202),
.B(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_208),
.B(n_218),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_245),
.Y(n_244)
);

XNOR2x2_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

OR2x6_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_222),
.B(n_224),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.C(n_230),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_225),
.B(n_228),
.Y(n_415)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_230),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.C(n_247),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_231),
.A2(n_232),
.B1(n_344),
.B2(n_346),
.Y(n_343)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_240),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_235),
.A2(n_240),
.B1(n_241),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_236),
.Y(n_333)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_244),
.A2(n_247),
.B1(n_248),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_244),
.Y(n_345)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_249),
.A2(n_250),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.C(n_256),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_256),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_254),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_256),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_257),
.Y(n_376)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2x1_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_417),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_351),
.B(n_410),
.C(n_411),
.D(n_416),
.Y(n_263)
);

NAND4xp25_ASAP7_75t_L g417 ( 
.A(n_264),
.B(n_411),
.C(n_418),
.D(n_420),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_337),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_265),
.B(n_337),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_310),
.C(n_314),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_266),
.A2(n_267),
.B1(n_311),
.B2(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_294),
.Y(n_267)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_268),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.C(n_279),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_269),
.B(n_402),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_273),
.A2(n_274),
.B1(n_279),
.B2(n_280),
.Y(n_402)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_274),
.A2(n_368),
.B(n_373),
.Y(n_367)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_287),
.C(n_291),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_291),
.Y(n_317)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_286),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_286),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_317),
.Y(n_316)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_305),
.B1(n_308),
.B2(n_309),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_295),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_298),
.B(n_299),
.C(n_302),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_298),
.B1(n_303),
.B2(n_304),
.Y(n_336)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_300),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_311),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_314),
.B(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_329),
.C(n_334),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_315),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.C(n_324),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_316),
.B(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_318),
.A2(n_319),
.B1(n_324),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_324),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_325),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_328),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_330),
.B(n_335),
.Y(n_399)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.C(n_341),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_342)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_344),
.Y(n_346)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_347),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_349),
.C(n_413),
.Y(n_412)
);

OAI21x1_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_404),
.B(n_409),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_397),
.Y(n_352)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_353),
.B(n_397),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_379),
.C(n_383),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_354),
.B(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_366),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_367),
.C(n_377),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.C(n_363),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_356),
.B(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_357),
.A2(n_358),
.B1(n_363),
.B2(n_364),
.Y(n_427)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_377),
.Y(n_366)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_379),
.A2(n_380),
.B1(n_383),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_383),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.C(n_388),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_384),
.B(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_388),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_395),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_389),
.B(n_395),
.Y(n_463)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_463),
.Y(n_462)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_398),
.B(n_401),
.C(n_403),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_419),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_406),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_414),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_443),
.B(n_525),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_440),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_422),
.B(n_440),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.C(n_428),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_423),
.A2(n_424),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_426),
.B(n_428),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.C(n_436),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_430),
.B1(n_431),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_436),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

AOI21x1_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_467),
.B(n_524),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_464),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_445),
.B(n_464),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.C(n_462),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_483),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_462),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_455),
.C(n_458),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_458),
.Y(n_472)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_484),
.B(n_523),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_482),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_469),
.B(n_482),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.C(n_480),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_471),
.B1(n_494),
.B2(n_496),
.Y(n_493)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_480),
.B1(n_481),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_473),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_474),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_487)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_497),
.B(n_522),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_493),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_486),
.B(n_493),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.C(n_492),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_506),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_488),
.A2(n_489),
.B1(n_492),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_492),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_494),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_498),
.A2(n_508),
.B(n_521),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_505),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_499),
.B(n_505),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_502),
.Y(n_514)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_515),
.B(n_520),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_514),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_510),
.B(n_514),
.Y(n_520)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);


endmodule