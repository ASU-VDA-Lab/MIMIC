module fake_netlist_6_279_n_69 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_69);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_69;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_37;
wire n_54;
wire n_33;
wire n_67;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_68;
wire n_55;
wire n_35;
wire n_58;
wire n_50;
wire n_49;
wire n_64;
wire n_43;
wire n_48;
wire n_47;
wire n_62;
wire n_31;
wire n_65;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_25),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_19),
.A2(n_29),
.B1(n_14),
.B2(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_0),
.Y(n_46)
);

AND2x6_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_32),
.B(n_38),
.Y(n_54)
);

O2A1O1Ixp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_45),
.B(n_42),
.C(n_35),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_44),
.B(n_43),
.Y(n_56)
);

OAI21x1_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_33),
.B(n_5),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_47),
.Y(n_59)
);

AO21x2_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_4),
.B(n_6),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

O2A1O1Ixp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_59),
.B(n_55),
.C(n_60),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_57),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_64)
);

NOR3x1_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_9),
.C(n_20),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OR2x6_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_64),
.Y(n_69)
);


endmodule