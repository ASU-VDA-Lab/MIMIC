module real_jpeg_12095_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_342, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_342;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_4),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_5),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_5),
.A2(n_45),
.B1(n_47),
.B2(n_124),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_59),
.B1(n_62),
.B2(n_124),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_5),
.A2(n_34),
.B1(n_40),
.B2(n_124),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_59),
.B1(n_62),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_6),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_173),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_6),
.A2(n_45),
.B1(n_47),
.B2(n_173),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_34),
.B1(n_40),
.B2(n_173),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_7),
.A2(n_44),
.B1(n_59),
.B2(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_7),
.A2(n_44),
.B1(n_64),
.B2(n_65),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_7),
.A2(n_34),
.B1(n_40),
.B2(n_44),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_8),
.A2(n_39),
.B1(n_59),
.B2(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_8),
.A2(n_39),
.B1(n_64),
.B2(n_65),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_9),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_9),
.A2(n_59),
.B1(n_62),
.B2(n_160),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_45),
.B1(n_47),
.B2(n_160),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_9),
.A2(n_34),
.B1(n_40),
.B2(n_160),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_10),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_45),
.B1(n_47),
.B2(n_68),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_34),
.B1(n_40),
.B2(n_68),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_12),
.A2(n_45),
.B1(n_47),
.B2(n_70),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_34),
.B1(n_40),
.B2(n_70),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_16),
.A2(n_45),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_16),
.A2(n_54),
.B1(n_59),
.B2(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_16),
.A2(n_34),
.B1(n_40),
.B2(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_16),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_17),
.A2(n_59),
.B1(n_62),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_17),
.A2(n_64),
.B1(n_65),
.B2(n_76),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_17),
.A2(n_45),
.B1(n_47),
.B2(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_17),
.A2(n_34),
.B1(n_40),
.B2(n_76),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_18),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_18),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_18),
.A2(n_64),
.B(n_200),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_18),
.A2(n_45),
.B1(n_47),
.B2(n_191),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_18),
.A2(n_47),
.B(n_50),
.C(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_18),
.B(n_83),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_18),
.B(n_37),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_18),
.B(n_55),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_18),
.A2(n_62),
.B(n_77),
.C(n_262),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_339),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_19),
.B(n_340),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_334),
.B(n_337),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_326),
.B(n_330),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_313),
.B(n_325),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_138),
.B(n_310),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_125),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_100),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_27),
.B(n_100),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_71),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_28),
.B(n_86),
.C(n_98),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_56),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_29),
.A2(n_30),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_31),
.A2(n_32),
.B1(n_56),
.B2(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_31),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_37),
.B(n_38),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_33),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_33),
.A2(n_37),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_33),
.A2(n_37),
.B1(n_180),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_33),
.A2(n_37),
.B1(n_151),
.B2(n_181),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_33),
.A2(n_37),
.B1(n_194),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_33),
.A2(n_37),
.B1(n_191),
.B2(n_247),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_33),
.A2(n_37),
.B1(n_240),
.B2(n_247),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_34),
.B(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_36),
.A2(n_114),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_36),
.A2(n_149),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_40),
.A2(n_51),
.B(n_191),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_43),
.A2(n_48),
.B1(n_55),
.B2(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_47),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_45),
.A2(n_62),
.A3(n_79),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_47),
.B(n_80),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_53),
.B1(n_55),
.B2(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_55),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_48),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_48),
.A2(n_55),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_48),
.A2(n_55),
.B1(n_154),
.B2(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_48),
.A2(n_55),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_48),
.A2(n_55),
.B1(n_226),
.B2(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_52),
.A2(n_118),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_52),
.A2(n_155),
.B1(n_184),
.B2(n_264),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_56),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_57),
.A2(n_58),
.B1(n_89),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_57),
.A2(n_58),
.B1(n_123),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_57),
.A2(n_58),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_57),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_58),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_62),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_59),
.B(n_191),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_201),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_60),
.B(n_62),
.Y(n_215)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_65),
.B(n_191),
.Y(n_201)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_86),
.B1(n_98),
.B2(n_99),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_73),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_84),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_81),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_82),
.B1(n_83),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_83),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_77),
.A2(n_83),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_77),
.A2(n_83),
.B(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_96),
.B1(n_120),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_81),
.A2(n_120),
.B1(n_121),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_81),
.A2(n_120),
.B1(n_175),
.B2(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_81),
.A2(n_172),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_88),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_92),
.C(n_94),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_88),
.B(n_128),
.C(n_131),
.Y(n_314)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_97),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_92),
.B(n_134),
.C(n_136),
.Y(n_324)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_108),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.C(n_122),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_110),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_295)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_122),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_125),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_126),
.B(n_127),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_135),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_137),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_163),
.B(n_309),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_161),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_140),
.B(n_161),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_145),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_141),
.B(n_144),
.Y(n_307)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_145),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.C(n_158),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_146),
.A2(n_147),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_148),
.B(n_152),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_156),
.B(n_158),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_157),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_159),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_304),
.B(n_308),
.Y(n_163)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_291),
.B1(n_302),
.B2(n_303),
.C(n_342),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_275),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_218),
.B(n_274),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_195),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_168),
.B(n_195),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_182),
.C(n_186),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_169),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_177),
.C(n_179),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_178),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_178),
.A2(n_288),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_178),
.A2(n_288),
.B1(n_321),
.B2(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_178),
.A2(n_288),
.B(n_328),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_190),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_209),
.B2(n_217),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_196),
.B(n_210),
.C(n_216),
.Y(n_276)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_198),
.B(n_204),
.C(n_208),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_202),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_211),
.B(n_214),
.Y(n_290)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_268),
.B(n_273),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_256),
.B(n_267),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_236),
.B(n_255),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_222),
.B(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_232),
.C(n_234),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_244),
.B(n_254),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_250),
.B(n_253),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_251),
.B(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_286),
.C(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_301),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_300),
.C(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_315),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_324),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_322),
.C(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_335),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_336),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);


endmodule