module fake_jpeg_7000_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_15),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_25),
.B1(n_16),
.B2(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_44),
.A2(n_48),
.B1(n_62),
.B2(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_51),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_26),
.C(n_32),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_53),
.C(n_18),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_25),
.B1(n_16),
.B2(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_54),
.B1(n_59),
.B2(n_11),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_22),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_31),
.B1(n_21),
.B2(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_10),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_67),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_83),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_11),
.B(n_15),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_87),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_69),
.B1(n_43),
.B2(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_56),
.B1(n_46),
.B2(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_71),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_73),
.Y(n_109)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_78),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_44),
.C(n_60),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_89),
.C(n_90),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_50),
.Y(n_82)
);

CKINVDCx10_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_94),
.B1(n_21),
.B2(n_19),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

OR2x4_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_53),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_22),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_42),
.B(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_44),
.B(n_62),
.C(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_112),
.B1(n_118),
.B2(n_78),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_73),
.B1(n_72),
.B2(n_81),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_63),
.B1(n_47),
.B2(n_49),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_19),
.B1(n_21),
.B2(n_2),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_93),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_120),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_22),
.C(n_17),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_82),
.C(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_22),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_17),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_131),
.C(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_64),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_132),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_138),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_65),
.B(n_84),
.C(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_145),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_17),
.B(n_22),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_136),
.B(n_149),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_17),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_17),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_91),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_147),
.B1(n_138),
.B2(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_86),
.C(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_0),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_1),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_1),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_9),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_121),
.B1(n_122),
.B2(n_118),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_112),
.B1(n_120),
.B2(n_117),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_19),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_152),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_75),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_105),
.B1(n_113),
.B2(n_10),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_109),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_175),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_122),
.B(n_114),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_173),
.B(n_177),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_164),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_176),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_170),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_114),
.B(n_101),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_95),
.B1(n_101),
.B2(n_110),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_101),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_95),
.B(n_116),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_105),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_113),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_148),
.C(n_136),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_181),
.C(n_172),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_188),
.B(n_194),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_149),
.B(n_95),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_144),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_183),
.B(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_204),
.C(n_180),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_141),
.B(n_96),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_156),
.B1(n_165),
.B2(n_167),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_119),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_206),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_172),
.B1(n_171),
.B2(n_153),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_184),
.B1(n_170),
.B2(n_169),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_1),
.C(n_2),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_1),
.B(n_3),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_164),
.B(n_3),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_9),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_159),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_217),
.C(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_182),
.C(n_173),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_176),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_166),
.C(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_186),
.C(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

XOR2x1_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_177),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_227),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_155),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_190),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_158),
.B1(n_165),
.B2(n_156),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_231),
.B1(n_195),
.B2(n_197),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_178),
.B1(n_174),
.B2(n_157),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_206),
.B1(n_203),
.B2(n_209),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_157),
.B1(n_12),
.B2(n_13),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_210),
.B(n_196),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_12),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_237),
.B1(n_218),
.B2(n_226),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_201),
.B(n_203),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_245),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_244),
.B1(n_248),
.B2(n_222),
.Y(n_256)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_189),
.B1(n_209),
.B2(n_200),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_189),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_250),
.C(n_251),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_207),
.B1(n_191),
.B2(n_186),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_207),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_216),
.B(n_229),
.C(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_256),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_228),
.B1(n_185),
.B2(n_220),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_262),
.B1(n_265),
.B2(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_213),
.C(n_250),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_243),
.C(n_240),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_185),
.B1(n_187),
.B2(n_212),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_232),
.B1(n_233),
.B2(n_196),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_188),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_214),
.B1(n_188),
.B2(n_211),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_239),
.C(n_245),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_214),
.B1(n_204),
.B2(n_188),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_270),
.C(n_277),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_261),
.A2(n_235),
.B1(n_247),
.B2(n_239),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_272),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_249),
.B1(n_240),
.B2(n_234),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_276),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_251),
.B(n_234),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_256),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_217),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_6),
.C(n_7),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_286),
.C(n_275),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_281),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_277),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_282),
.A2(n_252),
.B1(n_265),
.B2(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_291),
.C(n_293),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_292),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_13),
.C2(n_289),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_254),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_280),
.B(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_284),
.B(n_12),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_296),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_13),
.B(n_7),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_295),
.B(n_297),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_300),
.A2(n_299),
.B(n_7),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_6),
.B(n_8),
.Y(n_302)
);


endmodule