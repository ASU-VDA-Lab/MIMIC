module fake_ibex_1922_n_7571 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_854, n_1008, n_458, n_244, n_73, n_343, n_310, n_714, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_7571);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_7571;

wire n_4557;
wire n_6873;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_7170;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_7029;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_7042;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_7262;
wire n_7551;
wire n_6616;
wire n_6848;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_7063;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_6744;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_7147;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_7067;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_6842;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_7485;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_7450;
wire n_7492;
wire n_6760;
wire n_7396;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_7082;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_7313;
wire n_7305;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_7332;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_7151;
wire n_2839;
wire n_7013;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_1070;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_6602;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_7397;
wire n_3979;
wire n_7324;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_7105;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_7560;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_7187;
wire n_4854;
wire n_6732;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_7229;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_7099;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_7251;
wire n_7189;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_6868;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_7507;
wire n_1305;
wire n_2088;
wire n_6724;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_7097;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_7241;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_7264;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_7372;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_7521;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_6926;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_7358;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_6878;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_7316;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_7207;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_7112;
wire n_7083;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_7026;
wire n_3572;
wire n_6114;
wire n_6996;
wire n_1121;
wire n_4823;
wire n_7366;
wire n_5195;
wire n_5541;
wire n_7033;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_7103;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_6864;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_7445;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_6941;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_6824;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_7140;
wire n_4225;
wire n_7169;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_6912;
wire n_3455;
wire n_6940;
wire n_1591;
wire n_7048;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_7303;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_7192;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_6802;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_7394;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_6855;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_7003;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_7161;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_6958;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_7226;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6711;
wire n_6124;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_7356;
wire n_5199;
wire n_7377;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_7315;
wire n_7360;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_7081;
wire n_6136;
wire n_7559;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_7446;
wire n_1201;
wire n_5859;
wire n_7224;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_7541;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_7131;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_7155;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6971;
wire n_7553;
wire n_6128;
wire n_2361;
wire n_6804;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_7338;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_7221;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_6714;
wire n_4114;
wire n_6983;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_6857;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_6859;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_7101;
wire n_2954;
wire n_6379;
wire n_6911;
wire n_6766;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_7173;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6893;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_7530;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_7349;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6850;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_6827;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_7068;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_6699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_6901;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_6773;
wire n_4416;
wire n_7430;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6765;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_7391;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_7283;
wire n_2884;
wire n_3383;
wire n_7148;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_6704;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_7254;
wire n_2654;
wire n_7199;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_7509;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_6939;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_6727;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_6883;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_7457;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_6950;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_7327;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6915;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_7025;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_6922;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6731;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_7090;
wire n_1857;
wire n_1997;
wire n_7174;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_7250;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_6902;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_6837;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_6767;
wire n_7102;
wire n_4858;
wire n_6733;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_6723;
wire n_3339;
wire n_7177;
wire n_6900;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_7539;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_7233;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_7031;
wire n_1517;
wire n_5973;
wire n_7012;
wire n_7238;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_7030;
wire n_7110;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_6856;
wire n_5770;
wire n_1763;
wire n_6976;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_7517;
wire n_2516;
wire n_2031;
wire n_7121;
wire n_1348;
wire n_7317;
wire n_1191;
wire n_4099;
wire n_7190;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_7429;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_6777;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_7390;
wire n_2410;
wire n_7145;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_7561;
wire n_7529;
wire n_6185;
wire n_6706;
wire n_5342;
wire n_6884;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_7533;
wire n_2758;
wire n_5787;
wire n_6745;
wire n_7210;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_7563;
wire n_4022;
wire n_5843;
wire n_1072;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_7191;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_6881;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_7136;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_7213;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_7034;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_6990;
wire n_3650;
wire n_6948;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_6816;
wire n_7512;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_6712;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_7098;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_7323;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_7149;
wire n_7219;
wire n_4919;
wire n_7320;
wire n_7175;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_7357;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_7449;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_7218;
wire n_6863;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_7292;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_7142;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_7428;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_6805;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_7133;
wire n_2641;
wire n_7306;
wire n_1077;
wire n_7202;
wire n_6771;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_6695;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_7138;
wire n_7370;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_6978;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_6910;
wire n_2394;
wire n_1572;
wire n_7236;
wire n_1245;
wire n_4867;
wire n_7387;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_7122;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6925;
wire n_7024;
wire n_6483;
wire n_4686;
wire n_7466;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_6800;
wire n_7410;
wire n_5186;
wire n_7257;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6944;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_6980;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_7282;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_7495;
wire n_7334;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_7346;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_7532;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_5397;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_7401;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_7245;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_6946;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_6897;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_7075;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6847;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5265;
wire n_5087;
wire n_4401;
wire n_4727;
wire n_7367;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_6737;
wire n_3005;
wire n_4627;
wire n_6936;
wire n_5107;
wire n_6780;
wire n_4309;
wire n_4027;
wire n_7132;
wire n_7486;
wire n_6758;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_7419;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_7201;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_7555;
wire n_1736;
wire n_6176;
wire n_7265;
wire n_7232;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_7023;
wire n_3675;
wire n_7227;
wire n_2749;
wire n_2378;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_7273;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_6909;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_7070;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_6989;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_7046;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_7194;
wire n_5097;
wire n_4688;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_7527;
wire n_7290;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_7146;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_6960;
wire n_1226;
wire n_7253;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_7434;
wire n_4421;
wire n_2322;
wire n_7477;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_7452;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_6823;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_7414;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_6725;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_7475;
wire n_7184;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_6914;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_7152;
wire n_4771;
wire n_4970;
wire n_4652;
wire n_6927;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_6916;
wire n_6973;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_7554;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_7114;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_7354;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_6808;
wire n_7037;
wire n_2537;
wire n_1130;
wire n_4545;
wire n_2643;
wire n_4246;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_6747;
wire n_7335;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_6787;
wire n_1970;
wire n_3946;
wire n_7183;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_6784;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_7433;
wire n_2269;
wire n_6741;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_6807;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_6795;
wire n_7437;
wire n_6898;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_6785;
wire n_7384;
wire n_6738;
wire n_3030;
wire n_5631;
wire n_6818;
wire n_5983;
wire n_7516;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_7393;
wire n_4517;
wire n_6021;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_6966;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_6899;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_7503;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_6754;
wire n_4067;
wire n_6822;
wire n_6796;
wire n_6849;
wire n_6836;
wire n_4997;
wire n_5906;
wire n_7355;
wire n_6755;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_7084;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_7515;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_7483;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_6717;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_6988;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_7256;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_7172;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_7117;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_6790;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_6840;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_7287;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_6748;
wire n_3788;
wire n_3448;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_7301;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_7156;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_6993;
wire n_2390;
wire n_7544;
wire n_7203;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5488;
wire n_3107;
wire n_5465;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_1053;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_7408;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_7476;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_7566;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_7307;
wire n_2787;
wire n_4540;
wire n_6987;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_7409;
wire n_7087;
wire n_3503;
wire n_2441;
wire n_7280;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_7107;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_6984;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6701;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_7288;
wire n_7248;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_6907;
wire n_4554;
wire n_1260;
wire n_7038;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_6730;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_7153;
wire n_5194;
wire n_7230;
wire n_4579;
wire n_5628;
wire n_6994;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_7308;
wire n_1775;
wire n_6889;
wire n_6361;
wire n_6803;
wire n_7481;
wire n_2570;
wire n_4025;
wire n_6751;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_7403;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_7369;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_6696;
wire n_2395;
wire n_7089;
wire n_6062;
wire n_4059;
wire n_7258;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_6943;
wire n_1832;
wire n_1128;
wire n_3398;
wire n_2376;
wire n_3718;
wire n_4878;
wire n_6252;
wire n_7080;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_7002;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_6726;
wire n_3238;
wire n_6740;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_6799;
wire n_2463;
wire n_6932;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_7008;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_7049;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_7062;
wire n_7493;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_6716;
wire n_6797;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_7215;
wire n_7340;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_7154;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_6965;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_7279;
wire n_7499;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_6846;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_7052;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_6931;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_6700;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_6853;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5425;
wire n_5035;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_7158;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_7299;
wire n_1830;
wire n_6770;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_7095;
wire n_7464;
wire n_1662;
wire n_7426;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_7076;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_7246;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_7459;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_7570;
wire n_2075;
wire n_4816;
wire n_6951;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_6949;
wire n_5096;
wire n_6480;
wire n_7380;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_7167;
wire n_7537;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_7455;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_6819;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_6937;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_7474;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_6860;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_6833;
wire n_2159;
wire n_6865;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_7135;
wire n_6794;
wire n_3637;
wire n_7216;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_7487;
wire n_5277;
wire n_5900;
wire n_7421;
wire n_3647;
wire n_6240;
wire n_3928;
wire n_3619;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_7399;
wire n_1956;
wire n_7186;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_6498;
wire n_6720;
wire n_1669;
wire n_7562;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_6854;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_7197;
wire n_7015;
wire n_1175;
wire n_4408;
wire n_6832;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_7066;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_6779;
wire n_2567;
wire n_5645;
wire n_7044;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_7329;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_7438;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_6887;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_6769;
wire n_6903;
wire n_2433;
wire n_7255;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_6861;
wire n_2130;
wire n_4862;
wire n_7270;
wire n_5114;
wire n_7071;
wire n_6697;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_6826;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_7235;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_7129;
wire n_4242;
wire n_7243;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_7342;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_7547;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_7310;
wire n_2911;
wire n_1828;
wire n_6972;
wire n_1389;
wire n_6380;
wire n_7200;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_6703;
wire n_7116;
wire n_4562;
wire n_1584;
wire n_7540;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6719;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_7208;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_7337;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_7055;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_7073;
wire n_2637;
wire n_7417;
wire n_7159;
wire n_5047;
wire n_5504;
wire n_7494;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_7314;
wire n_3791;
wire n_6904;
wire n_6778;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_7294;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_7016;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_6444;
wire n_7422;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_6749;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_6985;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_7178;
wire n_7330;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_7388;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_5308;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5982;
wire n_6692;
wire n_7079;
wire n_6590;
wire n_7536;
wire n_3036;
wire n_7209;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_7467;
wire n_4038;
wire n_5503;
wire n_7206;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_6702;
wire n_3046;
wire n_7505;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_5644;
wire n_7501;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_7490;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_7051;
wire n_7278;
wire n_2791;
wire n_1450;
wire n_7416;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_7447;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_7520;
wire n_4442;
wire n_5700;
wire n_7274;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_6820;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_6952;
wire n_3261;
wire n_5324;
wire n_7534;
wire n_6547;
wire n_7065;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_6995;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_7461;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_7326;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_7423;
wire n_3270;
wire n_5168;
wire n_7443;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_7556;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_6879;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_7104;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2673;
wire n_2430;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_7106;
wire n_3615;
wire n_7198;
wire n_7381;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_7182;
wire n_6310;
wire n_6852;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_6961;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_7126;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_6956;
wire n_5184;
wire n_6440;
wire n_7564;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_7524;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_6643;
wire n_2687;
wire n_3456;
wire n_6569;
wire n_6814;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_7176;
wire n_4159;
wire n_7056;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_7535;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_7368;
wire n_5464;
wire n_6895;
wire n_6548;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_6890;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_6789;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_6867;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_6764;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_6935;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_7382;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_7130;
wire n_6942;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6772;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_7469;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_6955;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_7427;
wire n_6908;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_7506;
wire n_3822;
wire n_1276;
wire n_6874;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_6736;
wire n_4259;
wire n_1620;
wire n_7376;
wire n_5196;
wire n_5086;
wire n_7018;
wire n_6025;
wire n_6168;
wire n_7498;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_7134;
wire n_3967;
wire n_2373;
wire n_7456;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_7480;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_7348;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_7383;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_7053;
wire n_5483;
wire n_6713;
wire n_6919;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_7557;
wire n_3779;
wire n_3203;
wire n_7240;
wire n_7468;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_6750;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_6981;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_6828;
wire n_5123;
wire n_6160;
wire n_7043;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_7074;
wire n_7119;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_6875;
wire n_1701;
wire n_5236;
wire n_7567;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_6870;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_6715;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_7386;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_7007;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_7027;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_7432;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_7009;
wire n_6140;
wire n_5903;
wire n_7263;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_6663;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_6844;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_6999;
wire n_4571;
wire n_7214;
wire n_6982;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_6843;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_6877;
wire n_2821;
wire n_6892;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_7162;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_7510;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_7268;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_7465;
wire n_4337;
wire n_4826;
wire n_7398;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_7304;
wire n_7036;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_7462;
wire n_2490;
wire n_3127;
wire n_7171;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_7293;
wire n_1264;
wire n_6752;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_7568;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_7363;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_6698;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6977;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_7511;
wire n_7028;
wire n_1628;
wire n_6810;
wire n_1773;
wire n_7237;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_7039;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_6791;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_6967;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_7442;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_6768;
wire n_2458;
wire n_7489;
wire n_7144;
wire n_3401;
wire n_3032;
wire n_7362;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_6947;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6938;
wire n_6260;
wire n_5244;
wire n_7453;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_6906;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_7124;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_6918;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_7143;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_6834;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_6812;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_7123;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_7072;
wire n_4175;
wire n_4458;
wire n_7488;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_6762;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_6992;
wire n_7109;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_7325;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_6759;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_7137;
wire n_4621;
wire n_7526;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_7350;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_7311;
wire n_7458;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_7244;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_7339;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_7247;
wire n_2346;
wire n_4695;
wire n_7331;
wire n_7128;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_7284;
wire n_4163;
wire n_7321;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_7309;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_7163;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_6886;
wire n_4832;
wire n_5229;
wire n_7054;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_1587;
wire n_2555;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_6959;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_7413;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_7185;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_6710;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_6945;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_6776;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_7336;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_6905;
wire n_7120;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_7374;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_7491;
wire n_6964;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_7001;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_7111;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_7519;
wire n_1642;
wire n_5744;
wire n_6798;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_7538;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_7165;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_6888;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_7389;
wire n_1501;
wire n_7418;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_7375;
wire n_7096;
wire n_5257;
wire n_7281;
wire n_7300;
wire n_4397;
wire n_6920;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_6781;
wire n_4229;
wire n_4294;
wire n_7085;
wire n_1919;
wire n_4351;
wire n_6811;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_6921;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_7212;
wire n_7285;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_7032;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_7125;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_7160;
wire n_7100;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_7319;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_7504;
wire n_1586;
wire n_3497;
wire n_6722;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_7371;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_7361;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_7440;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_7010;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_7289;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_7004;
wire n_7021;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_7234;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_6975;
wire n_7266;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6573;
wire n_6786;
wire n_6774;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_6851;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_7211;
wire n_4335;
wire n_7141;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_6729;
wire n_7150;
wire n_6882;
wire n_1168;
wire n_5500;
wire n_7378;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_7470;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_7420;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_7558;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_6998;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_6721;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_7484;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_7271;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_7322;
wire n_7549;
wire n_7022;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_6885;
wire n_7217;
wire n_7166;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_6806;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_6933;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_7297;
wire n_3613;
wire n_1383;
wire n_7546;
wire n_2057;
wire n_7179;
wire n_5984;
wire n_6385;
wire n_7415;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_7057;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_6793;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_6746;
wire n_4702;
wire n_1341;
wire n_7411;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_7108;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_7220;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_7223;
wire n_2544;
wire n_7261;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_7092;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_6728;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_7275;
wire n_3768;
wire n_4224;
wire n_7272;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_7436;
wire n_3181;
wire n_7249;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_7168;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_7091;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_6858;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_7228;
wire n_3272;
wire n_7353;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_6841;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_6896;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_6954;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_7000;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_7040;
wire n_6132;
wire n_7196;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6872;
wire n_6089;
wire n_5211;
wire n_7205;
wire n_1668;
wire n_7260;
wire n_7500;
wire n_5861;
wire n_7086;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_7569;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_7047;
wire n_7412;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_7077;
wire n_2164;
wire n_7565;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6831;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6968;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_7523;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_7402;
wire n_2876;
wire n_6670;
wire n_7473;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_7405;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_7343;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_6046;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_7252;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_6991;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_6705;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_7451;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_7188;
wire n_6913;
wire n_5467;
wire n_2646;
wire n_7525;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_7528;
wire n_7113;
wire n_4435;
wire n_1235;
wire n_6355;
wire n_4755;
wire n_6329;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_6734;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_7471;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_7296;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_6825;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_6743;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_7345;
wire n_7472;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4542;
wire n_4122;
wire n_5021;
wire n_2819;
wire n_5523;
wire n_5456;
wire n_1985;
wire n_1140;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_7157;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_6809;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_7115;
wire n_1884;
wire n_6632;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_7286;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_6871;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_7344;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_6953;
wire n_3145;
wire n_5682;
wire n_6891;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_7127;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_6979;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_7050;
wire n_3554;
wire n_7431;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_6930;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_7118;
wire n_7259;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_6821;
wire n_4137;
wire n_1485;
wire n_7448;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_6775;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_7518;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6815;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_7069;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_7478;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_7011;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_7482;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_6763;
wire n_6782;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_7552;
wire n_6839;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_7164;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_7017;
wire n_7454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_6761;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_6974;
wire n_1898;
wire n_1254;
wire n_7312;
wire n_6894;
wire n_2524;
wire n_3927;
wire n_7045;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_7277;
wire n_6099;
wire n_5939;
wire n_7502;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_6997;
wire n_3747;
wire n_1323;
wire n_6753;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_7359;
wire n_3632;
wire n_5200;
wire n_7225;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_7020;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_7392;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2187;
wire n_2105;
wire n_5780;
wire n_2642;
wire n_6924;
wire n_5485;
wire n_5737;
wire n_6876;
wire n_7424;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_6962;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_7059;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_6970;
wire n_5185;
wire n_6829;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_7522;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_6830;
wire n_3290;
wire n_7365;
wire n_3585;
wire n_7094;
wire n_2878;
wire n_1810;
wire n_7439;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_7035;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_6838;
wire n_2698;
wire n_6869;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_6735;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_6866;
wire n_4383;
wire n_7395;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_7005;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_6742;
wire n_3063;
wire n_4543;
wire n_6969;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_7180;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_6929;
wire n_2255;
wire n_1820;
wire n_6986;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_6709;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_7385;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_7444;
wire n_6756;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_7441;
wire n_6250;
wire n_6718;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_7078;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_7093;
wire n_1167;
wire n_7333;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_7508;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_6757;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_7496;
wire n_3649;
wire n_1838;
wire n_6880;
wire n_3824;
wire n_7425;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_7550;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_7302;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_7548;
wire n_5142;
wire n_1433;
wire n_6934;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_7019;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_7088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_7542;
wire n_4487;
wire n_7204;
wire n_7014;
wire n_1165;
wire n_6708;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_7341;
wire n_7407;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_7514;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_6801;
wire n_1547;
wire n_1542;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_7193;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_7373;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_7291;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_6707;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_7239;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_6835;
wire n_7406;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_6792;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_7513;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_6928;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_7242;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_7181;
wire n_1161;
wire n_1103;
wire n_6739;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_7139;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_7404;
wire n_2870;
wire n_6862;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_7328;
wire n_6783;
wire n_4738;
wire n_7231;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3557;
wire n_3380;
wire n_7435;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_7058;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_7041;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_6788;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_7364;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_7006;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_6817;
wire n_1661;
wire n_6261;
wire n_7276;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_7269;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_6845;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_7531;
wire n_7222;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_7463;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_7347;
wire n_4944;
wire n_7060;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_7064;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_6917;
wire n_7545;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_7479;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_7400;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_6813;
wire n_2670;
wire n_7379;
wire n_1745;
wire n_7318;
wire n_7352;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_7295;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_7267;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_7497;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_6963;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_7543;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_6923;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_7460;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_7061;
wire n_7351;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_7298;
wire n_2497;
wire n_7195;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_6957;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_704),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_748),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_742),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_91),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_533),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_436),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_923),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_912),
.Y(n_1056)
);

BUFx2_ASAP7_75t_SL g1057 ( 
.A(n_296),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_302),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_818),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_525),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_511),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_896),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_582),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_299),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_920),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1004),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_212),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_4),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_377),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_1007),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_794),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_52),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1040),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_1009),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_90),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_136),
.Y(n_1076)
);

BUFx10_ASAP7_75t_L g1077 ( 
.A(n_219),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_1026),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_927),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1044),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_897),
.Y(n_1081)
);

BUFx5_ASAP7_75t_L g1082 ( 
.A(n_631),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_441),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_62),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_732),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_950),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_820),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_126),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_1003),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_581),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_895),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_1023),
.Y(n_1092)
);

BUFx5_ASAP7_75t_L g1093 ( 
.A(n_175),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_396),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_914),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_886),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_392),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_521),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1015),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_132),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_72),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_227),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_916),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_882),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_928),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1014),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1001),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_660),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_306),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_434),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_943),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_939),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_659),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_648),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_432),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_907),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_432),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_909),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_709),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_833),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_652),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_215),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_107),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_656),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_946),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1036),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_807),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_946),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_520),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_862),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_693),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_157),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_249),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_380),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_926),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_717),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_249),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1013),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_650),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_811),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_129),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_403),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_387),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_941),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_720),
.Y(n_1145)
);

BUFx10_ASAP7_75t_L g1146 ( 
.A(n_924),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_872),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_936),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_421),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1030),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_934),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_698),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_19),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_879),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_279),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_656),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_823),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_466),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_363),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_101),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_420),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_99),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_406),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_51),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_899),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_875),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_341),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_967),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_113),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_201),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_130),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_705),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_629),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_795),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1019),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_957),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_670),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_661),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_107),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_568),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_842),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_590),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_821),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_651),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_173),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_482),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_543),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_73),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_747),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_899),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_696),
.Y(n_1191)
);

CKINVDCx16_ASAP7_75t_R g1192 ( 
.A(n_12),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_786),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_913),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_343),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_888),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_772),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_728),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_62),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_830),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_760),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_127),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_978),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1039),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1025),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_166),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1037),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_383),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_419),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_843),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_982),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_252),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_626),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_661),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_604),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_887),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1012),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_985),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_225),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_925),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_905),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_407),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_238),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_642),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_600),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_617),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_377),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_123),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_84),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_405),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_574),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_365),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_155),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1042),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1030),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_0),
.Y(n_1237)
);

BUFx5_ASAP7_75t_L g1238 ( 
.A(n_180),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_515),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_896),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_278),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_673),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_750),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_670),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_149),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_258),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_202),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_871),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_694),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_59),
.Y(n_1250)
);

BUFx5_ASAP7_75t_L g1251 ( 
.A(n_144),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_893),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_266),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1013),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_490),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_992),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_601),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1031),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_482),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_804),
.Y(n_1260)
);

BUFx5_ASAP7_75t_L g1261 ( 
.A(n_224),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_491),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_272),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_161),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_19),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_433),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_601),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1036),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_353),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_872),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_182),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_259),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1017),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_413),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_986),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_25),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_887),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_570),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_989),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_887),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1016),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1011),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_431),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_742),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_97),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_949),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_336),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_403),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_19),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_246),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_157),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_746),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_919),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_219),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_741),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_775),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_747),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_941),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_428),
.Y(n_1299)
);

CKINVDCx16_ASAP7_75t_R g1300 ( 
.A(n_1043),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_503),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_344),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_199),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_646),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_559),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_930),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_9),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_653),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_901),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_624),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_747),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_299),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_917),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_970),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_757),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_190),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_440),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_189),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_806),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_283),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_929),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_217),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_77),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_142),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_904),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_510),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_348),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_590),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_874),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_263),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_496),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_541),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_805),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_318),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_510),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_852),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_300),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_853),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1038),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_632),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_298),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_179),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_345),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_758),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_886),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_570),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_540),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_876),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_409),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_515),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_931),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_320),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_805),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_135),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_782),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_881),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1028),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_882),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_5),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_879),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_122),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_35),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_933),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_203),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_557),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_443),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_3),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_791),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_598),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_351),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_998),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_379),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_783),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_358),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_14),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_874),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1022),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_789),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_815),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_834),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1010),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1029),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_79),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_251),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_575),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_926),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_294),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_60),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_558),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_635),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_152),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_721),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_930),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_802),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_663),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_886),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_514),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_484),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_493),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_175),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_992),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_381),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_704),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_287),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_910),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1032),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_612),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_526),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_104),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_113),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_55),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_51),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_185),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1047),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_891),
.Y(n_1415)
);

BUFx10_ASAP7_75t_L g1416 ( 
.A(n_102),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_630),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_435),
.Y(n_1418)
);

BUFx10_ASAP7_75t_L g1419 ( 
.A(n_838),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_748),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_674),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_890),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_469),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_714),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_511),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_453),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_916),
.Y(n_1427)
);

BUFx10_ASAP7_75t_L g1428 ( 
.A(n_1048),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_192),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_922),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_965),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_666),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_467),
.Y(n_1433)
);

BUFx10_ASAP7_75t_L g1434 ( 
.A(n_757),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_817),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_782),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_446),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_125),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_209),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_549),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_718),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_736),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1038),
.Y(n_1443)
);

CKINVDCx14_ASAP7_75t_R g1444 ( 
.A(n_909),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_818),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_307),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_711),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_354),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_185),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_880),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1028),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_423),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_39),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_541),
.Y(n_1454)
);

CKINVDCx16_ASAP7_75t_R g1455 ( 
.A(n_263),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_787),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_259),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_908),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_628),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_442),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1012),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_316),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_238),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_247),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_816),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_SL g1466 ( 
.A(n_366),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_894),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_714),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_583),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_613),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_490),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_639),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_113),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_574),
.Y(n_1474)
);

CKINVDCx14_ASAP7_75t_R g1475 ( 
.A(n_357),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_136),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_885),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_54),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_762),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_556),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_538),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1006),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_896),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_447),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_742),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1021),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_423),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_196),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_805),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_407),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_44),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1046),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_385),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_696),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_918),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_544),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_275),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_892),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1018),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_932),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_841),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_436),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1041),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_635),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_686),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_907),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_167),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_493),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_547),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_269),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_75),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_203),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_359),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_126),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_403),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_513),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_12),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_7),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_937),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_159),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_547),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_351),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_487),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_921),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_615),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1045),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_597),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1035),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_156),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_889),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_950),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_500),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_435),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_158),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_513),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_662),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_34),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_681),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_434),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_989),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_277),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_665),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_560),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_372),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_142),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1027),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_925),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_487),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1014),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_473),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_590),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_123),
.Y(n_1552)
);

BUFx5_ASAP7_75t_L g1553 ( 
.A(n_514),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1047),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_59),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_416),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_11),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_838),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_534),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_191),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_516),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_179),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_550),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_830),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_745),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_997),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_169),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_324),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_166),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_866),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_550),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_584),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1019),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_87),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_158),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_945),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_849),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_686),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1045),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_801),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_397),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1024),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_711),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_56),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_13),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_615),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_869),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_81),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_606),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_603),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1022),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_903),
.Y(n_1592)
);

BUFx10_ASAP7_75t_L g1593 ( 
.A(n_906),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_352),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_154),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_438),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_47),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_569),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_333),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_70),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_62),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_219),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_915),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_918),
.Y(n_1604)
);

BUFx5_ASAP7_75t_L g1605 ( 
.A(n_255),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_935),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_281),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_902),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_959),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_528),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_92),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_297),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_724),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_976),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_432),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_312),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_107),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_856),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_539),
.Y(n_1619)
);

CKINVDCx16_ASAP7_75t_R g1620 ( 
.A(n_135),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_865),
.Y(n_1621)
);

BUFx10_ASAP7_75t_L g1622 ( 
.A(n_883),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_375),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_268),
.Y(n_1624)
);

BUFx10_ASAP7_75t_L g1625 ( 
.A(n_438),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_909),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_900),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_97),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_302),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_677),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1006),
.Y(n_1631)
);

CKINVDCx16_ASAP7_75t_R g1632 ( 
.A(n_61),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_451),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_203),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_790),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_157),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1025),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_123),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_427),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_614),
.Y(n_1640)
);

BUFx10_ASAP7_75t_L g1641 ( 
.A(n_855),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_877),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_412),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_824),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_913),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_738),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_57),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_662),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_171),
.Y(n_1649)
);

CKINVDCx16_ASAP7_75t_R g1650 ( 
.A(n_818),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_721),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_53),
.Y(n_1652)
);

BUFx5_ASAP7_75t_L g1653 ( 
.A(n_457),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_884),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_109),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_206),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_179),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_356),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_228),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_9),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1034),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_662),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_872),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_336),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_911),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_878),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_111),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_968),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_898),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_229),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_359),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_553),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_16),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_898),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_586),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_885),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_371),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_230),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_710),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_187),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_764),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1033),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_475),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_474),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_537),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_241),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_330),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_854),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_252),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_452),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_229),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1184),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1156),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1317),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1527),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1070),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1082),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1059),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1444),
.B(n_0),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1444),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1250),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1403),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1445),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1598),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1475),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1184),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1689),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1079),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1133),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1191),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1318),
.Y(n_1712)
);

BUFx10_ASAP7_75t_L g1713 ( 
.A(n_1089),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1475),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1068),
.Y(n_1715)
);

INVxp33_ASAP7_75t_L g1716 ( 
.A(n_1372),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1120),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1052),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1082),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1065),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1082),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1085),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1077),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1082),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1082),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1088),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1077),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1192),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1579),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1120),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1097),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1100),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1359),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1148),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1455),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1102),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1105),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1579),
.Y(n_1738)
);

INVxp33_ASAP7_75t_SL g1739 ( 
.A(n_1256),
.Y(n_1739)
);

CKINVDCx16_ASAP7_75t_R g1740 ( 
.A(n_1620),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1109),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1632),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1650),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1119),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1049),
.Y(n_1745)
);

INVxp33_ASAP7_75t_SL g1746 ( 
.A(n_1050),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1121),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1134),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1142),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1166),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1167),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1170),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1148),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1485),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1082),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1171),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1173),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1174),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1178),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1082),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1179),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1519),
.B(n_0),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1182),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1077),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1185),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1186),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1187),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1190),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1070),
.Y(n_1769)
);

CKINVDCx16_ASAP7_75t_R g1770 ( 
.A(n_1113),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1193),
.Y(n_1771)
);

INVxp33_ASAP7_75t_L g1772 ( 
.A(n_1466),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1196),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1113),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1485),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1510),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1419),
.Y(n_1777)
);

INVxp33_ASAP7_75t_L g1778 ( 
.A(n_1066),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1579),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1198),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1051),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1206),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1113),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1419),
.Y(n_1784)
);

NOR2xp67_ASAP7_75t_L g1785 ( 
.A(n_1201),
.B(n_1),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1212),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_1061),
.Y(n_1787)
);

CKINVDCx14_ASAP7_75t_R g1788 ( 
.A(n_1131),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1213),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1215),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1093),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1216),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1510),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1226),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1227),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1101),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1229),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1629),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1259),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1053),
.Y(n_1800)
);

BUFx2_ASAP7_75t_SL g1801 ( 
.A(n_1131),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1104),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1625),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1230),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1241),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1054),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1055),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1243),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1629),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1093),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1245),
.Y(n_1811)
);

CKINVDCx16_ASAP7_75t_R g1812 ( 
.A(n_1131),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1247),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1253),
.Y(n_1814)
);

CKINVDCx16_ASAP7_75t_R g1815 ( 
.A(n_1146),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1257),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1056),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1283),
.Y(n_1818)
);

CKINVDCx16_ASAP7_75t_R g1819 ( 
.A(n_1146),
.Y(n_1819)
);

INVxp33_ASAP7_75t_L g1820 ( 
.A(n_1073),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1287),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1060),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1288),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1302),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1146),
.Y(n_1825)
);

BUFx10_ASAP7_75t_L g1826 ( 
.A(n_1303),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1093),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1696),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1723),
.B(n_1203),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1717),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1717),
.Y(n_1831)
);

NOR2xp67_ASAP7_75t_L g1832 ( 
.A(n_1723),
.B(n_1292),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1788),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1770),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1734),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1734),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1812),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1815),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1775),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1819),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1774),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1775),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1692),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1746),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1716),
.Y(n_1845)
);

INVxp67_ASAP7_75t_SL g1846 ( 
.A(n_1712),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1740),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1742),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1730),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_1787),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1745),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_1796),
.Y(n_1852)
);

CKINVDCx20_ASAP7_75t_R g1853 ( 
.A(n_1802),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1753),
.Y(n_1854)
);

NOR2xp67_ASAP7_75t_L g1855 ( 
.A(n_1774),
.B(n_1316),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1754),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1769),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1781),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1714),
.Y(n_1859)
);

INVxp33_ASAP7_75t_SL g1860 ( 
.A(n_1727),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1776),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1793),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1715),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1693),
.B(n_1300),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1728),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1800),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1806),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1798),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1694),
.B(n_1326),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1695),
.B(n_1361),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1809),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1807),
.Y(n_1872)
);

CKINVDCx20_ASAP7_75t_R g1873 ( 
.A(n_1733),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1822),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1735),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1764),
.B(n_1555),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1706),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1707),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1708),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1817),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1743),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1718),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1697),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1720),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1719),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1722),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1783),
.B(n_1640),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1727),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1713),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1726),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1729),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1700),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1705),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1801),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1799),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1731),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1721),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1825),
.B(n_1062),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1713),
.B(n_1777),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1739),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1732),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1709),
.B(n_1063),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1736),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1699),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1826),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1737),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1741),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1710),
.B(n_1064),
.Y(n_1908)
);

NOR2xp67_ASAP7_75t_L g1909 ( 
.A(n_1784),
.B(n_1306),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1744),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1826),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1803),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1747),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1748),
.Y(n_1914)
);

CKINVDCx16_ASAP7_75t_R g1915 ( 
.A(n_1711),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1749),
.B(n_1067),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1724),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1750),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1751),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1752),
.Y(n_1920)
);

INVxp67_ASAP7_75t_SL g1921 ( 
.A(n_1756),
.Y(n_1921)
);

INVxp33_ASAP7_75t_SL g1922 ( 
.A(n_1698),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1701),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1702),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1757),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1703),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1704),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1758),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1759),
.Y(n_1929)
);

CKINVDCx20_ASAP7_75t_R g1930 ( 
.A(n_1772),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1761),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1763),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1765),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1762),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1766),
.Y(n_1935)
);

CKINVDCx20_ASAP7_75t_R g1936 ( 
.A(n_1767),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1768),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1771),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1773),
.Y(n_1939)
);

CKINVDCx20_ASAP7_75t_R g1940 ( 
.A(n_1780),
.Y(n_1940)
);

CKINVDCx20_ASAP7_75t_R g1941 ( 
.A(n_1782),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1786),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1789),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1785),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1790),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1792),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1794),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1795),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1797),
.Y(n_1949)
);

INVxp33_ASAP7_75t_SL g1950 ( 
.A(n_1785),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1725),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1804),
.Y(n_1952)
);

INVxp33_ASAP7_75t_SL g1953 ( 
.A(n_1805),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1808),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1811),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1813),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1814),
.Y(n_1957)
);

CKINVDCx20_ASAP7_75t_R g1958 ( 
.A(n_1816),
.Y(n_1958)
);

CKINVDCx20_ASAP7_75t_R g1959 ( 
.A(n_1818),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1821),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1823),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1824),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1755),
.Y(n_1963)
);

CKINVDCx20_ASAP7_75t_R g1964 ( 
.A(n_1778),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1760),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1820),
.Y(n_1966)
);

NOR2xp67_ASAP7_75t_L g1967 ( 
.A(n_1791),
.B(n_1307),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1810),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1827),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1779),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1779),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1729),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1729),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1738),
.B(n_1416),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1738),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1738),
.Y(n_1976)
);

CKINVDCx20_ASAP7_75t_R g1977 ( 
.A(n_1779),
.Y(n_1977)
);

INVxp33_ASAP7_75t_SL g1978 ( 
.A(n_1714),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1788),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1788),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1717),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1714),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1717),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1717),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1717),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1717),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1788),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1717),
.Y(n_1988)
);

BUFx10_ASAP7_75t_L g1989 ( 
.A(n_1714),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1770),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1717),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1717),
.Y(n_1992)
);

NOR2xp67_ASAP7_75t_L g1993 ( 
.A(n_1723),
.B(n_1308),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1717),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1717),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1788),
.Y(n_1996)
);

CKINVDCx16_ASAP7_75t_R g1997 ( 
.A(n_1770),
.Y(n_1997)
);

NOR2xp67_ASAP7_75t_L g1998 ( 
.A(n_1723),
.B(n_1312),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1717),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1717),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1714),
.B(n_1069),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1714),
.B(n_1072),
.Y(n_2002)
);

CKINVDCx20_ASAP7_75t_R g2003 ( 
.A(n_1770),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1717),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1717),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1696),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1696),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1714),
.B(n_1075),
.Y(n_2008)
);

CKINVDCx20_ASAP7_75t_R g2009 ( 
.A(n_1770),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1717),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1717),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1717),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1717),
.Y(n_2013)
);

INVxp67_ASAP7_75t_SL g2014 ( 
.A(n_1717),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1717),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1788),
.Y(n_2016)
);

CKINVDCx16_ASAP7_75t_R g2017 ( 
.A(n_1770),
.Y(n_2017)
);

XOR2xp5_ASAP7_75t_L g2018 ( 
.A(n_1787),
.B(n_1115),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1717),
.Y(n_2019)
);

INVxp33_ASAP7_75t_L g2020 ( 
.A(n_1716),
.Y(n_2020)
);

INVxp67_ASAP7_75t_SL g2021 ( 
.A(n_1717),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1788),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1770),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1717),
.Y(n_2024)
);

CKINVDCx16_ASAP7_75t_R g2025 ( 
.A(n_1770),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1723),
.B(n_1076),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1717),
.Y(n_2027)
);

INVxp33_ASAP7_75t_SL g2028 ( 
.A(n_1714),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1723),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1788),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1717),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1717),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1770),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1717),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1723),
.B(n_1081),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1723),
.B(n_1083),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1770),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1717),
.Y(n_2038)
);

BUFx2_ASAP7_75t_L g2039 ( 
.A(n_1788),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1770),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1788),
.Y(n_2041)
);

INVxp67_ASAP7_75t_L g2042 ( 
.A(n_1714),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1788),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1717),
.Y(n_2044)
);

CKINVDCx20_ASAP7_75t_R g2045 ( 
.A(n_1770),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1788),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1788),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1717),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1717),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_1717),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1717),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1770),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1717),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1788),
.Y(n_2054)
);

CKINVDCx16_ASAP7_75t_R g2055 ( 
.A(n_1770),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1717),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1717),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1788),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_1770),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1717),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2014),
.B(n_1093),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2014),
.B(n_1093),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1974),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_2039),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2020),
.B(n_1416),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1860),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2021),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2021),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1928),
.B(n_1416),
.Y(n_2069)
);

INVx4_ASAP7_75t_L g2070 ( 
.A(n_1905),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1953),
.B(n_1084),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_1964),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1929),
.B(n_1434),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1921),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_SL g2075 ( 
.A1(n_1850),
.A2(n_1853),
.B1(n_1852),
.B2(n_2018),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2050),
.B(n_1093),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1921),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1961),
.B(n_1093),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1966),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1961),
.B(n_1238),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1880),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_SL g2082 ( 
.A1(n_1895),
.A2(n_1222),
.B1(n_1228),
.B2(n_1163),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1911),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1828),
.Y(n_2084)
);

AOI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1846),
.A2(n_1087),
.B1(n_1094),
.B2(n_1090),
.Y(n_2085)
);

AND2x6_ASAP7_75t_L g2086 ( 
.A(n_1849),
.B(n_1056),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1848),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1845),
.B(n_1434),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1857),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1939),
.B(n_1434),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1989),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1877),
.Y(n_2092)
);

BUFx8_ASAP7_75t_L g2093 ( 
.A(n_1889),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1888),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1989),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1878),
.Y(n_2096)
);

OA21x2_ASAP7_75t_L g2097 ( 
.A1(n_1963),
.A2(n_1321),
.B(n_1320),
.Y(n_2097)
);

INVx5_ASAP7_75t_L g2098 ( 
.A(n_1841),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_2029),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1879),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1841),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1942),
.B(n_1593),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1979),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1997),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1899),
.B(n_1095),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1854),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1856),
.Y(n_2107)
);

OA21x2_ASAP7_75t_L g2108 ( 
.A1(n_1965),
.A2(n_1968),
.B(n_1885),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_1915),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2006),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1980),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1861),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1830),
.B(n_1238),
.Y(n_2113)
);

CKINVDCx20_ASAP7_75t_R g2114 ( 
.A(n_2017),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1831),
.B(n_1238),
.Y(n_2115)
);

INVx4_ASAP7_75t_L g2116 ( 
.A(n_1987),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1996),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1862),
.Y(n_2118)
);

INVx4_ASAP7_75t_L g2119 ( 
.A(n_2016),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1935),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2007),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_2025),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1868),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_1833),
.B(n_1242),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1835),
.B(n_1238),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1836),
.B(n_1238),
.Y(n_2126)
);

INVx5_ASAP7_75t_L g2127 ( 
.A(n_1891),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1969),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1871),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1936),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1843),
.Y(n_2131)
);

CKINVDCx16_ASAP7_75t_R g2132 ( 
.A(n_2055),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_1940),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_2022),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1993),
.Y(n_2135)
);

OA21x2_ASAP7_75t_L g2136 ( 
.A1(n_1883),
.A2(n_1327),
.B(n_1322),
.Y(n_2136)
);

BUFx2_ASAP7_75t_L g2137 ( 
.A(n_1941),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1846),
.B(n_1593),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1998),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_1958),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1839),
.B(n_1238),
.Y(n_2141)
);

CKINVDCx16_ASAP7_75t_R g2142 ( 
.A(n_1834),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1882),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1959),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1884),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_1947),
.A2(n_1096),
.B1(n_1108),
.B2(n_1098),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1886),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1890),
.Y(n_2148)
);

BUFx6f_ASAP7_75t_L g2149 ( 
.A(n_2030),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1949),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1952),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1896),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1962),
.A2(n_1110),
.B1(n_1116),
.B2(n_1114),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1950),
.B(n_1593),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1901),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_2041),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1842),
.B(n_1238),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1903),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_2043),
.Y(n_2159)
);

CKINVDCx20_ASAP7_75t_R g2160 ( 
.A(n_1838),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_1982),
.B(n_1622),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1981),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1983),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2058),
.B(n_2046),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1906),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1907),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1982),
.B(n_1622),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_2047),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_1922),
.A2(n_1118),
.B1(n_1122),
.B2(n_1117),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1910),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_2054),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2042),
.B(n_1622),
.Y(n_2172)
);

BUFx6f_ASAP7_75t_L g2173 ( 
.A(n_1894),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1913),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1984),
.B(n_1251),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_2042),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_1900),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_2001),
.B(n_1123),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1844),
.B(n_1641),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1914),
.Y(n_2180)
);

INVx6_ASAP7_75t_L g2181 ( 
.A(n_1891),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1985),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1986),
.B(n_1251),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_1924),
.A2(n_1127),
.B1(n_1129),
.B2(n_1124),
.Y(n_2184)
);

XNOR2xp5_ASAP7_75t_L g2185 ( 
.A(n_1990),
.B(n_1269),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1988),
.B(n_1251),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1976),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1918),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1919),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1851),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1991),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1992),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1837),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_SL g2194 ( 
.A1(n_2003),
.A2(n_1293),
.B1(n_1309),
.B2(n_1291),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1840),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1994),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1902),
.B(n_1641),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1995),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1999),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_1970),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_2009),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1858),
.Y(n_2202)
);

BUFx3_ASAP7_75t_L g2203 ( 
.A(n_1971),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1909),
.B(n_1310),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_L g2205 ( 
.A1(n_1920),
.A2(n_1071),
.B(n_1058),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2000),
.B(n_1251),
.Y(n_2206)
);

CKINVDCx20_ASAP7_75t_R g2207 ( 
.A(n_2023),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_2033),
.Y(n_2208)
);

AND2x6_ASAP7_75t_L g2209 ( 
.A(n_2004),
.B(n_1058),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1927),
.A2(n_1136),
.B1(n_1137),
.B2(n_1130),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2005),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2010),
.B(n_1251),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1925),
.Y(n_2213)
);

CKINVDCx20_ASAP7_75t_R g2214 ( 
.A(n_2037),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1931),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1932),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_1866),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2011),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2012),
.Y(n_2219)
);

INVx5_ASAP7_75t_L g2220 ( 
.A(n_1891),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_SL g2221 ( 
.A1(n_2040),
.A2(n_1331),
.B1(n_1340),
.B2(n_1328),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_1908),
.B(n_1641),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1933),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2013),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_2045),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1867),
.Y(n_2226)
);

AND2x2_ASAP7_75t_SL g2227 ( 
.A(n_2052),
.B(n_1071),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2015),
.Y(n_2228)
);

CKINVDCx20_ASAP7_75t_R g2229 ( 
.A(n_2059),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2019),
.B(n_1251),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_1912),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1934),
.A2(n_1139),
.B1(n_1141),
.B2(n_1140),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1937),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_1847),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_2002),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_1859),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_1832),
.B(n_1365),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1876),
.A2(n_1145),
.B1(n_1147),
.B2(n_1143),
.Y(n_2238)
);

INVx6_ASAP7_75t_L g2239 ( 
.A(n_1975),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_1872),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1938),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1943),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1945),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1855),
.B(n_1369),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1946),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2024),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_SL g2247 ( 
.A1(n_1923),
.A2(n_1399),
.B1(n_1410),
.B2(n_1392),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_2027),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2031),
.B(n_1251),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1887),
.B(n_1625),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2032),
.B(n_1261),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_1930),
.B(n_1438),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1948),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1874),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1875),
.B(n_1447),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2034),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1881),
.B(n_1472),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_2038),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_2008),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2044),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1954),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1916),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1955),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1863),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_1865),
.B(n_1483),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1978),
.B(n_1149),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1956),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_1904),
.A2(n_1151),
.B1(n_1153),
.B2(n_1152),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2048),
.B(n_1261),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1873),
.B(n_1490),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1957),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2049),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1960),
.Y(n_2273)
);

INVxp67_ASAP7_75t_L g2274 ( 
.A(n_1898),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2026),
.B(n_1091),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2051),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_1892),
.B(n_1508),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2053),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2056),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1897),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2057),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_2060),
.Y(n_2282)
);

OA21x2_ASAP7_75t_L g2283 ( 
.A1(n_1917),
.A2(n_1332),
.B(n_1330),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_1893),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1967),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1944),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_1829),
.B(n_1509),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2035),
.B(n_2036),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1869),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1951),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2028),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1870),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1864),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1926),
.B(n_1261),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1977),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_1972),
.B(n_1261),
.Y(n_2296)
);

OA21x2_ASAP7_75t_L g2297 ( 
.A1(n_1973),
.A2(n_1347),
.B(n_1345),
.Y(n_2297)
);

AND2x6_ASAP7_75t_L g2298 ( 
.A(n_1849),
.B(n_1091),
.Y(n_2298)
);

OAI21x1_ASAP7_75t_L g2299 ( 
.A1(n_1882),
.A2(n_1132),
.B(n_1103),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2014),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2014),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2014),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1989),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2014),
.Y(n_2304)
);

AND2x6_ASAP7_75t_L g2305 ( 
.A(n_1849),
.B(n_1103),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_1964),
.Y(n_2306)
);

INVx3_ASAP7_75t_L g2307 ( 
.A(n_1989),
.Y(n_2307)
);

BUFx3_ASAP7_75t_L g2308 ( 
.A(n_1964),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1860),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1860),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2039),
.B(n_1517),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_1989),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1860),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2014),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_1964),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1860),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1974),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2039),
.B(n_1545),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2014),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2014),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2039),
.B(n_1551),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2014),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2014),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2014),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2020),
.B(n_1428),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_1953),
.B(n_1155),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1974),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2014),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_2039),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1974),
.Y(n_2330)
);

AND2x6_ASAP7_75t_L g2331 ( 
.A(n_1849),
.B(n_1132),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1974),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2014),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2014),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_1860),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1974),
.Y(n_2336)
);

INVx4_ASAP7_75t_L g2337 ( 
.A(n_2039),
.Y(n_2337)
);

CKINVDCx16_ASAP7_75t_R g2338 ( 
.A(n_1997),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2014),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2014),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_SL g2341 ( 
.A1(n_1850),
.A2(n_1603),
.B1(n_1604),
.B2(n_1564),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_1974),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_1964),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2014),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_R g2345 ( 
.A(n_1847),
.B(n_1158),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2014),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_1964),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_1974),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_1860),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2014),
.B(n_1261),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_2039),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2014),
.Y(n_2352)
);

INVx4_ASAP7_75t_L g2353 ( 
.A(n_2039),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1860),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2014),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2020),
.B(n_1428),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2014),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2014),
.B(n_1261),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2020),
.B(n_1159),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2014),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1860),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_1860),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_SL g2363 ( 
.A1(n_1850),
.A2(n_1611),
.B1(n_1642),
.B2(n_1607),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2039),
.B(n_1678),
.Y(n_2364)
);

BUFx6f_ASAP7_75t_L g2365 ( 
.A(n_2039),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_1860),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2014),
.B(n_1261),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2039),
.B(n_1074),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2108),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2108),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_2176),
.B(n_1160),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2136),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2136),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2205),
.Y(n_2374)
);

BUFx3_ASAP7_75t_L g2375 ( 
.A(n_2091),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_2299),
.Y(n_2376)
);

BUFx6f_ASAP7_75t_L g2377 ( 
.A(n_2283),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2143),
.Y(n_2378)
);

NAND3x1_ASAP7_75t_L g2379 ( 
.A(n_2291),
.B(n_1207),
.C(n_1078),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2283),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2087),
.B(n_1211),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2145),
.Y(n_2382)
);

NAND3xp33_ASAP7_75t_L g2383 ( 
.A(n_2071),
.B(n_1162),
.C(n_1161),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2147),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2148),
.Y(n_2385)
);

OAI22xp33_ASAP7_75t_SL g2386 ( 
.A1(n_2066),
.A2(n_1165),
.B1(n_1172),
.B2(n_1164),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2274),
.B(n_1177),
.Y(n_2387)
);

AOI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2288),
.A2(n_1356),
.B(n_1353),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2091),
.B(n_1180),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2152),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_2098),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2155),
.Y(n_2392)
);

OAI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2309),
.A2(n_1503),
.B1(n_1554),
.B2(n_1486),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2158),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2235),
.B(n_1183),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2165),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2166),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2170),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2174),
.Y(n_2399)
);

INVx2_ASAP7_75t_SL g2400 ( 
.A(n_2095),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2180),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2188),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2138),
.B(n_1189),
.Y(n_2403)
);

CKINVDCx6p67_ASAP7_75t_R g2404 ( 
.A(n_2095),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2093),
.Y(n_2405)
);

BUFx10_ASAP7_75t_L g2406 ( 
.A(n_2164),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2189),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2213),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2215),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2140),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2216),
.Y(n_2411)
);

AOI21x1_ASAP7_75t_L g2412 ( 
.A1(n_2078),
.A2(n_1360),
.B(n_1358),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2223),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2109),
.B(n_1154),
.Y(n_2414)
);

INVxp33_ASAP7_75t_L g2415 ( 
.A(n_2094),
.Y(n_2415)
);

INVx5_ASAP7_75t_L g2416 ( 
.A(n_2303),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2081),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2161),
.B(n_1194),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2120),
.B(n_1181),
.Y(n_2419)
);

BUFx3_ASAP7_75t_L g2420 ( 
.A(n_2239),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2233),
.Y(n_2421)
);

BUFx3_ASAP7_75t_L g2422 ( 
.A(n_2239),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2241),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2310),
.Y(n_2424)
);

OR2x2_ASAP7_75t_L g2425 ( 
.A(n_2120),
.B(n_1223),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2242),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2243),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2131),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2074),
.B(n_1195),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2245),
.Y(n_2430)
);

INVx8_ASAP7_75t_L g2431 ( 
.A(n_2064),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2253),
.Y(n_2432)
);

INVx8_ASAP7_75t_L g2433 ( 
.A(n_2064),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2261),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2172),
.B(n_1197),
.Y(n_2435)
);

INVx2_ASAP7_75t_SL g2436 ( 
.A(n_2329),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2077),
.B(n_1199),
.Y(n_2437)
);

NOR2x1p5_ASAP7_75t_L g2438 ( 
.A(n_2313),
.B(n_1200),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2263),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2267),
.Y(n_2440)
);

OR2x6_ASAP7_75t_L g2441 ( 
.A(n_2082),
.B(n_1057),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2316),
.B(n_2335),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2271),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_2259),
.B(n_1208),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2106),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2273),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2259),
.B(n_1209),
.Y(n_2447)
);

INVxp67_ASAP7_75t_L g2448 ( 
.A(n_2236),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2197),
.B(n_1217),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_SL g2450 ( 
.A(n_2306),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2101),
.Y(n_2451)
);

AOI21x1_ASAP7_75t_L g2452 ( 
.A1(n_2080),
.A2(n_2296),
.B(n_2062),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2084),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2089),
.Y(n_2454)
);

NOR2x1p5_ASAP7_75t_L g2455 ( 
.A(n_2349),
.B(n_1220),
.Y(n_2455)
);

NOR2x1p5_ASAP7_75t_L g2456 ( 
.A(n_2354),
.B(n_1224),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2110),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2280),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2307),
.B(n_1225),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2312),
.B(n_1231),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2361),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2290),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2107),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2222),
.B(n_1232),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2112),
.Y(n_2465)
);

INVx2_ASAP7_75t_SL g2466 ( 
.A(n_2329),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2092),
.Y(n_2467)
);

BUFx10_ASAP7_75t_L g2468 ( 
.A(n_2190),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2096),
.Y(n_2469)
);

BUFx2_ASAP7_75t_L g2470 ( 
.A(n_2362),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2097),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2366),
.B(n_2326),
.Y(n_2472)
);

BUFx4f_ASAP7_75t_L g2473 ( 
.A(n_2103),
.Y(n_2473)
);

AND3x2_ASAP7_75t_L g2474 ( 
.A(n_2130),
.B(n_1367),
.C(n_1362),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2100),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2097),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2262),
.B(n_1237),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2262),
.B(n_1239),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2113),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2118),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2130),
.B(n_1277),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2123),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2128),
.Y(n_2483)
);

BUFx6f_ASAP7_75t_L g2484 ( 
.A(n_2099),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2129),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2150),
.B(n_1240),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2067),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2266),
.B(n_1244),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2063),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2293),
.B(n_1249),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2068),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2098),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2359),
.B(n_1252),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2137),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2300),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2317),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2179),
.B(n_1255),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2301),
.Y(n_2498)
);

BUFx2_ASAP7_75t_L g2499 ( 
.A(n_2133),
.Y(n_2499)
);

INVx2_ASAP7_75t_SL g2500 ( 
.A(n_2351),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2327),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2151),
.B(n_1260),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2289),
.B(n_1262),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2330),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2332),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2302),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2304),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2336),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_SL g2509 ( 
.A(n_2264),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2342),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2314),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2098),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2167),
.B(n_1263),
.Y(n_2513)
);

BUFx10_ASAP7_75t_L g2514 ( 
.A(n_2190),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2319),
.Y(n_2515)
);

INVx1_ASAP7_75t_SL g2516 ( 
.A(n_2200),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2320),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_L g2518 ( 
.A(n_2086),
.B(n_1553),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2348),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2115),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2204),
.B(n_1264),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2322),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2323),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2248),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2070),
.B(n_1265),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2258),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2324),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2250),
.B(n_1266),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2282),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2292),
.B(n_1267),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2069),
.B(n_1270),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2297),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2125),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2073),
.B(n_1274),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2126),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2297),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_2088),
.B(n_1278),
.Y(n_2537)
);

BUFx3_ASAP7_75t_L g2538 ( 
.A(n_2351),
.Y(n_2538)
);

INVx2_ASAP7_75t_SL g2539 ( 
.A(n_2365),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2141),
.Y(n_2540)
);

INVx3_ASAP7_75t_L g2541 ( 
.A(n_2099),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2157),
.Y(n_2542)
);

INVx3_ASAP7_75t_L g2543 ( 
.A(n_2121),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2328),
.B(n_1280),
.Y(n_2544)
);

INVxp33_ASAP7_75t_L g2545 ( 
.A(n_2185),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2333),
.B(n_1284),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_2173),
.B(n_1285),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2175),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2183),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2334),
.Y(n_2550)
);

INVxp67_ASAP7_75t_R g2551 ( 
.A(n_2247),
.Y(n_2551)
);

INVx3_ASAP7_75t_L g2552 ( 
.A(n_2339),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2144),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2340),
.B(n_1289),
.Y(n_2554)
);

AOI21x1_ASAP7_75t_L g2555 ( 
.A1(n_2061),
.A2(n_1376),
.B(n_1375),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2344),
.B(n_1290),
.Y(n_2556)
);

INVxp67_ASAP7_75t_SL g2557 ( 
.A(n_2203),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2346),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2186),
.Y(n_2559)
);

INVx2_ASAP7_75t_SL g2560 ( 
.A(n_2365),
.Y(n_2560)
);

AND3x2_ASAP7_75t_L g2561 ( 
.A(n_2177),
.B(n_1386),
.C(n_1383),
.Y(n_2561)
);

INVx3_ASAP7_75t_L g2562 ( 
.A(n_2352),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2355),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2206),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_SL g2565 ( 
.A(n_2308),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2357),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2212),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2230),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2090),
.B(n_1294),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2360),
.Y(n_2570)
);

CKINVDCx6p67_ASAP7_75t_R g2571 ( 
.A(n_2132),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2162),
.Y(n_2572)
);

CKINVDCx20_ASAP7_75t_R g2573 ( 
.A(n_2160),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2163),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2182),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2191),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2249),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2192),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2251),
.Y(n_2579)
);

CKINVDCx6p67_ASAP7_75t_R g2580 ( 
.A(n_2338),
.Y(n_2580)
);

BUFx6f_ASAP7_75t_L g2581 ( 
.A(n_2127),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2196),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2065),
.B(n_1295),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2269),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2198),
.Y(n_2585)
);

INVxp33_ASAP7_75t_L g2586 ( 
.A(n_2185),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2178),
.B(n_1296),
.Y(n_2587)
);

AND3x2_ASAP7_75t_L g2588 ( 
.A(n_2265),
.B(n_1402),
.C(n_1387),
.Y(n_2588)
);

BUFx8_ASAP7_75t_SL g2589 ( 
.A(n_2201),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2199),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2127),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2350),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2211),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2358),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2173),
.B(n_1304),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2218),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2169),
.B(n_1305),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2367),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2076),
.Y(n_2599)
);

XOR2x2_ASAP7_75t_L g2600 ( 
.A(n_2075),
.B(n_1),
.Y(n_2600)
);

INVxp67_ASAP7_75t_SL g2601 ( 
.A(n_2268),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2219),
.Y(n_2602)
);

BUFx3_ASAP7_75t_L g2603 ( 
.A(n_2103),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2224),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2086),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2228),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2246),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2256),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2086),
.B(n_1313),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2260),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2298),
.B(n_2305),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2272),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2127),
.Y(n_2613)
);

INVx4_ASAP7_75t_L g2614 ( 
.A(n_2337),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2276),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2278),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2353),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2279),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2281),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2135),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2232),
.A2(n_1319),
.B1(n_1323),
.B2(n_1315),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2146),
.B(n_2153),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2285),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2139),
.Y(n_2624)
);

INVx5_ASAP7_75t_L g2625 ( 
.A(n_2187),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2298),
.B(n_1324),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2220),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2220),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2220),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2181),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2181),
.Y(n_2631)
);

BUFx10_ASAP7_75t_L g2632 ( 
.A(n_2202),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2286),
.Y(n_2633)
);

INVx2_ASAP7_75t_SL g2634 ( 
.A(n_2187),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2298),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2275),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2305),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2305),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2331),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2227),
.B(n_1325),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2331),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2085),
.B(n_1329),
.Y(n_2642)
);

OAI22xp5_ASAP7_75t_SL g2643 ( 
.A1(n_2341),
.A2(n_1334),
.B1(n_1335),
.B2(n_1333),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2331),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2209),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2209),
.B(n_1336),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2209),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2294),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2102),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2154),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2184),
.B(n_1337),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2238),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2210),
.B(n_1338),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_2105),
.B(n_1342),
.Y(n_2654)
);

INVx5_ASAP7_75t_L g2655 ( 
.A(n_2231),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2202),
.B(n_1343),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2287),
.B(n_1344),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2217),
.Y(n_2658)
);

INVx2_ASAP7_75t_SL g2659 ( 
.A(n_2079),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2325),
.Y(n_2660)
);

AO21x2_ASAP7_75t_L g2661 ( 
.A1(n_2237),
.A2(n_1415),
.B(n_1411),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2356),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2244),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2295),
.Y(n_2664)
);

NAND3xp33_ASAP7_75t_L g2665 ( 
.A(n_2345),
.B(n_1348),
.C(n_1346),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2134),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2156),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2072),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2116),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2072),
.Y(n_2670)
);

CKINVDCx6p67_ASAP7_75t_R g2671 ( 
.A(n_2142),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_L g2672 ( 
.A(n_2311),
.B(n_1350),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2119),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2347),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2347),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_2318),
.B(n_1351),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2284),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2284),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2217),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2111),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2111),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2226),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2117),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2117),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2226),
.Y(n_2685)
);

INVx1_ASAP7_75t_SL g2686 ( 
.A(n_2315),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2240),
.B(n_1352),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_L g2688 ( 
.A(n_2321),
.B(n_1354),
.Y(n_2688)
);

INVx3_ASAP7_75t_L g2689 ( 
.A(n_2149),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2149),
.Y(n_2690)
);

NAND3xp33_ASAP7_75t_L g2691 ( 
.A(n_2254),
.B(n_1364),
.C(n_1363),
.Y(n_2691)
);

AND3x2_ASAP7_75t_L g2692 ( 
.A(n_2270),
.B(n_1425),
.C(n_1420),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2193),
.A2(n_1368),
.B1(n_1373),
.B2(n_1366),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2159),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2159),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2343),
.Y(n_2696)
);

INVxp33_ASAP7_75t_SL g2697 ( 
.A(n_2083),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2124),
.Y(n_2698)
);

BUFx10_ASAP7_75t_L g2699 ( 
.A(n_2104),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2364),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2195),
.B(n_1378),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2368),
.Y(n_2702)
);

INVx3_ASAP7_75t_L g2703 ( 
.A(n_2168),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2255),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2257),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2363),
.B(n_1341),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2122),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2252),
.B(n_1379),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2234),
.B(n_1380),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2194),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2171),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2277),
.B(n_1384),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2114),
.Y(n_2713)
);

OAI22xp33_ASAP7_75t_SL g2714 ( 
.A1(n_2208),
.A2(n_1388),
.B1(n_1389),
.B2(n_1385),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2221),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2225),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2207),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2214),
.B(n_1390),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2229),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2108),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2108),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2081),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2081),
.Y(n_2723)
);

OR2x2_ASAP7_75t_L g2724 ( 
.A(n_2087),
.B(n_1349),
.Y(n_2724)
);

INVx2_ASAP7_75t_SL g2725 ( 
.A(n_2087),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2108),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2108),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2108),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2087),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2176),
.B(n_1391),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2108),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2138),
.B(n_1393),
.Y(n_2732)
);

AOI21x1_ASAP7_75t_L g2733 ( 
.A1(n_2288),
.A2(n_1459),
.B(n_1446),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2087),
.B(n_1394),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2108),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2108),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2108),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2087),
.Y(n_2738)
);

AOI21x1_ASAP7_75t_L g2739 ( 
.A1(n_2288),
.A2(n_1463),
.B(n_1460),
.Y(n_2739)
);

BUFx6f_ASAP7_75t_L g2740 ( 
.A(n_2108),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2108),
.Y(n_2741)
);

AOI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2176),
.A2(n_1397),
.B1(n_1398),
.B2(n_1395),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2108),
.Y(n_2743)
);

NOR2x1p5_ASAP7_75t_L g2744 ( 
.A(n_2066),
.B(n_1400),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2091),
.B(n_1404),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2108),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2108),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2108),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2108),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2108),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2108),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_2091),
.B(n_1405),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2176),
.B(n_1407),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2108),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_2176),
.B(n_1408),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2176),
.B(n_1409),
.Y(n_2756)
);

NAND2xp33_ASAP7_75t_SL g2757 ( 
.A(n_2091),
.B(n_1413),
.Y(n_2757)
);

INVx8_ASAP7_75t_L g2758 ( 
.A(n_2091),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2108),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2087),
.B(n_1355),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_SL g2761 ( 
.A(n_2091),
.B(n_1417),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2108),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2138),
.B(n_1418),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2415),
.B(n_1421),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2417),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2731),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2731),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2428),
.Y(n_2768)
);

INVx2_ASAP7_75t_SL g2769 ( 
.A(n_2758),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2734),
.B(n_1422),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2735),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2445),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2463),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2652),
.B(n_1423),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_2589),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_L g2776 ( 
.A(n_2448),
.B(n_1424),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2465),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2735),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2729),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_2738),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2740),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2736),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2480),
.Y(n_2783)
);

BUFx6f_ASAP7_75t_L g2784 ( 
.A(n_2740),
.Y(n_2784)
);

INVx4_ASAP7_75t_L g2785 ( 
.A(n_2758),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2736),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2467),
.B(n_1427),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2467),
.B(n_1429),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2737),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2482),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2485),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2737),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2743),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2743),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2747),
.Y(n_2795)
);

INVx1_ASAP7_75t_SL g2796 ( 
.A(n_2410),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2686),
.B(n_1430),
.Y(n_2797)
);

INVx4_ASAP7_75t_L g2798 ( 
.A(n_2404),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2747),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2725),
.B(n_1432),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2431),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2748),
.Y(n_2802)
);

INVx3_ASAP7_75t_L g2803 ( 
.A(n_2581),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2748),
.Y(n_2804)
);

INVx3_ASAP7_75t_L g2805 ( 
.A(n_2581),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2750),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2722),
.Y(n_2807)
);

OR2x6_ASAP7_75t_L g2808 ( 
.A(n_2405),
.B(n_1106),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2750),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2700),
.B(n_1433),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2751),
.A2(n_1437),
.B1(n_1439),
.B2(n_1436),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2723),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2751),
.Y(n_2813)
);

AND2x6_ASAP7_75t_L g2814 ( 
.A(n_2635),
.B(n_1157),
.Y(n_2814)
);

AND2x6_ASAP7_75t_L g2815 ( 
.A(n_2635),
.B(n_1157),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2724),
.B(n_2760),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2698),
.B(n_1440),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2712),
.B(n_1441),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2469),
.B(n_2475),
.Y(n_2819)
);

OR2x2_ASAP7_75t_L g2820 ( 
.A(n_2414),
.B(n_1374),
.Y(n_2820)
);

INVx5_ASAP7_75t_L g2821 ( 
.A(n_2658),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_2571),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2469),
.B(n_2475),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2572),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2635),
.B(n_1442),
.Y(n_2825)
);

AOI22xp33_ASAP7_75t_L g2826 ( 
.A1(n_2715),
.A2(n_1448),
.B1(n_1450),
.B2(n_1449),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2494),
.Y(n_2827)
);

CKINVDCx16_ASAP7_75t_R g2828 ( 
.A(n_2573),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2369),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2370),
.Y(n_2830)
);

INVx8_ASAP7_75t_L g2831 ( 
.A(n_2431),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2576),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2602),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2381),
.B(n_1452),
.Y(n_2834)
);

INVxp67_ASAP7_75t_SL g2835 ( 
.A(n_2740),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2604),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2614),
.B(n_1080),
.Y(n_2837)
);

INVx6_ASAP7_75t_L g2838 ( 
.A(n_2468),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2607),
.Y(n_2839)
);

INVx4_ASAP7_75t_L g2840 ( 
.A(n_2433),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2493),
.B(n_1453),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_2614),
.B(n_1456),
.Y(n_2842)
);

AND2x4_ASAP7_75t_L g2843 ( 
.A(n_2655),
.B(n_1107),
.Y(n_2843)
);

NAND3xp33_ASAP7_75t_L g2844 ( 
.A(n_2654),
.B(n_1691),
.C(n_1690),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2655),
.B(n_1111),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2597),
.B(n_1457),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2612),
.B(n_1458),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2720),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2581),
.Y(n_2849)
);

INVx1_ASAP7_75t_SL g2850 ( 
.A(n_2433),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2591),
.Y(n_2851)
);

BUFx2_ASAP7_75t_L g2852 ( 
.A(n_2499),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_2658),
.B(n_1462),
.Y(n_2853)
);

OR2x6_ASAP7_75t_L g2854 ( 
.A(n_2441),
.B(n_1106),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_L g2855 ( 
.A(n_2591),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2580),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2615),
.Y(n_2857)
);

BUFx6f_ASAP7_75t_L g2858 ( 
.A(n_2591),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2616),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2574),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2575),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2704),
.B(n_2705),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2710),
.A2(n_1465),
.B1(n_1467),
.B2(n_1464),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2655),
.B(n_1214),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2721),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2468),
.Y(n_2866)
);

AND2x6_ASAP7_75t_L g2867 ( 
.A(n_2605),
.B(n_1157),
.Y(n_2867)
);

INVx1_ASAP7_75t_SL g2868 ( 
.A(n_2375),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_2658),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2387),
.B(n_1469),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2578),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2726),
.Y(n_2872)
);

BUFx10_ASAP7_75t_L g2873 ( 
.A(n_2450),
.Y(n_2873)
);

AND2x6_ASAP7_75t_L g2874 ( 
.A(n_2605),
.B(n_1157),
.Y(n_2874)
);

INVxp67_ASAP7_75t_SL g2875 ( 
.A(n_2727),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2671),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2582),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2585),
.Y(n_2878)
);

AND2x4_ASAP7_75t_L g2879 ( 
.A(n_2416),
.B(n_1236),
.Y(n_2879)
);

INVx4_ASAP7_75t_L g2880 ( 
.A(n_2625),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2590),
.Y(n_2881)
);

BUFx3_ASAP7_75t_L g2882 ( 
.A(n_2625),
.Y(n_2882)
);

AND2x6_ASAP7_75t_L g2883 ( 
.A(n_2372),
.B(n_1169),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2651),
.B(n_1471),
.Y(n_2884)
);

AND2x2_ASAP7_75t_SL g2885 ( 
.A(n_2473),
.B(n_2706),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2728),
.Y(n_2886)
);

OAI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2741),
.A2(n_1477),
.B1(n_1478),
.B2(n_1473),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2702),
.B(n_2622),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2746),
.Y(n_2889)
);

AND2x6_ASAP7_75t_L g2890 ( 
.A(n_2372),
.B(n_1169),
.Y(n_2890)
);

BUFx3_ASAP7_75t_L g2891 ( 
.A(n_2625),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2488),
.B(n_1480),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2416),
.B(n_1254),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2749),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2593),
.B(n_1484),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2596),
.B(n_1487),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2640),
.B(n_1488),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2606),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2416),
.B(n_1491),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2754),
.Y(n_2900)
);

AND2x6_ASAP7_75t_L g2901 ( 
.A(n_2373),
.B(n_2380),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2583),
.B(n_1496),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2528),
.B(n_1497),
.Y(n_2903)
);

INVx2_ASAP7_75t_SL g2904 ( 
.A(n_2514),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2608),
.Y(n_2905)
);

AND2x4_ASAP7_75t_L g2906 ( 
.A(n_2617),
.B(n_1273),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2759),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2742),
.B(n_2395),
.Y(n_2908)
);

HB1xp67_ASAP7_75t_L g2909 ( 
.A(n_2553),
.Y(n_2909)
);

BUFx3_ASAP7_75t_L g2910 ( 
.A(n_2514),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2610),
.Y(n_2911)
);

BUFx4f_ASAP7_75t_L g2912 ( 
.A(n_2441),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2762),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_2419),
.B(n_1656),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2618),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2619),
.B(n_1498),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2719),
.B(n_1500),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2392),
.Y(n_2918)
);

NAND2x1_ASAP7_75t_L g2919 ( 
.A(n_2613),
.B(n_1169),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2392),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_2400),
.B(n_1275),
.Y(n_2921)
);

BUFx6f_ASAP7_75t_L g2922 ( 
.A(n_2613),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2601),
.B(n_1504),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2397),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2397),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2399),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2524),
.B(n_1401),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2399),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2552),
.Y(n_2929)
);

AOI22xp33_ASAP7_75t_L g2930 ( 
.A1(n_2657),
.A2(n_1512),
.B1(n_1513),
.B2(n_1505),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2371),
.B(n_1521),
.Y(n_2931)
);

NAND3xp33_ASAP7_75t_L g2932 ( 
.A(n_2521),
.B(n_1675),
.C(n_1674),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2730),
.B(n_1522),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2552),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2401),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2487),
.B(n_1524),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_L g2937 ( 
.A(n_2660),
.B(n_1525),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2662),
.B(n_1529),
.Y(n_2938)
);

CKINVDCx5p33_ASAP7_75t_R g2939 ( 
.A(n_2509),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2538),
.Y(n_2940)
);

BUFx3_ASAP7_75t_L g2941 ( 
.A(n_2632),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2753),
.B(n_2755),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2401),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2409),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2562),
.Y(n_2945)
);

BUFx10_ASAP7_75t_L g2946 ( 
.A(n_2450),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2621),
.B(n_1532),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2693),
.B(n_2756),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2409),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2562),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2491),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2472),
.B(n_1535),
.Y(n_2952)
);

OR2x2_ASAP7_75t_L g2953 ( 
.A(n_2425),
.B(n_1396),
.Y(n_2953)
);

OR2x2_ASAP7_75t_L g2954 ( 
.A(n_2481),
.B(n_1673),
.Y(n_2954)
);

AND2x6_ASAP7_75t_L g2955 ( 
.A(n_2373),
.B(n_1169),
.Y(n_2955)
);

BUFx6f_ASAP7_75t_L g2956 ( 
.A(n_2613),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2526),
.B(n_1406),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2484),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2495),
.B(n_1536),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_L g2960 ( 
.A(n_2497),
.B(n_1537),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2377),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2498),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2377),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2506),
.B(n_1541),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2377),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2393),
.B(n_1454),
.Y(n_2966)
);

AND2x6_ASAP7_75t_L g2967 ( 
.A(n_2380),
.B(n_1202),
.Y(n_2967)
);

AND2x4_ASAP7_75t_L g2968 ( 
.A(n_2529),
.B(n_1451),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2672),
.B(n_1544),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2550),
.Y(n_2970)
);

AND2x6_ASAP7_75t_L g2971 ( 
.A(n_2637),
.B(n_1202),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2507),
.Y(n_2972)
);

INVx2_ASAP7_75t_SL g2973 ( 
.A(n_2632),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2511),
.B(n_1548),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2418),
.B(n_1552),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2515),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2484),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2558),
.Y(n_2978)
);

OAI22xp5_ASAP7_75t_L g2979 ( 
.A1(n_2592),
.A2(n_1557),
.B1(n_1560),
.B2(n_1556),
.Y(n_2979)
);

AND2x6_ASAP7_75t_L g2980 ( 
.A(n_2638),
.B(n_1202),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2563),
.Y(n_2981)
);

INVx3_ASAP7_75t_L g2982 ( 
.A(n_2484),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2517),
.B(n_1562),
.Y(n_2983)
);

INVx4_ASAP7_75t_L g2984 ( 
.A(n_2473),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_2676),
.B(n_1565),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2522),
.B(n_1569),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2523),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2391),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2566),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2527),
.B(n_1570),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2391),
.Y(n_2991)
);

AO22x2_ASAP7_75t_L g2992 ( 
.A1(n_2471),
.A2(n_1561),
.B1(n_1680),
.B2(n_1583),
.Y(n_2992)
);

NOR2xp33_ASAP7_75t_L g2993 ( 
.A(n_2688),
.B(n_1571),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2633),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2435),
.B(n_1572),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2403),
.B(n_1574),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2570),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2378),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2763),
.B(n_2732),
.Y(n_2999)
);

INVx1_ASAP7_75t_SL g3000 ( 
.A(n_2516),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2661),
.B(n_1578),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2376),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2429),
.B(n_1584),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2382),
.Y(n_3004)
);

AND2x4_ASAP7_75t_L g3005 ( 
.A(n_2669),
.B(n_1492),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2384),
.Y(n_3006)
);

INVx4_ASAP7_75t_L g3007 ( 
.A(n_2603),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2673),
.B(n_1546),
.Y(n_3008)
);

INVx3_ASAP7_75t_L g3009 ( 
.A(n_2492),
.Y(n_3009)
);

BUFx4f_ASAP7_75t_L g3010 ( 
.A(n_2703),
.Y(n_3010)
);

AND2x6_ASAP7_75t_L g3011 ( 
.A(n_2639),
.B(n_2641),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2649),
.B(n_1549),
.Y(n_3012)
);

AOI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_2668),
.A2(n_1587),
.B1(n_1590),
.B2(n_1585),
.Y(n_3013)
);

BUFx6f_ASAP7_75t_L g3014 ( 
.A(n_2376),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_2697),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2659),
.B(n_1592),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2696),
.B(n_1594),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2437),
.B(n_1595),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2385),
.Y(n_3019)
);

NAND2x1p5_ASAP7_75t_L g3020 ( 
.A(n_2420),
.B(n_1540),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2490),
.B(n_1597),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2449),
.B(n_1601),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2390),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2394),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2396),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_L g3026 ( 
.A(n_2376),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2398),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2670),
.B(n_1602),
.Y(n_3028)
);

BUFx3_ASAP7_75t_L g3029 ( 
.A(n_2422),
.Y(n_3029)
);

CKINVDCx5p33_ASAP7_75t_R g3030 ( 
.A(n_2565),
.Y(n_3030)
);

OR2x6_ASAP7_75t_L g3031 ( 
.A(n_2379),
.B(n_1431),
.Y(n_3031)
);

INVx3_ASAP7_75t_L g3032 ( 
.A(n_2492),
.Y(n_3032)
);

INVx3_ASAP7_75t_L g3033 ( 
.A(n_2512),
.Y(n_3033)
);

CKINVDCx5p33_ASAP7_75t_R g3034 ( 
.A(n_2565),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2402),
.Y(n_3035)
);

AND2x6_ASAP7_75t_L g3036 ( 
.A(n_2645),
.B(n_2647),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2674),
.B(n_1612),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_2386),
.B(n_2461),
.Y(n_3038)
);

AND2x6_ASAP7_75t_L g3039 ( 
.A(n_2644),
.B(n_1202),
.Y(n_3039)
);

INVx3_ASAP7_75t_L g3040 ( 
.A(n_2512),
.Y(n_3040)
);

BUFx8_ASAP7_75t_SL g3041 ( 
.A(n_2424),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2464),
.B(n_1616),
.Y(n_3042)
);

INVx3_ASAP7_75t_L g3043 ( 
.A(n_2541),
.Y(n_3043)
);

INVx4_ASAP7_75t_L g3044 ( 
.A(n_2406),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2503),
.B(n_1617),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2407),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2408),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2411),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_2699),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2413),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2530),
.B(n_2544),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2442),
.B(n_1623),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2675),
.B(n_1624),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2421),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_2663),
.B(n_1628),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2423),
.Y(n_3056)
);

AND2x4_ASAP7_75t_L g3057 ( 
.A(n_2678),
.B(n_1573),
.Y(n_3057)
);

BUFx3_ASAP7_75t_L g3058 ( 
.A(n_2689),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2426),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2427),
.Y(n_3060)
);

AND3x4_ASAP7_75t_L g3061 ( 
.A(n_2713),
.B(n_1218),
.C(n_1204),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2406),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2643),
.A2(n_1634),
.B1(n_1636),
.B2(n_1630),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2646),
.B(n_1639),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2537),
.B(n_1643),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2430),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2699),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2546),
.B(n_1644),
.Y(n_3068)
);

INVxp33_ASAP7_75t_L g3069 ( 
.A(n_2470),
.Y(n_3069)
);

BUFx6f_ASAP7_75t_L g3070 ( 
.A(n_2476),
.Y(n_3070)
);

INVxp67_ASAP7_75t_SL g3071 ( 
.A(n_2703),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2708),
.B(n_1648),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2717),
.B(n_2653),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2532),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2554),
.B(n_1649),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2432),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2556),
.B(n_1651),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_2689),
.B(n_1582),
.Y(n_3078)
);

AND2x2_ASAP7_75t_L g3079 ( 
.A(n_2551),
.B(n_1652),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_2436),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_2541),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2434),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2438),
.B(n_2455),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2439),
.Y(n_3084)
);

HB1xp67_ASAP7_75t_L g3085 ( 
.A(n_2466),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_SL g3086 ( 
.A(n_2600),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2634),
.B(n_2680),
.Y(n_3087)
);

INVx2_ASAP7_75t_SL g3088 ( 
.A(n_2500),
.Y(n_3088)
);

INVx4_ASAP7_75t_L g3089 ( 
.A(n_2561),
.Y(n_3089)
);

INVx1_ASAP7_75t_SL g3090 ( 
.A(n_2757),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2456),
.B(n_1654),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2440),
.Y(n_3092)
);

AND2x6_ASAP7_75t_L g3093 ( 
.A(n_2592),
.B(n_2594),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_2536),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2443),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2744),
.B(n_1655),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2446),
.Y(n_3097)
);

INVx2_ASAP7_75t_SL g3098 ( 
.A(n_2539),
.Y(n_3098)
);

INVx2_ASAP7_75t_SL g3099 ( 
.A(n_2560),
.Y(n_3099)
);

OAI21xp33_ASAP7_75t_SL g3100 ( 
.A1(n_2479),
.A2(n_1683),
.B(n_1679),
.Y(n_3100)
);

XNOR2xp5_ASAP7_75t_L g3101 ( 
.A(n_2545),
.B(n_1659),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2489),
.B(n_1660),
.Y(n_3102)
);

AOI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_2711),
.A2(n_1663),
.B1(n_1664),
.B2(n_1662),
.Y(n_3103)
);

BUFx3_ASAP7_75t_L g3104 ( 
.A(n_2681),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2496),
.Y(n_3105)
);

AND2x6_ASAP7_75t_L g3106 ( 
.A(n_2594),
.B(n_1210),
.Y(n_3106)
);

HB1xp67_ASAP7_75t_L g3107 ( 
.A(n_2557),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2501),
.B(n_2504),
.Y(n_3108)
);

AND2x4_ASAP7_75t_L g3109 ( 
.A(n_2683),
.B(n_1204),
.Y(n_3109)
);

AND2x2_ASAP7_75t_SL g3110 ( 
.A(n_2518),
.B(n_1135),
.Y(n_3110)
);

INVx4_ASAP7_75t_L g3111 ( 
.A(n_2474),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2505),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2508),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_L g3114 ( 
.A(n_2707),
.B(n_1665),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2609),
.B(n_2626),
.Y(n_3115)
);

AND2x4_ASAP7_75t_L g3116 ( 
.A(n_2684),
.B(n_1218),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2510),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2519),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2587),
.B(n_1666),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2388),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2733),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2716),
.B(n_1667),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2664),
.B(n_1670),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2739),
.Y(n_3124)
);

INVx5_ASAP7_75t_L g3125 ( 
.A(n_2543),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2458),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2462),
.Y(n_3127)
);

AND2x6_ASAP7_75t_L g3128 ( 
.A(n_2598),
.B(n_1210),
.Y(n_3128)
);

OR2x2_ASAP7_75t_L g3129 ( 
.A(n_2586),
.B(n_1671),
.Y(n_3129)
);

BUFx3_ASAP7_75t_L g3130 ( 
.A(n_2690),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2453),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_2665),
.B(n_1672),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2451),
.Y(n_3133)
);

OR2x6_ASAP7_75t_L g3134 ( 
.A(n_2694),
.B(n_2695),
.Y(n_3134)
);

AND2x6_ASAP7_75t_L g3135 ( 
.A(n_2598),
.B(n_1210),
.Y(n_3135)
);

INVx4_ASAP7_75t_L g3136 ( 
.A(n_2588),
.Y(n_3136)
);

AOI22xp33_ASAP7_75t_L g3137 ( 
.A1(n_2599),
.A2(n_1676),
.B1(n_1685),
.B2(n_1684),
.Y(n_3137)
);

AND2x2_ASAP7_75t_SL g3138 ( 
.A(n_2611),
.B(n_2677),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2691),
.B(n_1686),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2513),
.B(n_1687),
.Y(n_3140)
);

INVx2_ASAP7_75t_SL g3141 ( 
.A(n_2666),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2454),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_2642),
.B(n_1086),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_2718),
.B(n_1576),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2457),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2636),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2620),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2555),
.Y(n_3148)
);

INVx4_ASAP7_75t_L g3149 ( 
.A(n_2692),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2623),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2531),
.B(n_1092),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2534),
.B(n_1099),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2648),
.B(n_1468),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2569),
.B(n_1112),
.Y(n_3154)
);

INVx4_ASAP7_75t_L g3155 ( 
.A(n_2543),
.Y(n_3155)
);

BUFx10_ASAP7_75t_L g3156 ( 
.A(n_2679),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2714),
.B(n_1637),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2412),
.Y(n_3158)
);

AND2x6_ASAP7_75t_L g3159 ( 
.A(n_2599),
.B(n_1210),
.Y(n_3159)
);

INVx3_ASAP7_75t_L g3160 ( 
.A(n_2627),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2624),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2483),
.Y(n_3162)
);

BUFx6f_ASAP7_75t_L g3163 ( 
.A(n_2374),
.Y(n_3163)
);

NAND2xp33_ASAP7_75t_R g3164 ( 
.A(n_2682),
.B(n_1),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2650),
.B(n_1470),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2479),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_2383),
.B(n_1125),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_SL g3168 ( 
.A(n_2667),
.B(n_1682),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2520),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_2685),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2477),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2520),
.Y(n_3172)
);

INVx2_ASAP7_75t_SL g3173 ( 
.A(n_2389),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2478),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2533),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2533),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2535),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_2628),
.Y(n_3178)
);

NAND2x1p5_ASAP7_75t_L g3179 ( 
.A(n_2525),
.B(n_1461),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2444),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_2629),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2447),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2535),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2540),
.B(n_1474),
.Y(n_3184)
);

AND2x6_ASAP7_75t_L g3185 ( 
.A(n_2540),
.B(n_1271),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2542),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2542),
.Y(n_3187)
);

INVxp33_ASAP7_75t_L g3188 ( 
.A(n_2687),
.Y(n_3188)
);

INVx5_ASAP7_75t_L g3189 ( 
.A(n_2630),
.Y(n_3189)
);

NAND2xp33_ASAP7_75t_L g3190 ( 
.A(n_2548),
.B(n_1553),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2486),
.B(n_1126),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2701),
.B(n_1128),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2548),
.Y(n_3193)
);

CKINVDCx5p33_ASAP7_75t_R g3194 ( 
.A(n_2709),
.Y(n_3194)
);

AND2x4_ASAP7_75t_SL g3195 ( 
.A(n_2549),
.B(n_1271),
.Y(n_3195)
);

INVxp33_ASAP7_75t_L g3196 ( 
.A(n_2656),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_L g3197 ( 
.A(n_2631),
.Y(n_3197)
);

INVx5_ASAP7_75t_L g3198 ( 
.A(n_2745),
.Y(n_3198)
);

INVx4_ASAP7_75t_L g3199 ( 
.A(n_2549),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_2502),
.B(n_1138),
.Y(n_3200)
);

BUFx10_ASAP7_75t_L g3201 ( 
.A(n_2559),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2559),
.B(n_2564),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2564),
.B(n_2567),
.Y(n_3203)
);

INVx4_ASAP7_75t_L g3204 ( 
.A(n_2567),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2568),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2568),
.Y(n_3206)
);

AND2x4_ASAP7_75t_L g3207 ( 
.A(n_2547),
.B(n_1461),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2577),
.Y(n_3208)
);

OR2x2_ASAP7_75t_L g3209 ( 
.A(n_2752),
.B(n_2761),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_SL g3210 ( 
.A(n_2577),
.B(n_1144),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_2459),
.B(n_1150),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2579),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_2579),
.B(n_2584),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_2584),
.B(n_1168),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_2460),
.Y(n_3215)
);

CKINVDCx20_ASAP7_75t_R g3216 ( 
.A(n_2595),
.Y(n_3216)
);

NAND3xp33_ASAP7_75t_L g3217 ( 
.A(n_2452),
.B(n_1272),
.C(n_1271),
.Y(n_3217)
);

HB1xp67_ASAP7_75t_L g3218 ( 
.A(n_2729),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2417),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2417),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2731),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2652),
.B(n_1476),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2652),
.B(n_1481),
.Y(n_3223)
);

INVx1_ASAP7_75t_SL g3224 ( 
.A(n_2729),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2417),
.Y(n_3225)
);

INVxp67_ASAP7_75t_L g3226 ( 
.A(n_2725),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2652),
.B(n_1489),
.Y(n_3227)
);

INVxp33_ASAP7_75t_L g3228 ( 
.A(n_2381),
.Y(n_3228)
);

NOR2xp67_ASAP7_75t_L g3229 ( 
.A(n_2614),
.B(n_2),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2417),
.Y(n_3230)
);

BUFx6f_ASAP7_75t_L g3231 ( 
.A(n_2740),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2417),
.Y(n_3232)
);

INVx4_ASAP7_75t_L g3233 ( 
.A(n_2758),
.Y(n_3233)
);

INVx1_ASAP7_75t_SL g3234 ( 
.A(n_2729),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_2731),
.Y(n_3235)
);

INVx4_ASAP7_75t_L g3236 ( 
.A(n_2758),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2652),
.B(n_1493),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2758),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2417),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2731),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2740),
.Y(n_3241)
);

OR2x2_ASAP7_75t_L g3242 ( 
.A(n_2724),
.B(n_1175),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2581),
.Y(n_3243)
);

BUFx6f_ASAP7_75t_L g3244 ( 
.A(n_2740),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2731),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2417),
.Y(n_3246)
);

BUFx6f_ASAP7_75t_L g3247 ( 
.A(n_2740),
.Y(n_3247)
);

INVx5_ASAP7_75t_L g3248 ( 
.A(n_2758),
.Y(n_3248)
);

INVxp67_ASAP7_75t_L g3249 ( 
.A(n_2725),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_2614),
.B(n_1494),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2731),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_2415),
.B(n_1176),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2734),
.B(n_1205),
.Y(n_3253)
);

NAND2x1p5_ASAP7_75t_L g3254 ( 
.A(n_2375),
.B(n_1271),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_2415),
.B(n_1219),
.Y(n_3255)
);

BUFx8_ASAP7_75t_SL g3256 ( 
.A(n_2589),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2417),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2652),
.B(n_1495),
.Y(n_3258)
);

NOR2xp33_ASAP7_75t_L g3259 ( 
.A(n_2415),
.B(n_1235),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2415),
.B(n_1258),
.Y(n_3260)
);

BUFx10_ASAP7_75t_L g3261 ( 
.A(n_2658),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2734),
.B(n_1268),
.Y(n_3262)
);

BUFx3_ASAP7_75t_L g3263 ( 
.A(n_2758),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2731),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_SL g3265 ( 
.A(n_2729),
.B(n_1279),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2652),
.B(n_1501),
.Y(n_3266)
);

BUFx6f_ASAP7_75t_L g3267 ( 
.A(n_2740),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2581),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_2415),
.B(n_1281),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2731),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_2415),
.B(n_1282),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_2614),
.B(n_1502),
.Y(n_3272)
);

AND2x6_ASAP7_75t_L g3273 ( 
.A(n_2635),
.B(n_1272),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_2734),
.B(n_1286),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_2731),
.Y(n_3275)
);

NOR2x1p5_ASAP7_75t_L g3276 ( 
.A(n_2405),
.B(n_1298),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_2581),
.Y(n_3277)
);

NOR2xp33_ASAP7_75t_L g3278 ( 
.A(n_2415),
.B(n_1314),
.Y(n_3278)
);

BUFx6f_ASAP7_75t_L g3279 ( 
.A(n_2740),
.Y(n_3279)
);

INVx3_ASAP7_75t_L g3280 ( 
.A(n_2581),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2417),
.Y(n_3281)
);

AND2x2_ASAP7_75t_SL g3282 ( 
.A(n_2635),
.B(n_1135),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2417),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_2415),
.B(n_1339),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_2758),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_2415),
.B(n_1357),
.Y(n_3286)
);

INVx4_ASAP7_75t_L g3287 ( 
.A(n_2758),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2417),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2417),
.Y(n_3289)
);

BUFx6f_ASAP7_75t_L g3290 ( 
.A(n_2740),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2417),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2417),
.Y(n_3292)
);

INVx5_ASAP7_75t_L g3293 ( 
.A(n_2758),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2417),
.Y(n_3294)
);

BUFx3_ASAP7_75t_L g3295 ( 
.A(n_2758),
.Y(n_3295)
);

BUFx4f_ASAP7_75t_L g3296 ( 
.A(n_2571),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_2734),
.B(n_1371),
.Y(n_3297)
);

BUFx2_ASAP7_75t_L g3298 ( 
.A(n_2729),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2417),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2734),
.B(n_1377),
.Y(n_3300)
);

AND2x4_ASAP7_75t_L g3301 ( 
.A(n_2614),
.B(n_1507),
.Y(n_3301)
);

BUFx6f_ASAP7_75t_L g3302 ( 
.A(n_2740),
.Y(n_3302)
);

INVx4_ASAP7_75t_SL g3303 ( 
.A(n_2405),
.Y(n_3303)
);

INVx4_ASAP7_75t_L g3304 ( 
.A(n_2758),
.Y(n_3304)
);

INVxp67_ASAP7_75t_L g3305 ( 
.A(n_2725),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_2415),
.B(n_1381),
.Y(n_3306)
);

AOI22xp33_ASAP7_75t_L g3307 ( 
.A1(n_2715),
.A2(n_1382),
.B1(n_1443),
.B2(n_1414),
.Y(n_3307)
);

BUFx6f_ASAP7_75t_L g3308 ( 
.A(n_2740),
.Y(n_3308)
);

BUFx2_ASAP7_75t_L g3309 ( 
.A(n_2729),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2652),
.B(n_1511),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_2415),
.B(n_1482),
.Y(n_3311)
);

INVx4_ASAP7_75t_L g3312 ( 
.A(n_2758),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2652),
.B(n_1514),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2731),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2731),
.Y(n_3315)
);

AO22x2_ASAP7_75t_L g3316 ( 
.A1(n_2731),
.A2(n_1515),
.B1(n_1518),
.B2(n_1516),
.Y(n_3316)
);

AND2x6_ASAP7_75t_L g3317 ( 
.A(n_2635),
.B(n_1272),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_2415),
.B(n_1499),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_2734),
.B(n_1526),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_2731),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_2731),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2731),
.Y(n_3322)
);

INVx4_ASAP7_75t_L g3323 ( 
.A(n_2758),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_L g3324 ( 
.A(n_2415),
.B(n_1528),
.Y(n_3324)
);

INVx3_ASAP7_75t_L g3325 ( 
.A(n_2581),
.Y(n_3325)
);

OR2x2_ASAP7_75t_L g3326 ( 
.A(n_2724),
.B(n_1531),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2417),
.Y(n_3327)
);

INVx4_ASAP7_75t_L g3328 ( 
.A(n_2758),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2731),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2731),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_2731),
.Y(n_3331)
);

OR2x2_ASAP7_75t_L g3332 ( 
.A(n_2724),
.B(n_1566),
.Y(n_3332)
);

NOR2xp33_ASAP7_75t_L g3333 ( 
.A(n_2415),
.B(n_1591),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2417),
.Y(n_3334)
);

INVx1_ASAP7_75t_SL g3335 ( 
.A(n_2729),
.Y(n_3335)
);

NOR2xp33_ASAP7_75t_L g3336 ( 
.A(n_2415),
.B(n_1609),
.Y(n_3336)
);

INVx8_ASAP7_75t_L g3337 ( 
.A(n_2758),
.Y(n_3337)
);

NAND3xp33_ASAP7_75t_L g3338 ( 
.A(n_2654),
.B(n_1426),
.C(n_1272),
.Y(n_3338)
);

NAND2x1p5_ASAP7_75t_L g3339 ( 
.A(n_2375),
.B(n_1426),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_SL g3340 ( 
.A(n_2405),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2731),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2417),
.Y(n_3342)
);

AOI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_2729),
.A2(n_1631),
.B1(n_1661),
.B2(n_1614),
.Y(n_3343)
);

BUFx6f_ASAP7_75t_L g3344 ( 
.A(n_2740),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2417),
.Y(n_3345)
);

INVx4_ASAP7_75t_L g3346 ( 
.A(n_2758),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2417),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2415),
.B(n_1668),
.Y(n_3348)
);

INVx3_ASAP7_75t_L g3349 ( 
.A(n_2581),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_2731),
.Y(n_3350)
);

INVxp33_ASAP7_75t_L g3351 ( 
.A(n_2381),
.Y(n_3351)
);

OAI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_2731),
.A2(n_1221),
.B1(n_1233),
.B2(n_1188),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2417),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2417),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_2729),
.B(n_1653),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_2734),
.B(n_1520),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2417),
.Y(n_3357)
);

AND2x2_ASAP7_75t_SL g3358 ( 
.A(n_2635),
.B(n_1188),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_2417),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2417),
.Y(n_3360)
);

BUFx2_ASAP7_75t_L g3361 ( 
.A(n_2729),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2652),
.B(n_1523),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_2729),
.B(n_1653),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2417),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_2715),
.A2(n_1605),
.B1(n_1653),
.B2(n_1553),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_2614),
.B(n_1530),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_2652),
.B(n_1533),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_2734),
.B(n_1534),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2415),
.B(n_1538),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_2729),
.B(n_1653),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2731),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2731),
.Y(n_3372)
);

CKINVDCx5p33_ASAP7_75t_R g3373 ( 
.A(n_2589),
.Y(n_3373)
);

INVx4_ASAP7_75t_L g3374 ( 
.A(n_2758),
.Y(n_3374)
);

INVx2_ASAP7_75t_SL g3375 ( 
.A(n_2758),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_2415),
.B(n_1539),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_2415),
.B(n_1543),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2652),
.B(n_1547),
.Y(n_3378)
);

HB1xp67_ASAP7_75t_L g3379 ( 
.A(n_2729),
.Y(n_3379)
);

INVx3_ASAP7_75t_L g3380 ( 
.A(n_2581),
.Y(n_3380)
);

BUFx3_ASAP7_75t_L g3381 ( 
.A(n_2758),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2417),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2652),
.B(n_1550),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_2729),
.B(n_1553),
.Y(n_3384)
);

NOR2x1p5_ASAP7_75t_L g3385 ( 
.A(n_2405),
.B(n_1669),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_2729),
.B(n_1553),
.Y(n_3386)
);

INVxp67_ASAP7_75t_SL g3387 ( 
.A(n_2725),
.Y(n_3387)
);

INVx1_ASAP7_75t_SL g3388 ( 
.A(n_2729),
.Y(n_3388)
);

NAND3x1_ASAP7_75t_L g3389 ( 
.A(n_2710),
.B(n_1559),
.C(n_1558),
.Y(n_3389)
);

AND2x6_ASAP7_75t_L g3390 ( 
.A(n_2635),
.B(n_1426),
.Y(n_3390)
);

BUFx2_ASAP7_75t_L g3391 ( 
.A(n_2729),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_2652),
.B(n_1563),
.Y(n_3392)
);

INVx4_ASAP7_75t_SL g3393 ( 
.A(n_2405),
.Y(n_3393)
);

BUFx6f_ASAP7_75t_L g3394 ( 
.A(n_2740),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_2415),
.B(n_1567),
.Y(n_3395)
);

INVx4_ASAP7_75t_L g3396 ( 
.A(n_2758),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_L g3397 ( 
.A1(n_2715),
.A2(n_1605),
.B1(n_1653),
.B2(n_1553),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_2734),
.B(n_1568),
.Y(n_3398)
);

AND2x4_ASAP7_75t_L g3399 ( 
.A(n_2614),
.B(n_1575),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2417),
.Y(n_3400)
);

INVx4_ASAP7_75t_L g3401 ( 
.A(n_2758),
.Y(n_3401)
);

INVx2_ASAP7_75t_SL g3402 ( 
.A(n_2758),
.Y(n_3402)
);

INVx3_ASAP7_75t_L g3403 ( 
.A(n_2581),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2731),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_2731),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_2417),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2417),
.Y(n_3407)
);

AND2x6_ASAP7_75t_L g3408 ( 
.A(n_2635),
.B(n_1426),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_2758),
.Y(n_3409)
);

INVx4_ASAP7_75t_L g3410 ( 
.A(n_2758),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_2731),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2417),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_2734),
.B(n_1577),
.Y(n_3413)
);

BUFx3_ASAP7_75t_L g3414 ( 
.A(n_2758),
.Y(n_3414)
);

CKINVDCx5p33_ASAP7_75t_R g3415 ( 
.A(n_2589),
.Y(n_3415)
);

OR2x2_ASAP7_75t_L g3416 ( 
.A(n_2724),
.B(n_1580),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_SL g3417 ( 
.A(n_2729),
.B(n_1221),
.Y(n_3417)
);

AOI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_2729),
.A2(n_1581),
.B1(n_1588),
.B2(n_1586),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2652),
.B(n_1589),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2417),
.Y(n_3420)
);

INVx4_ASAP7_75t_L g3421 ( 
.A(n_2758),
.Y(n_3421)
);

INVx2_ASAP7_75t_SL g3422 ( 
.A(n_2758),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_2740),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3417),
.B(n_1479),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2816),
.B(n_1596),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_SL g3426 ( 
.A(n_3201),
.B(n_1479),
.Y(n_3426)
);

INVx2_ASAP7_75t_SL g3427 ( 
.A(n_3337),
.Y(n_3427)
);

NAND2x1_ASAP7_75t_L g3428 ( 
.A(n_3093),
.B(n_1479),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3201),
.B(n_1479),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_2884),
.B(n_1599),
.Y(n_3430)
);

AOI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_3061),
.A2(n_1600),
.B1(n_1613),
.B2(n_1606),
.Y(n_3431)
);

CKINVDCx20_ASAP7_75t_R g3432 ( 
.A(n_3256),
.Y(n_3432)
);

INVx1_ASAP7_75t_SL g3433 ( 
.A(n_2796),
.Y(n_3433)
);

BUFx6f_ASAP7_75t_L g3434 ( 
.A(n_2781),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_SL g3435 ( 
.A(n_3199),
.B(n_1506),
.Y(n_3435)
);

OAI22xp33_ASAP7_75t_L g3436 ( 
.A1(n_3031),
.A2(n_1618),
.B1(n_1619),
.B2(n_1615),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2994),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_2765),
.Y(n_3438)
);

NAND2xp33_ASAP7_75t_L g3439 ( 
.A(n_3093),
.B(n_1553),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_3199),
.B(n_1506),
.Y(n_3440)
);

A2O1A1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_3100),
.A2(n_1234),
.B(n_1246),
.C(n_1233),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_L g3442 ( 
.A(n_2781),
.Y(n_3442)
);

AND2x6_ASAP7_75t_L g3443 ( 
.A(n_3202),
.B(n_1506),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_3204),
.B(n_1506),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3166),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_2768),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_2772),
.Y(n_3447)
);

NAND3xp33_ASAP7_75t_L g3448 ( 
.A(n_3338),
.B(n_1681),
.C(n_1579),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_2773),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_2846),
.B(n_1621),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3169),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_2999),
.B(n_1626),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_L g3453 ( 
.A(n_3228),
.B(n_1627),
.Y(n_3453)
);

NOR3xp33_ASAP7_75t_L g3454 ( 
.A(n_2948),
.B(n_1635),
.C(n_1633),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3172),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3175),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3413),
.B(n_1638),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_2777),
.Y(n_3458)
);

INVxp67_ASAP7_75t_L g3459 ( 
.A(n_2852),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3176),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3356),
.B(n_1645),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2783),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3368),
.B(n_1646),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2790),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3177),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_3204),
.B(n_1681),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_3351),
.B(n_1647),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3398),
.B(n_1657),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_2912),
.B(n_1681),
.Y(n_3469)
);

NAND2x1_ASAP7_75t_L g3470 ( 
.A(n_3093),
.B(n_1681),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_2912),
.B(n_1605),
.Y(n_3471)
);

BUFx8_ASAP7_75t_L g3472 ( 
.A(n_3340),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_2908),
.B(n_1658),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3193),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_2942),
.B(n_1688),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_2885),
.B(n_1605),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3183),
.B(n_1431),
.Y(n_3477)
);

INVx4_ASAP7_75t_L g3478 ( 
.A(n_3337),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_2909),
.Y(n_3479)
);

OAI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3203),
.A2(n_1246),
.B1(n_1248),
.B2(n_1234),
.Y(n_3480)
);

INVx3_ASAP7_75t_L g3481 ( 
.A(n_3093),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3186),
.B(n_3187),
.Y(n_3482)
);

BUFx5_ASAP7_75t_L g3483 ( 
.A(n_2901),
.Y(n_3483)
);

INVxp67_ASAP7_75t_L g3484 ( 
.A(n_2779),
.Y(n_3484)
);

NAND2xp33_ASAP7_75t_SL g3485 ( 
.A(n_2880),
.B(n_1248),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3205),
.Y(n_3486)
);

NAND2xp33_ASAP7_75t_L g3487 ( 
.A(n_2901),
.B(n_1605),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_2897),
.A2(n_1297),
.B1(n_1299),
.B2(n_1276),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3069),
.B(n_1276),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3206),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3208),
.B(n_1297),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3129),
.B(n_1299),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3282),
.B(n_1653),
.Y(n_3493)
);

AND2x4_ASAP7_75t_L g3494 ( 
.A(n_3212),
.B(n_1301),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2791),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3358),
.B(n_1653),
.Y(n_3496)
);

INVxp67_ASAP7_75t_L g3497 ( 
.A(n_3298),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3051),
.B(n_1301),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_2829),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_2821),
.B(n_1605),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2807),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2888),
.B(n_1311),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_2830),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_2848),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_2821),
.B(n_1605),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2821),
.B(n_1311),
.Y(n_3506)
);

OAI221xp5_ASAP7_75t_L g3507 ( 
.A1(n_2774),
.A2(n_1435),
.B1(n_1542),
.B2(n_1412),
.C(n_1370),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_2951),
.B(n_1370),
.Y(n_3508)
);

AOI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_2960),
.A2(n_1435),
.B1(n_1542),
.B2(n_1412),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2812),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_SL g3511 ( 
.A(n_3195),
.B(n_1608),
.Y(n_3511)
);

INVx2_ASAP7_75t_SL g3512 ( 
.A(n_2831),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_2962),
.B(n_1608),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_2972),
.B(n_1610),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_2824),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_2976),
.B(n_1610),
.Y(n_3516)
);

O2A1O1Ixp33_ASAP7_75t_L g3517 ( 
.A1(n_2995),
.A2(n_1677),
.B(n_4),
.C(n_2),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_2832),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_SL g3519 ( 
.A(n_3309),
.B(n_1677),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_2987),
.B(n_2833),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_2836),
.B(n_2),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_2865),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_2839),
.B(n_3),
.Y(n_3523)
);

INVx3_ASAP7_75t_L g3524 ( 
.A(n_3261),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3188),
.B(n_3),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_2857),
.B(n_4),
.Y(n_3526)
);

NOR2xp33_ASAP7_75t_L g3527 ( 
.A(n_3218),
.B(n_5),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_2859),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3219),
.Y(n_3529)
);

INVx2_ASAP7_75t_SL g3530 ( 
.A(n_2831),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_2770),
.B(n_2841),
.Y(n_3531)
);

OR2x2_ASAP7_75t_L g3532 ( 
.A(n_2820),
.B(n_5),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3220),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3238),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3225),
.B(n_6),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3230),
.B(n_6),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3232),
.B(n_6),
.Y(n_3537)
);

NOR2xp33_ASAP7_75t_L g3538 ( 
.A(n_3379),
.B(n_7),
.Y(n_3538)
);

INVxp67_ASAP7_75t_SL g3539 ( 
.A(n_2875),
.Y(n_3539)
);

INVx1_ASAP7_75t_SL g3540 ( 
.A(n_3000),
.Y(n_3540)
);

BUFx5_ASAP7_75t_L g3541 ( 
.A(n_2901),
.Y(n_3541)
);

BUFx6f_ASAP7_75t_L g3542 ( 
.A(n_2781),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_2872),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_2902),
.B(n_7),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3239),
.B(n_8),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3246),
.B(n_8),
.Y(n_3546)
);

INVxp33_ASAP7_75t_L g3547 ( 
.A(n_3361),
.Y(n_3547)
);

AND2x4_ASAP7_75t_L g3548 ( 
.A(n_3248),
.B(n_8),
.Y(n_3548)
);

INVxp67_ASAP7_75t_L g3549 ( 
.A(n_3391),
.Y(n_3549)
);

AND2x4_ASAP7_75t_L g3550 ( 
.A(n_3248),
.B(n_9),
.Y(n_3550)
);

OR2x6_ASAP7_75t_L g3551 ( 
.A(n_2798),
.B(n_10),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3257),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_2886),
.Y(n_3553)
);

AND2x2_ASAP7_75t_L g3554 ( 
.A(n_2892),
.B(n_10),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3020),
.B(n_937),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3281),
.B(n_10),
.Y(n_3556)
);

AOI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_2952),
.A2(n_2797),
.B1(n_2992),
.B2(n_3016),
.Y(n_3557)
);

BUFx6f_ASAP7_75t_SL g3558 ( 
.A(n_2873),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3283),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_2889),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_2914),
.B(n_11),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_2953),
.B(n_11),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3288),
.B(n_12),
.Y(n_3563)
);

OAI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3110),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3289),
.Y(n_3565)
);

INVx4_ASAP7_75t_L g3566 ( 
.A(n_3248),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_2894),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_2854),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_SL g3569 ( 
.A(n_2780),
.B(n_3224),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_2900),
.Y(n_3570)
);

OAI22xp5_ASAP7_75t_L g3571 ( 
.A1(n_2992),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_3571)
);

OR2x6_ASAP7_75t_L g3572 ( 
.A(n_2798),
.B(n_16),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3291),
.B(n_17),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3292),
.B(n_17),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3294),
.B(n_3299),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3234),
.B(n_938),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3327),
.B(n_18),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3334),
.B(n_18),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3342),
.B(n_3345),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_2907),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3347),
.B(n_18),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3353),
.B(n_3354),
.Y(n_3582)
);

AOI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_3052),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3357),
.B(n_20),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3359),
.B(n_20),
.Y(n_3585)
);

INVxp67_ASAP7_75t_L g3586 ( 
.A(n_2827),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_SL g3587 ( 
.A(n_3335),
.B(n_938),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_2954),
.B(n_21),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_3388),
.B(n_21),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3360),
.B(n_22),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3364),
.B(n_22),
.Y(n_3591)
);

INVxp67_ASAP7_75t_L g3592 ( 
.A(n_3164),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_3293),
.B(n_939),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3382),
.B(n_23),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3400),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2913),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_3293),
.B(n_940),
.Y(n_3597)
);

NOR2xp33_ASAP7_75t_L g3598 ( 
.A(n_3196),
.B(n_23),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3406),
.B(n_23),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3407),
.B(n_24),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_3293),
.B(n_940),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_2766),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_2767),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3412),
.B(n_24),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3101),
.B(n_24),
.Y(n_3605)
);

INVx2_ASAP7_75t_SL g3606 ( 
.A(n_3296),
.Y(n_3606)
);

AOI221xp5_ASAP7_75t_L g3607 ( 
.A1(n_3369),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.C(n_28),
.Y(n_3607)
);

INVx8_ASAP7_75t_L g3608 ( 
.A(n_3340),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3420),
.Y(n_3609)
);

INVx1_ASAP7_75t_SL g3610 ( 
.A(n_2850),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_2771),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_2849),
.B(n_942),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_2996),
.B(n_25),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3022),
.B(n_26),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3042),
.B(n_26),
.Y(n_3615)
);

NAND2xp33_ASAP7_75t_L g3616 ( 
.A(n_2901),
.B(n_27),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_2849),
.B(n_2855),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_2860),
.Y(n_3618)
);

AOI22xp5_ASAP7_75t_L g3619 ( 
.A1(n_2776),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_3619)
);

INVx2_ASAP7_75t_SL g3620 ( 
.A(n_3296),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_2819),
.B(n_2823),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_2834),
.B(n_28),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_2969),
.B(n_29),
.Y(n_3623)
);

AOI22xp5_ASAP7_75t_L g3624 ( 
.A1(n_2764),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_3624)
);

NAND2xp33_ASAP7_75t_L g3625 ( 
.A(n_2883),
.B(n_30),
.Y(n_3625)
);

OAI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3031),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3416),
.B(n_31),
.Y(n_3627)
);

CKINVDCx5p33_ASAP7_75t_R g3628 ( 
.A(n_2775),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_2778),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_2782),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_2975),
.B(n_32),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_2979),
.B(n_32),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_2903),
.B(n_33),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3222),
.B(n_33),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_2985),
.B(n_33),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3223),
.B(n_34),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3227),
.B(n_34),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_2880),
.B(n_35),
.Y(n_3638)
);

NAND3xp33_ASAP7_75t_L g3639 ( 
.A(n_3365),
.B(n_35),
.C(n_36),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_2849),
.B(n_942),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_2861),
.Y(n_3641)
);

INVx3_ASAP7_75t_L g3642 ( 
.A(n_3261),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3190),
.A2(n_3213),
.B(n_3217),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3237),
.B(n_36),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_2993),
.B(n_36),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_SL g3646 ( 
.A(n_2855),
.B(n_2858),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_2871),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_2786),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_2784),
.Y(n_3649)
);

A2O1A1Ixp33_ASAP7_75t_L g3650 ( 
.A1(n_3120),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_2789),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3258),
.B(n_37),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3266),
.B(n_37),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_2799),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_2877),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3310),
.B(n_38),
.Y(n_3656)
);

INVx4_ASAP7_75t_L g3657 ( 
.A(n_2785),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_SL g3658 ( 
.A(n_2855),
.B(n_943),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_2878),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_2881),
.Y(n_3660)
);

AND2x6_ASAP7_75t_SL g3661 ( 
.A(n_3083),
.B(n_38),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_2804),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_2806),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_2966),
.B(n_39),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_2858),
.B(n_944),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_2898),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_L g3667 ( 
.A(n_3226),
.B(n_40),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3313),
.B(n_40),
.Y(n_3668)
);

INVxp67_ASAP7_75t_L g3669 ( 
.A(n_3041),
.Y(n_3669)
);

NAND2x1_ASAP7_75t_L g3670 ( 
.A(n_2814),
.B(n_40),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3362),
.B(n_3367),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_2809),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_2813),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2905),
.Y(n_3674)
);

INVx2_ASAP7_75t_SL g3675 ( 
.A(n_3263),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3378),
.B(n_41),
.Y(n_3676)
);

NAND3xp33_ASAP7_75t_SL g3677 ( 
.A(n_3015),
.B(n_3415),
.C(n_3373),
.Y(n_3677)
);

BUFx8_ASAP7_75t_L g3678 ( 
.A(n_3295),
.Y(n_3678)
);

OAI22xp5_ASAP7_75t_L g3679 ( 
.A1(n_3316),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_3679)
);

AOI22xp5_ASAP7_75t_L g3680 ( 
.A1(n_2870),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_2911),
.Y(n_3681)
);

AND2x4_ASAP7_75t_L g3682 ( 
.A(n_2785),
.B(n_42),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_2915),
.Y(n_3683)
);

HB1xp67_ASAP7_75t_L g3684 ( 
.A(n_3249),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_SL g3685 ( 
.A1(n_3111),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_2858),
.B(n_944),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_SL g3687 ( 
.A(n_2922),
.B(n_945),
.Y(n_3687)
);

INVx4_ASAP7_75t_L g3688 ( 
.A(n_3233),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_2922),
.B(n_947),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_2922),
.B(n_947),
.Y(n_3690)
);

BUFx8_ASAP7_75t_L g3691 ( 
.A(n_3381),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3383),
.B(n_3392),
.Y(n_3692)
);

INVx2_ASAP7_75t_SL g3693 ( 
.A(n_3414),
.Y(n_3693)
);

INVx4_ASAP7_75t_L g3694 ( 
.A(n_3233),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3419),
.B(n_44),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3305),
.B(n_45),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3221),
.Y(n_3697)
);

CKINVDCx5p33_ASAP7_75t_R g3698 ( 
.A(n_2828),
.Y(n_3698)
);

NOR2xp67_ASAP7_75t_L g3699 ( 
.A(n_2869),
.B(n_46),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3102),
.B(n_45),
.Y(n_3700)
);

BUFx8_ASAP7_75t_L g3701 ( 
.A(n_2769),
.Y(n_3701)
);

INVxp67_ASAP7_75t_L g3702 ( 
.A(n_3107),
.Y(n_3702)
);

INVxp67_ASAP7_75t_L g3703 ( 
.A(n_3387),
.Y(n_3703)
);

BUFx3_ASAP7_75t_L g3704 ( 
.A(n_2910),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3123),
.B(n_46),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3012),
.B(n_46),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_SL g3707 ( 
.A(n_2956),
.B(n_948),
.Y(n_3707)
);

NAND3xp33_ASAP7_75t_L g3708 ( 
.A(n_3397),
.B(n_2844),
.C(n_3229),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3235),
.Y(n_3709)
);

AND2x6_ASAP7_75t_SL g3710 ( 
.A(n_2854),
.B(n_2808),
.Y(n_3710)
);

AND3x1_ASAP7_75t_L g3711 ( 
.A(n_3079),
.B(n_47),
.C(n_48),
.Y(n_3711)
);

INVx5_ASAP7_75t_L g3712 ( 
.A(n_2814),
.Y(n_3712)
);

BUFx3_ASAP7_75t_L g3713 ( 
.A(n_2941),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3240),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3012),
.B(n_47),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3140),
.B(n_48),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3245),
.Y(n_3717)
);

AOI22xp33_ASAP7_75t_L g3718 ( 
.A1(n_2931),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3105),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3112),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3251),
.Y(n_3721)
);

NOR2xp67_ASAP7_75t_L g3722 ( 
.A(n_2869),
.B(n_50),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_L g3723 ( 
.A(n_2784),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3113),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_L g3725 ( 
.A(n_2932),
.B(n_49),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_2933),
.B(n_49),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3137),
.B(n_50),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_L g3728 ( 
.A(n_2800),
.B(n_51),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_2918),
.B(n_2920),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3117),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_2924),
.B(n_52),
.Y(n_3731)
);

AOI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3253),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3118),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3316),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_2925),
.B(n_53),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_2926),
.B(n_54),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_2928),
.B(n_55),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_2956),
.B(n_948),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3264),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3148),
.A2(n_55),
.B(n_56),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3108),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_2935),
.B(n_2943),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_2944),
.B(n_56),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_2949),
.B(n_57),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3046),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3262),
.B(n_3274),
.Y(n_3746)
);

BUFx6f_ASAP7_75t_L g3747 ( 
.A(n_2784),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_2923),
.B(n_57),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3270),
.Y(n_3749)
);

NOR2xp67_ASAP7_75t_L g3750 ( 
.A(n_2792),
.B(n_59),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3297),
.B(n_3300),
.Y(n_3751)
);

INVxp33_ASAP7_75t_L g3752 ( 
.A(n_2940),
.Y(n_3752)
);

INVx2_ASAP7_75t_SL g3753 ( 
.A(n_2838),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3319),
.B(n_58),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3275),
.Y(n_3755)
);

OAI221xp5_ASAP7_75t_L g3756 ( 
.A1(n_3418),
.A2(n_61),
.B1(n_58),
.B2(n_60),
.C(n_63),
.Y(n_3756)
);

INVxp67_ASAP7_75t_L g3757 ( 
.A(n_3250),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3046),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_2956),
.B(n_949),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3147),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_2998),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3073),
.B(n_58),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_2862),
.B(n_60),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_2811),
.B(n_61),
.Y(n_3764)
);

A2O1A1Ixp33_ASAP7_75t_L g3765 ( 
.A1(n_3121),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3184),
.B(n_63),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_SL g3767 ( 
.A(n_3010),
.B(n_951),
.Y(n_3767)
);

INVxp67_ASAP7_75t_L g3768 ( 
.A(n_3250),
.Y(n_3768)
);

BUFx6f_ASAP7_75t_L g3769 ( 
.A(n_3231),
.Y(n_3769)
);

NOR2xp67_ASAP7_75t_L g3770 ( 
.A(n_2792),
.B(n_65),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3072),
.B(n_64),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_SL g3772 ( 
.A(n_3010),
.B(n_2906),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3320),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_2937),
.B(n_2938),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_2787),
.B(n_64),
.Y(n_3775)
);

INVxp67_ASAP7_75t_L g3776 ( 
.A(n_3272),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3019),
.Y(n_3777)
);

OAI22xp5_ASAP7_75t_L g3778 ( 
.A1(n_3242),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3326),
.B(n_66),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_2906),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_3170),
.B(n_951),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3332),
.B(n_67),
.Y(n_3782)
);

NAND3xp33_ASAP7_75t_L g3783 ( 
.A(n_3124),
.B(n_68),
.C(n_69),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3321),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3272),
.B(n_68),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_SL g3786 ( 
.A(n_3089),
.B(n_952),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3023),
.Y(n_3787)
);

INVx5_ASAP7_75t_L g3788 ( 
.A(n_2814),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_3158),
.A2(n_69),
.B(n_70),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3152),
.B(n_69),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3331),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_2788),
.B(n_70),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3153),
.B(n_3021),
.Y(n_3793)
);

INVx2_ASAP7_75t_SL g3794 ( 
.A(n_2838),
.Y(n_3794)
);

BUFx6f_ASAP7_75t_SL g3795 ( 
.A(n_2873),
.Y(n_3795)
);

OAI221xp5_ASAP7_75t_L g3796 ( 
.A1(n_2930),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.C(n_74),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3045),
.B(n_71),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3341),
.Y(n_3798)
);

NOR3xp33_ASAP7_75t_L g3799 ( 
.A(n_3136),
.B(n_71),
.C(n_72),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3003),
.B(n_3018),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3350),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3068),
.B(n_73),
.Y(n_3802)
);

INVxp67_ASAP7_75t_L g3803 ( 
.A(n_3301),
.Y(n_3803)
);

AND2x4_ASAP7_75t_L g3804 ( 
.A(n_3236),
.B(n_74),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3024),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3075),
.B(n_3077),
.Y(n_3806)
);

NOR2xp33_ASAP7_75t_L g3807 ( 
.A(n_3154),
.B(n_74),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3371),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3028),
.B(n_75),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3025),
.Y(n_3810)
);

OAI22xp5_ASAP7_75t_L g3811 ( 
.A1(n_3372),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3811)
);

AND2x2_ASAP7_75t_SL g3812 ( 
.A(n_3089),
.B(n_76),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3027),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3037),
.B(n_76),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_SL g3815 ( 
.A(n_3111),
.B(n_952),
.Y(n_3815)
);

AOI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3114),
.A2(n_3017),
.B1(n_3063),
.B2(n_3252),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3035),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3404),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_SL g3819 ( 
.A(n_2879),
.B(n_953),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3301),
.B(n_77),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3053),
.B(n_78),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3001),
.B(n_78),
.Y(n_3822)
);

OAI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3405),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_2879),
.B(n_953),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_2893),
.B(n_954),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3047),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_SL g3827 ( 
.A(n_2893),
.B(n_954),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3048),
.Y(n_3828)
);

OAI22xp33_ASAP7_75t_L g3829 ( 
.A1(n_3136),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_2921),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3830)
);

INVx4_ASAP7_75t_L g3831 ( 
.A(n_3236),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3050),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_SL g3833 ( 
.A(n_3149),
.B(n_955),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3119),
.B(n_82),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_SL g3835 ( 
.A(n_3287),
.B(n_82),
.Y(n_3835)
);

NOR2x1p5_ASAP7_75t_L g3836 ( 
.A(n_3149),
.B(n_83),
.Y(n_3836)
);

AOI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3255),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3376),
.B(n_83),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3054),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3411),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3056),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_2921),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3377),
.B(n_85),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3395),
.B(n_86),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3165),
.B(n_86),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_SL g3846 ( 
.A(n_3044),
.B(n_955),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_2936),
.B(n_87),
.Y(n_3847)
);

NAND2x1p5_ASAP7_75t_L g3848 ( 
.A(n_3287),
.B(n_87),
.Y(n_3848)
);

INVx4_ASAP7_75t_L g3849 ( 
.A(n_3304),
.Y(n_3849)
);

OAI22xp33_ASAP7_75t_L g3850 ( 
.A1(n_2808),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_2959),
.B(n_88),
.Y(n_3851)
);

NOR2xp33_ASAP7_75t_L g3852 ( 
.A(n_2818),
.B(n_88),
.Y(n_3852)
);

INVxp67_ASAP7_75t_L g3853 ( 
.A(n_3366),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3059),
.Y(n_3854)
);

AOI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3366),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_2964),
.B(n_89),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_2974),
.B(n_91),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_2983),
.B(n_92),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_2986),
.B(n_92),
.Y(n_3859)
);

BUFx2_ASAP7_75t_L g3860 ( 
.A(n_3304),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_SL g3861 ( 
.A(n_3044),
.B(n_956),
.Y(n_3861)
);

AOI22xp5_ASAP7_75t_L g3862 ( 
.A1(n_3259),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3862)
);

INVx4_ASAP7_75t_L g3863 ( 
.A(n_3312),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3060),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_2990),
.B(n_2847),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3082),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3084),
.Y(n_3867)
);

INVx2_ASAP7_75t_SL g3868 ( 
.A(n_3312),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_3399),
.B(n_956),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3399),
.B(n_957),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3151),
.B(n_93),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_2895),
.B(n_93),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_2896),
.B(n_94),
.Y(n_3873)
);

AOI22xp5_ASAP7_75t_L g3874 ( 
.A1(n_3260),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_3874)
);

INVxp67_ASAP7_75t_L g3875 ( 
.A(n_3269),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_2916),
.B(n_95),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3122),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_2843),
.B(n_958),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_2927),
.B(n_96),
.Y(n_3879)
);

INVx2_ASAP7_75t_SL g3880 ( 
.A(n_3323),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_SL g3881 ( 
.A(n_2843),
.B(n_2845),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_2845),
.B(n_2864),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_SL g3883 ( 
.A(n_2864),
.B(n_958),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_SL g3884 ( 
.A(n_2887),
.B(n_959),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3138),
.B(n_960),
.Y(n_3885)
);

AO22x2_ASAP7_75t_L g3886 ( 
.A1(n_2793),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_2970),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_2927),
.B(n_98),
.Y(n_3888)
);

AOI22xp33_ASAP7_75t_L g3889 ( 
.A1(n_2837),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3092),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_2984),
.B(n_960),
.Y(n_3891)
);

CKINVDCx5p33_ASAP7_75t_R g3892 ( 
.A(n_2822),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_2984),
.B(n_961),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3133),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_2978),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3103),
.B(n_100),
.Y(n_3896)
);

INVx2_ASAP7_75t_SL g3897 ( 
.A(n_3323),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_2957),
.B(n_101),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3144),
.B(n_102),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_2981),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3013),
.B(n_102),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_2837),
.B(n_961),
.Y(n_3902)
);

BUFx5_ASAP7_75t_L g3903 ( 
.A(n_2883),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_2868),
.B(n_3125),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3125),
.B(n_962),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_2957),
.B(n_103),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2968),
.B(n_103),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3125),
.B(n_962),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3070),
.B(n_963),
.Y(n_3909)
);

AOI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3271),
.A2(n_3284),
.B1(n_3286),
.B2(n_3278),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3306),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_3911)
);

AO22x2_ASAP7_75t_L g3912 ( 
.A1(n_2793),
.A2(n_2795),
.B1(n_2802),
.B2(n_2794),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_2989),
.Y(n_3913)
);

AND2x2_ASAP7_75t_SL g3914 ( 
.A(n_3328),
.B(n_104),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_SL g3915 ( 
.A(n_3070),
.B(n_963),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_2968),
.B(n_105),
.Y(n_3916)
);

BUFx2_ASAP7_75t_SL g3917 ( 
.A(n_3328),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_SL g3918 ( 
.A(n_3070),
.B(n_964),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_2997),
.Y(n_3919)
);

NOR2xp33_ASAP7_75t_L g3920 ( 
.A(n_3209),
.B(n_105),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3055),
.B(n_106),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_2794),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3150),
.Y(n_3923)
);

OAI22xp5_ASAP7_75t_L g3924 ( 
.A1(n_2795),
.A2(n_109),
.B1(n_106),
.B2(n_108),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3005),
.B(n_106),
.Y(n_3925)
);

NOR3xp33_ASAP7_75t_L g3926 ( 
.A(n_3157),
.B(n_108),
.C(n_109),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3161),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3127),
.Y(n_3928)
);

NAND2xp33_ASAP7_75t_L g3929 ( 
.A(n_2883),
.B(n_108),
.Y(n_3929)
);

NAND3xp33_ASAP7_75t_L g3930 ( 
.A(n_3352),
.B(n_2917),
.C(n_3115),
.Y(n_3930)
);

INVx2_ASAP7_75t_SL g3931 ( 
.A(n_3346),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3005),
.B(n_110),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3008),
.B(n_110),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3131),
.Y(n_3934)
);

NAND2x1p5_ASAP7_75t_L g3935 ( 
.A(n_3346),
.B(n_110),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3142),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_SL g3937 ( 
.A(n_3074),
.B(n_964),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3145),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3008),
.B(n_111),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_2802),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_2826),
.B(n_111),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_2817),
.B(n_112),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_SL g3943 ( 
.A(n_3074),
.B(n_965),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3162),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_2947),
.B(n_112),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3374),
.Y(n_3946)
);

INVx2_ASAP7_75t_L g3947 ( 
.A(n_3314),
.Y(n_3947)
);

OAI221xp5_ASAP7_75t_L g3948 ( 
.A1(n_2863),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.C(n_116),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_2810),
.B(n_114),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3074),
.B(n_966),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3314),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3315),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_L g3953 ( 
.A(n_3091),
.B(n_114),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3004),
.Y(n_3954)
);

AOI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3311),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3006),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3318),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3065),
.B(n_117),
.Y(n_3958)
);

BUFx3_ASAP7_75t_L g3959 ( 
.A(n_3374),
.Y(n_3959)
);

INVxp67_ASAP7_75t_SL g3960 ( 
.A(n_3094),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3096),
.B(n_118),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3071),
.B(n_3171),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3094),
.B(n_966),
.Y(n_3963)
);

NOR2xp67_ASAP7_75t_L g3964 ( 
.A(n_3315),
.B(n_119),
.Y(n_3964)
);

INVx2_ASAP7_75t_SL g3965 ( 
.A(n_3396),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3066),
.Y(n_3966)
);

INVx6_ASAP7_75t_L g3967 ( 
.A(n_3396),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3174),
.B(n_118),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3094),
.B(n_967),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3180),
.B(n_118),
.Y(n_3970)
);

HB1xp67_ASAP7_75t_L g3971 ( 
.A(n_3401),
.Y(n_3971)
);

AND2x4_ASAP7_75t_L g3972 ( 
.A(n_3401),
.B(n_119),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3385),
.B(n_119),
.Y(n_3973)
);

INVxp67_ASAP7_75t_L g3974 ( 
.A(n_3324),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3076),
.Y(n_3975)
);

NAND2xp33_ASAP7_75t_L g3976 ( 
.A(n_2883),
.B(n_120),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3095),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3097),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_L g3979 ( 
.A(n_3215),
.B(n_120),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3182),
.B(n_3057),
.Y(n_3980)
);

INVxp67_ASAP7_75t_L g3981 ( 
.A(n_3333),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3192),
.B(n_120),
.Y(n_3982)
);

AND2x2_ASAP7_75t_L g3983 ( 
.A(n_3211),
.B(n_3343),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_2882),
.B(n_968),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3322),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3126),
.Y(n_3986)
);

AOI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3336),
.A2(n_124),
.B1(n_121),
.B2(n_122),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3322),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3038),
.A2(n_124),
.B1(n_121),
.B2(n_122),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3057),
.B(n_121),
.Y(n_3990)
);

AND2x2_ASAP7_75t_SL g3991 ( 
.A(n_3410),
.B(n_124),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_2891),
.B(n_969),
.Y(n_3992)
);

OR2x2_ASAP7_75t_L g3993 ( 
.A(n_3410),
.B(n_125),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3329),
.Y(n_3994)
);

NOR2xp67_ASAP7_75t_L g3995 ( 
.A(n_3329),
.B(n_3330),
.Y(n_3995)
);

INVx8_ASAP7_75t_L g3996 ( 
.A(n_2856),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3173),
.B(n_125),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_3478),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3486),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3531),
.B(n_3389),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3490),
.Y(n_4001)
);

INVx1_ASAP7_75t_SL g4002 ( 
.A(n_3917),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3912),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3912),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3671),
.B(n_3330),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3437),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3746),
.B(n_3914),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3712),
.B(n_3198),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_3712),
.B(n_3198),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3692),
.B(n_3430),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3991),
.B(n_3078),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_SL g4012 ( 
.A(n_3712),
.B(n_3198),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3450),
.B(n_3475),
.Y(n_4013)
);

OAI22xp5_ASAP7_75t_L g4014 ( 
.A1(n_3621),
.A2(n_3086),
.B1(n_3216),
.B2(n_2929),
.Y(n_4014)
);

INVx4_ASAP7_75t_L g4015 ( 
.A(n_3478),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3438),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3446),
.Y(n_4017)
);

NAND3xp33_ASAP7_75t_SL g4018 ( 
.A(n_3835),
.B(n_3067),
.C(n_3049),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3454),
.A2(n_3207),
.B1(n_3078),
.B2(n_3159),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3447),
.Y(n_4020)
);

BUFx6f_ASAP7_75t_L g4021 ( 
.A(n_3959),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3734),
.B(n_3085),
.Y(n_4022)
);

AND2x6_ASAP7_75t_L g4023 ( 
.A(n_3481),
.B(n_3231),
.Y(n_4023)
);

BUFx6f_ASAP7_75t_L g4024 ( 
.A(n_3704),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3445),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3449),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3458),
.Y(n_4027)
);

INVx2_ASAP7_75t_SL g4028 ( 
.A(n_3678),
.Y(n_4028)
);

BUFx3_ASAP7_75t_L g4029 ( 
.A(n_3678),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_SL g4030 ( 
.A1(n_3812),
.A2(n_2955),
.B1(n_2967),
.B2(n_2890),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3751),
.B(n_3087),
.Y(n_4031)
);

OR2x2_ASAP7_75t_L g4032 ( 
.A(n_3433),
.B(n_2866),
.Y(n_4032)
);

BUFx6f_ASAP7_75t_L g4033 ( 
.A(n_3713),
.Y(n_4033)
);

A2O1A1Ixp33_ASAP7_75t_L g4034 ( 
.A1(n_3616),
.A2(n_3143),
.B(n_3207),
.C(n_3178),
.Y(n_4034)
);

BUFx4f_ASAP7_75t_L g4035 ( 
.A(n_3608),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3664),
.B(n_3452),
.Y(n_4036)
);

AOI22xp5_ASAP7_75t_L g4037 ( 
.A1(n_3436),
.A2(n_3348),
.B1(n_3276),
.B2(n_3191),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3462),
.B(n_3464),
.Y(n_4038)
);

NAND2x1p5_ASAP7_75t_L g4039 ( 
.A(n_3657),
.B(n_3688),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3495),
.B(n_3501),
.Y(n_4040)
);

NOR2xp33_ASAP7_75t_L g4041 ( 
.A(n_3547),
.B(n_3265),
.Y(n_4041)
);

OAI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_3557),
.A2(n_2934),
.B1(n_2950),
.B2(n_2945),
.Y(n_4042)
);

AND2x4_ASAP7_75t_L g4043 ( 
.A(n_3481),
.B(n_2803),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_3451),
.Y(n_4044)
);

INVx2_ASAP7_75t_SL g4045 ( 
.A(n_3691),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3510),
.B(n_3087),
.Y(n_4046)
);

BUFx3_ASAP7_75t_L g4047 ( 
.A(n_3691),
.Y(n_4047)
);

AND2x2_ASAP7_75t_SL g4048 ( 
.A(n_3625),
.B(n_3421),
.Y(n_4048)
);

AOI21xp5_ASAP7_75t_L g4049 ( 
.A1(n_3439),
.A2(n_2835),
.B(n_3231),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_SL g4050 ( 
.A(n_3788),
.B(n_3699),
.Y(n_4050)
);

OAI22xp5_ASAP7_75t_SL g4051 ( 
.A1(n_3551),
.A2(n_2939),
.B1(n_2876),
.B2(n_3030),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3515),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_SL g4053 ( 
.A1(n_3443),
.A2(n_2955),
.B1(n_2967),
.B2(n_2890),
.Y(n_4053)
);

NAND2x1p5_ASAP7_75t_L g4054 ( 
.A(n_3657),
.B(n_3421),
.Y(n_4054)
);

INVx1_ASAP7_75t_SL g4055 ( 
.A(n_3860),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3518),
.B(n_3194),
.Y(n_4056)
);

AOI22xp33_ASAP7_75t_L g4057 ( 
.A1(n_3926),
.A2(n_3159),
.B1(n_3106),
.B2(n_3135),
.Y(n_4057)
);

INVx2_ASAP7_75t_SL g4058 ( 
.A(n_3967),
.Y(n_4058)
);

AOI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3790),
.A2(n_3159),
.B1(n_3106),
.B2(n_3135),
.Y(n_4059)
);

BUFx5_ASAP7_75t_L g4060 ( 
.A(n_3443),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3528),
.B(n_3062),
.Y(n_4061)
);

AOI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3431),
.A2(n_3200),
.B1(n_3214),
.B2(n_3210),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_3788),
.B(n_2803),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_R g4064 ( 
.A(n_3432),
.B(n_3034),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3455),
.Y(n_4065)
);

AOI22xp5_ASAP7_75t_SL g4066 ( 
.A1(n_3592),
.A2(n_2840),
.B1(n_2801),
.B2(n_3159),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3529),
.Y(n_4067)
);

INVx4_ASAP7_75t_L g4068 ( 
.A(n_3688),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3701),
.Y(n_4069)
);

BUFx3_ASAP7_75t_L g4070 ( 
.A(n_3701),
.Y(n_4070)
);

BUFx12f_ASAP7_75t_L g4071 ( 
.A(n_3472),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_3785),
.B(n_3007),
.Y(n_4072)
);

AND2x4_ASAP7_75t_L g4073 ( 
.A(n_3788),
.B(n_2805),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3533),
.B(n_3307),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3552),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3559),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3565),
.Y(n_4077)
);

BUFx6f_ASAP7_75t_L g4078 ( 
.A(n_3534),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3595),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3456),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3460),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3609),
.B(n_2904),
.Y(n_4082)
);

NOR2xp33_ASAP7_75t_L g4083 ( 
.A(n_3875),
.B(n_2842),
.Y(n_4083)
);

BUFx3_ASAP7_75t_L g4084 ( 
.A(n_3967),
.Y(n_4084)
);

CKINVDCx5p33_ASAP7_75t_R g4085 ( 
.A(n_3472),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3760),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3465),
.Y(n_4087)
);

INVx1_ASAP7_75t_SL g4088 ( 
.A(n_3971),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3520),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3474),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3575),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3579),
.Y(n_4092)
);

AO22x2_ASAP7_75t_L g4093 ( 
.A1(n_3571),
.A2(n_3090),
.B1(n_3155),
.B2(n_2961),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_3499),
.Y(n_4094)
);

AND2x4_ASAP7_75t_L g4095 ( 
.A(n_3995),
.B(n_2805),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3582),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3618),
.Y(n_4097)
);

BUFx6f_ASAP7_75t_L g4098 ( 
.A(n_3434),
.Y(n_4098)
);

AOI22xp5_ASAP7_75t_L g4099 ( 
.A1(n_3816),
.A2(n_3064),
.B1(n_3139),
.B2(n_3128),
.Y(n_4099)
);

AOI22xp33_ASAP7_75t_SL g4100 ( 
.A1(n_3443),
.A2(n_2955),
.B1(n_2967),
.B2(n_2890),
.Y(n_4100)
);

CKINVDCx5p33_ASAP7_75t_R g4101 ( 
.A(n_3628),
.Y(n_4101)
);

BUFx6f_ASAP7_75t_L g4102 ( 
.A(n_3434),
.Y(n_4102)
);

BUFx2_ASAP7_75t_L g4103 ( 
.A(n_3539),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3482),
.B(n_2973),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3641),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_L g4106 ( 
.A(n_3974),
.B(n_3029),
.Y(n_4106)
);

INVx2_ASAP7_75t_SL g4107 ( 
.A(n_3694),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3647),
.Y(n_4108)
);

INVxp67_ASAP7_75t_L g4109 ( 
.A(n_3684),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3981),
.B(n_3007),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3699),
.B(n_3241),
.Y(n_4111)
);

BUFx6f_ASAP7_75t_L g4112 ( 
.A(n_3434),
.Y(n_4112)
);

AND2x4_ASAP7_75t_L g4113 ( 
.A(n_3995),
.B(n_2851),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3807),
.A2(n_3128),
.B1(n_3135),
.B2(n_3106),
.Y(n_4114)
);

INVx4_ASAP7_75t_L g4115 ( 
.A(n_3694),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3503),
.Y(n_4116)
);

INVx2_ASAP7_75t_SL g4117 ( 
.A(n_3831),
.Y(n_4117)
);

AND2x4_ASAP7_75t_L g4118 ( 
.A(n_3741),
.B(n_2851),
.Y(n_4118)
);

BUFx3_ASAP7_75t_L g4119 ( 
.A(n_3427),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3504),
.Y(n_4120)
);

INVx3_ASAP7_75t_L g4121 ( 
.A(n_3831),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_3820),
.B(n_3058),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3655),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3659),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_SL g4125 ( 
.A(n_3722),
.B(n_3241),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3522),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_SL g4127 ( 
.A(n_3722),
.B(n_3241),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3543),
.Y(n_4128)
);

INVx2_ASAP7_75t_SL g4129 ( 
.A(n_3849),
.Y(n_4129)
);

CKINVDCx5p33_ASAP7_75t_R g4130 ( 
.A(n_3608),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_3544),
.B(n_3622),
.Y(n_4131)
);

INVx2_ASAP7_75t_SL g4132 ( 
.A(n_3849),
.Y(n_4132)
);

BUFx3_ASAP7_75t_L g4133 ( 
.A(n_3512),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_3558),
.Y(n_4134)
);

INVx4_ASAP7_75t_L g4135 ( 
.A(n_3863),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_3553),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_SL g4137 ( 
.A(n_3903),
.B(n_3244),
.Y(n_4137)
);

INVx3_ASAP7_75t_L g4138 ( 
.A(n_3863),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_SL g4139 ( 
.A(n_3903),
.B(n_3244),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3457),
.B(n_3461),
.Y(n_4140)
);

BUFx4f_ASAP7_75t_SL g4141 ( 
.A(n_3530),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3463),
.B(n_3146),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_SL g4143 ( 
.A(n_3903),
.B(n_3244),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3468),
.B(n_3080),
.Y(n_4144)
);

INVxp67_ASAP7_75t_L g4145 ( 
.A(n_3993),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3560),
.Y(n_4146)
);

INVxp67_ASAP7_75t_SL g4147 ( 
.A(n_3929),
.Y(n_4147)
);

INVx3_ASAP7_75t_L g4148 ( 
.A(n_3566),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_SL g4149 ( 
.A(n_3903),
.B(n_3247),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_3425),
.B(n_3088),
.Y(n_4150)
);

CKINVDCx5p33_ASAP7_75t_R g4151 ( 
.A(n_3558),
.Y(n_4151)
);

AND2x4_ASAP7_75t_L g4152 ( 
.A(n_3745),
.B(n_3243),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3660),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_3567),
.Y(n_4154)
);

AND2x4_ASAP7_75t_L g4155 ( 
.A(n_3758),
.B(n_3243),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_SL g4156 ( 
.A(n_3903),
.B(n_3750),
.Y(n_4156)
);

INVx4_ASAP7_75t_L g4157 ( 
.A(n_3996),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3774),
.B(n_3098),
.Y(n_4158)
);

NOR2x2_ASAP7_75t_L g4159 ( 
.A(n_3551),
.B(n_3303),
.Y(n_4159)
);

BUFx3_ASAP7_75t_L g4160 ( 
.A(n_3996),
.Y(n_4160)
);

NOR2xp33_ASAP7_75t_R g4161 ( 
.A(n_3710),
.B(n_2946),
.Y(n_4161)
);

OR2x6_ASAP7_75t_L g4162 ( 
.A(n_3572),
.B(n_2801),
.Y(n_4162)
);

INVx2_ASAP7_75t_SL g4163 ( 
.A(n_3868),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_3623),
.A2(n_3128),
.B1(n_3135),
.B2(n_3106),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3635),
.A2(n_3128),
.B1(n_3185),
.B2(n_3116),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3473),
.B(n_3099),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3666),
.Y(n_4167)
);

AND2x4_ASAP7_75t_L g4168 ( 
.A(n_3988),
.B(n_3268),
.Y(n_4168)
);

AND2x4_ASAP7_75t_L g4169 ( 
.A(n_3994),
.B(n_3268),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3865),
.B(n_3141),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3674),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3570),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3800),
.B(n_3160),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_3580),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_SL g4175 ( 
.A(n_3750),
.B(n_3247),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_SL g4176 ( 
.A(n_3770),
.B(n_3247),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3681),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_3683),
.B(n_3277),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3923),
.Y(n_4179)
);

NAND3xp33_ASAP7_75t_SL g4180 ( 
.A(n_3848),
.B(n_3179),
.C(n_2840),
.Y(n_4180)
);

BUFx4f_ASAP7_75t_SL g4181 ( 
.A(n_3606),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_3566),
.Y(n_4182)
);

BUFx2_ASAP7_75t_L g4183 ( 
.A(n_3443),
.Y(n_4183)
);

BUFx6f_ASAP7_75t_L g4184 ( 
.A(n_3442),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3596),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_SL g4186 ( 
.A(n_3770),
.B(n_3267),
.Y(n_4186)
);

AND2x4_ASAP7_75t_L g4187 ( 
.A(n_3927),
.B(n_3277),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3719),
.Y(n_4188)
);

AND2x4_ASAP7_75t_L g4189 ( 
.A(n_3720),
.B(n_3280),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_3645),
.A2(n_3185),
.B1(n_3116),
.B2(n_3109),
.Y(n_4190)
);

NAND2xp33_ASAP7_75t_L g4191 ( 
.A(n_3483),
.B(n_3185),
.Y(n_4191)
);

INVx3_ASAP7_75t_L g4192 ( 
.A(n_3880),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3806),
.B(n_3160),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_3561),
.B(n_3178),
.Y(n_4194)
);

NOR2xp33_ASAP7_75t_L g4195 ( 
.A(n_3910),
.B(n_2899),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3554),
.B(n_3109),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3588),
.B(n_3104),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_3602),
.Y(n_4198)
);

INVx4_ASAP7_75t_L g4199 ( 
.A(n_3795),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3724),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_3730),
.Y(n_4201)
);

AOI21xp5_ASAP7_75t_L g4202 ( 
.A1(n_3487),
.A2(n_3279),
.B(n_3267),
.Y(n_4202)
);

INVx2_ASAP7_75t_SL g4203 ( 
.A(n_3897),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3733),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3761),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_3603),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_SL g4207 ( 
.A(n_3964),
.B(n_3267),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3562),
.B(n_3130),
.Y(n_4208)
);

INVx2_ASAP7_75t_SL g4209 ( 
.A(n_3931),
.Y(n_4209)
);

INVx5_ASAP7_75t_L g4210 ( 
.A(n_3572),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_SL g4211 ( 
.A(n_3964),
.B(n_3279),
.Y(n_4211)
);

BUFx2_ASAP7_75t_L g4212 ( 
.A(n_3483),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_3611),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3453),
.B(n_3375),
.Y(n_4214)
);

OR2x6_ASAP7_75t_L g4215 ( 
.A(n_3669),
.B(n_3285),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3777),
.Y(n_4216)
);

INVxp67_ASAP7_75t_L g4217 ( 
.A(n_3667),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3787),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_3702),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3805),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3810),
.Y(n_4221)
);

INVxp67_ASAP7_75t_L g4222 ( 
.A(n_3696),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3813),
.Y(n_4223)
);

INVx1_ASAP7_75t_SL g4224 ( 
.A(n_3610),
.Y(n_4224)
);

CKINVDCx5p33_ASAP7_75t_R g4225 ( 
.A(n_3795),
.Y(n_4225)
);

OAI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_3930),
.A2(n_3339),
.B1(n_3254),
.B2(n_3325),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3817),
.Y(n_4227)
);

OAI22xp5_ASAP7_75t_SL g4228 ( 
.A1(n_3711),
.A2(n_3409),
.B1(n_3422),
.B2(n_3402),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3467),
.B(n_3189),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_3483),
.B(n_3279),
.Y(n_4230)
);

NOR2xp33_ASAP7_75t_L g4231 ( 
.A(n_3484),
.B(n_3132),
.Y(n_4231)
);

AND2x6_ASAP7_75t_L g4232 ( 
.A(n_3638),
.B(n_3290),
.Y(n_4232)
);

CKINVDCx5p33_ASAP7_75t_R g4233 ( 
.A(n_3892),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_3793),
.B(n_3983),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3779),
.B(n_3156),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_3782),
.B(n_3156),
.Y(n_4236)
);

BUFx3_ASAP7_75t_L g4237 ( 
.A(n_3946),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3826),
.Y(n_4238)
);

AND3x2_ASAP7_75t_SL g4239 ( 
.A(n_3836),
.B(n_3393),
.C(n_3303),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_3828),
.Y(n_4240)
);

AOI22xp33_ASAP7_75t_L g4241 ( 
.A1(n_3852),
.A2(n_3185),
.B1(n_3363),
.B2(n_3355),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_3953),
.A2(n_3384),
.B1(n_3386),
.B2(n_3370),
.Y(n_4242)
);

NOR2xp33_ASAP7_75t_L g4243 ( 
.A(n_3497),
.B(n_3549),
.Y(n_4243)
);

AND2x4_ASAP7_75t_L g4244 ( 
.A(n_3832),
.B(n_3280),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3839),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3629),
.Y(n_4246)
);

OAI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_3492),
.A2(n_3167),
.B(n_2853),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_R g4248 ( 
.A(n_3677),
.B(n_2946),
.Y(n_4248)
);

BUFx6f_ASAP7_75t_L g4249 ( 
.A(n_3965),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_SL g4250 ( 
.A(n_3483),
.B(n_3290),
.Y(n_4250)
);

AND2x4_ASAP7_75t_L g4251 ( 
.A(n_3841),
.B(n_3854),
.Y(n_4251)
);

A2O1A1Ixp33_ASAP7_75t_SL g4252 ( 
.A1(n_3725),
.A2(n_3349),
.B(n_3380),
.C(n_3325),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_3630),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3899),
.B(n_3189),
.Y(n_4254)
);

OAI21xp33_ASAP7_75t_SL g4255 ( 
.A1(n_3435),
.A2(n_2955),
.B(n_2890),
.Y(n_4255)
);

INVx5_ASAP7_75t_L g4256 ( 
.A(n_3548),
.Y(n_4256)
);

INVx2_ASAP7_75t_SL g4257 ( 
.A(n_3675),
.Y(n_4257)
);

NAND2xp33_ASAP7_75t_SL g4258 ( 
.A(n_3428),
.B(n_3290),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3864),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_3961),
.A2(n_2967),
.B1(n_3181),
.B2(n_2825),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_3627),
.B(n_3189),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3757),
.B(n_2988),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_3698),
.Y(n_4263)
);

OAI22xp5_ASAP7_75t_L g4264 ( 
.A1(n_3680),
.A2(n_3380),
.B1(n_3403),
.B2(n_3349),
.Y(n_4264)
);

NOR2x2_ASAP7_75t_L g4265 ( 
.A(n_3661),
.B(n_3393),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_3866),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_3648),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3768),
.B(n_2988),
.Y(n_4268)
);

INVx2_ASAP7_75t_SL g4269 ( 
.A(n_3693),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3776),
.B(n_2991),
.Y(n_4270)
);

AND2x4_ASAP7_75t_L g4271 ( 
.A(n_3867),
.B(n_3403),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3803),
.B(n_2991),
.Y(n_4272)
);

NAND2x1p5_ASAP7_75t_L g4273 ( 
.A(n_3620),
.B(n_2958),
.Y(n_4273)
);

OAI21xp33_ASAP7_75t_SL g4274 ( 
.A1(n_3440),
.A2(n_3466),
.B(n_3444),
.Y(n_4274)
);

INVxp67_ASAP7_75t_SL g4275 ( 
.A(n_3976),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_3853),
.B(n_3009),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3890),
.Y(n_4277)
);

INVx3_ASAP7_75t_L g4278 ( 
.A(n_3524),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3488),
.B(n_3634),
.Y(n_4279)
);

AOI22xp5_ASAP7_75t_L g4280 ( 
.A1(n_3762),
.A2(n_3168),
.B1(n_3134),
.B2(n_2815),
.Y(n_4280)
);

INVx1_ASAP7_75t_SL g4281 ( 
.A(n_3540),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3928),
.Y(n_4282)
);

AO22x1_ASAP7_75t_L g4283 ( 
.A1(n_3548),
.A2(n_2815),
.B1(n_3273),
.B2(n_2814),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3934),
.Y(n_4284)
);

INVx3_ASAP7_75t_L g4285 ( 
.A(n_3524),
.Y(n_4285)
);

NAND2x1p5_ASAP7_75t_L g4286 ( 
.A(n_3550),
.B(n_2958),
.Y(n_4286)
);

AND2x6_ASAP7_75t_L g4287 ( 
.A(n_3638),
.B(n_3302),
.Y(n_4287)
);

INVx4_ASAP7_75t_L g4288 ( 
.A(n_3550),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3636),
.B(n_3009),
.Y(n_4289)
);

INVx1_ASAP7_75t_SL g4290 ( 
.A(n_3569),
.Y(n_4290)
);

NOR2xp67_ASAP7_75t_L g4291 ( 
.A(n_3479),
.B(n_3155),
.Y(n_4291)
);

INVx2_ASAP7_75t_SL g4292 ( 
.A(n_3682),
.Y(n_4292)
);

OR2x2_ASAP7_75t_SL g4293 ( 
.A(n_3532),
.B(n_3181),
.Y(n_4293)
);

OR2x6_ASAP7_75t_L g4294 ( 
.A(n_3935),
.B(n_3134),
.Y(n_4294)
);

BUFx3_ASAP7_75t_L g4295 ( 
.A(n_3753),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_3483),
.B(n_3302),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_3936),
.Y(n_4297)
);

AND2x2_ASAP7_75t_SL g4298 ( 
.A(n_3682),
.B(n_3302),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3938),
.Y(n_4299)
);

NAND2xp33_ASAP7_75t_L g4300 ( 
.A(n_3541),
.B(n_2815),
.Y(n_4300)
);

OR2x2_ASAP7_75t_L g4301 ( 
.A(n_3459),
.B(n_3032),
.Y(n_4301)
);

NOR2x2_ASAP7_75t_L g4302 ( 
.A(n_3922),
.B(n_2963),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_3637),
.B(n_3032),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_3644),
.B(n_3033),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_3652),
.B(n_3033),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3944),
.Y(n_4306)
);

BUFx6f_ASAP7_75t_L g4307 ( 
.A(n_3442),
.Y(n_4307)
);

AOI22xp5_ASAP7_75t_L g4308 ( 
.A1(n_3920),
.A2(n_3273),
.B1(n_3317),
.B2(n_2815),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_3894),
.Y(n_4309)
);

O2A1O1Ixp33_ASAP7_75t_L g4310 ( 
.A1(n_3771),
.A2(n_3838),
.B(n_3844),
.C(n_3843),
.Y(n_4310)
);

INVx2_ASAP7_75t_SL g4311 ( 
.A(n_3804),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3895),
.Y(n_4312)
);

OAI221xp5_ASAP7_75t_L g4313 ( 
.A1(n_3799),
.A2(n_3040),
.B1(n_3081),
.B2(n_3043),
.C(n_2919),
.Y(n_4313)
);

NAND2xp33_ASAP7_75t_L g4314 ( 
.A(n_3541),
.B(n_3273),
.Y(n_4314)
);

CKINVDCx20_ASAP7_75t_R g4315 ( 
.A(n_3794),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_3653),
.B(n_3040),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_3541),
.B(n_3308),
.Y(n_4317)
);

AOI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_3896),
.A2(n_3317),
.B1(n_3390),
.B2(n_3273),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_3651),
.Y(n_4319)
);

INVx5_ASAP7_75t_L g4320 ( 
.A(n_3442),
.Y(n_4320)
);

AND2x4_ASAP7_75t_L g4321 ( 
.A(n_3470),
.B(n_2977),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_SL g4322 ( 
.A(n_3541),
.B(n_3308),
.Y(n_4322)
);

O2A1O1Ixp33_ASAP7_75t_L g4323 ( 
.A1(n_3555),
.A2(n_3043),
.B(n_3081),
.C(n_2965),
.Y(n_4323)
);

AND2x4_ASAP7_75t_L g4324 ( 
.A(n_3940),
.B(n_2977),
.Y(n_4324)
);

AOI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_3728),
.A2(n_3390),
.B1(n_3408),
.B2(n_3317),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_3541),
.B(n_3308),
.Y(n_4326)
);

INVxp67_ASAP7_75t_L g4327 ( 
.A(n_3489),
.Y(n_4327)
);

INVx2_ASAP7_75t_SL g4328 ( 
.A(n_3804),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_3485),
.B(n_3511),
.Y(n_4329)
);

NOR2xp67_ASAP7_75t_L g4330 ( 
.A(n_3703),
.B(n_2982),
.Y(n_4330)
);

INVx3_ASAP7_75t_L g4331 ( 
.A(n_3642),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3656),
.B(n_3668),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_SL g4333 ( 
.A(n_3626),
.B(n_3344),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_3676),
.B(n_3181),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_3900),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_3695),
.B(n_3498),
.Y(n_4336)
);

INVx2_ASAP7_75t_SL g4337 ( 
.A(n_3972),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_3654),
.Y(n_4338)
);

HB1xp67_ASAP7_75t_L g4339 ( 
.A(n_3586),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_3901),
.B(n_3197),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_3729),
.B(n_3197),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_3919),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3742),
.B(n_3197),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_SL g4344 ( 
.A(n_3642),
.B(n_3344),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_3982),
.B(n_126),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_3613),
.B(n_2982),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_3886),
.Y(n_4347)
);

INVx3_ASAP7_75t_L g4348 ( 
.A(n_3972),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_3886),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3614),
.B(n_3036),
.Y(n_4350)
);

INVx5_ASAP7_75t_L g4351 ( 
.A(n_3542),
.Y(n_4351)
);

BUFx2_ASAP7_75t_L g4352 ( 
.A(n_3960),
.Y(n_4352)
);

AND2x4_ASAP7_75t_L g4353 ( 
.A(n_3947),
.B(n_3390),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_3615),
.B(n_3036),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_SL g4355 ( 
.A(n_3426),
.B(n_3344),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_3662),
.Y(n_4356)
);

AOI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_3979),
.A2(n_3390),
.B1(n_3408),
.B2(n_3317),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3954),
.Y(n_4358)
);

AOI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_3945),
.A2(n_3036),
.B1(n_3011),
.B2(n_2874),
.Y(n_4359)
);

OR2x6_ASAP7_75t_L g4360 ( 
.A(n_3772),
.B(n_3394),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_3663),
.Y(n_4361)
);

BUFx2_ASAP7_75t_L g4362 ( 
.A(n_3542),
.Y(n_4362)
);

NOR2xp33_ASAP7_75t_L g4363 ( 
.A(n_3881),
.B(n_3882),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_3887),
.Y(n_4364)
);

INVx5_ASAP7_75t_L g4365 ( 
.A(n_3542),
.Y(n_4365)
);

BUFx6f_ASAP7_75t_L g4366 ( 
.A(n_3649),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_SL g4367 ( 
.A(n_3429),
.B(n_3394),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_3766),
.B(n_3036),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3956),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_3966),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_3975),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_3705),
.B(n_3011),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_3672),
.Y(n_4373)
);

NOR2xp33_ASAP7_75t_L g4374 ( 
.A(n_3752),
.B(n_127),
.Y(n_4374)
);

AND2x4_ASAP7_75t_L g4375 ( 
.A(n_3951),
.B(n_3408),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_3977),
.Y(n_4376)
);

INVx3_ASAP7_75t_L g4377 ( 
.A(n_3913),
.Y(n_4377)
);

INVxp67_ASAP7_75t_L g4378 ( 
.A(n_3527),
.Y(n_4378)
);

AO22x1_ASAP7_75t_L g4379 ( 
.A1(n_3973),
.A2(n_3408),
.B1(n_2874),
.B2(n_2867),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_3525),
.A2(n_2874),
.B1(n_2867),
.B2(n_3011),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3978),
.Y(n_4381)
);

AND2x4_ASAP7_75t_L g4382 ( 
.A(n_3952),
.B(n_3394),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_3673),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_3986),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_3809),
.B(n_3011),
.Y(n_4385)
);

NAND2x1_ASAP7_75t_L g4386 ( 
.A(n_3649),
.B(n_3423),
.Y(n_4386)
);

OAI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_3583),
.A2(n_3423),
.B1(n_3163),
.B2(n_3014),
.Y(n_4387)
);

INVx3_ASAP7_75t_L g4388 ( 
.A(n_3985),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_3697),
.Y(n_4389)
);

INVx1_ASAP7_75t_SL g4390 ( 
.A(n_3904),
.Y(n_4390)
);

NOR2xp33_ASAP7_75t_L g4391 ( 
.A(n_3519),
.B(n_127),
.Y(n_4391)
);

BUFx6f_ASAP7_75t_L g4392 ( 
.A(n_3649),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_L g4393 ( 
.A(n_3726),
.B(n_3958),
.Y(n_4393)
);

AND2x2_ASAP7_75t_SL g4394 ( 
.A(n_3568),
.B(n_3423),
.Y(n_4394)
);

BUFx3_ASAP7_75t_L g4395 ( 
.A(n_3709),
.Y(n_4395)
);

AND2x4_ASAP7_75t_L g4396 ( 
.A(n_3714),
.B(n_2867),
.Y(n_4396)
);

INVx1_ASAP7_75t_SL g4397 ( 
.A(n_3494),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_SL g4398 ( 
.A(n_3885),
.B(n_3163),
.Y(n_4398)
);

INVx4_ASAP7_75t_L g4399 ( 
.A(n_3723),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_3717),
.Y(n_4400)
);

BUFx6f_ASAP7_75t_L g4401 ( 
.A(n_3723),
.Y(n_4401)
);

HB1xp67_ASAP7_75t_L g4402 ( 
.A(n_3721),
.Y(n_4402)
);

BUFx8_ASAP7_75t_SL g4403 ( 
.A(n_3494),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3521),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_SL g4405 ( 
.A(n_3564),
.B(n_3163),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_3523),
.Y(n_4406)
);

INVx5_ASAP7_75t_L g4407 ( 
.A(n_3723),
.Y(n_4407)
);

BUFx4f_ASAP7_75t_L g4408 ( 
.A(n_3739),
.Y(n_4408)
);

BUFx6f_ASAP7_75t_L g4409 ( 
.A(n_3747),
.Y(n_4409)
);

BUFx12f_ASAP7_75t_L g4410 ( 
.A(n_3747),
.Y(n_4410)
);

AND2x4_ASAP7_75t_L g4411 ( 
.A(n_3749),
.B(n_2867),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_3814),
.B(n_128),
.Y(n_4412)
);

INVx3_ASAP7_75t_L g4413 ( 
.A(n_3755),
.Y(n_4413)
);

BUFx6f_ASAP7_75t_L g4414 ( 
.A(n_3747),
.Y(n_4414)
);

CKINVDCx5p33_ASAP7_75t_R g4415 ( 
.A(n_3605),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_3821),
.B(n_128),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_3526),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_3631),
.B(n_128),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_3633),
.B(n_129),
.Y(n_4419)
);

NOR2xp33_ASAP7_75t_L g4420 ( 
.A(n_3754),
.B(n_129),
.Y(n_4420)
);

NOR2x1p5_ASAP7_75t_L g4421 ( 
.A(n_3670),
.B(n_2874),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_3535),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_3536),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_3537),
.Y(n_4424)
);

INVx2_ASAP7_75t_SL g4425 ( 
.A(n_3469),
.Y(n_4425)
);

INVx4_ASAP7_75t_L g4426 ( 
.A(n_3769),
.Y(n_4426)
);

AND2x6_ASAP7_75t_SL g4427 ( 
.A(n_3589),
.B(n_3538),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_SL g4428 ( 
.A(n_3850),
.B(n_3002),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_3773),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_3685),
.B(n_130),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_3727),
.B(n_130),
.Y(n_4431)
);

AOI22xp33_ASAP7_75t_L g4432 ( 
.A1(n_3756),
.A2(n_2971),
.B1(n_2980),
.B2(n_3039),
.Y(n_4432)
);

O2A1O1Ixp5_ASAP7_75t_L g4433 ( 
.A1(n_3424),
.A2(n_2980),
.B(n_2971),
.C(n_3039),
.Y(n_4433)
);

BUFx3_ASAP7_75t_L g4434 ( 
.A(n_3784),
.Y(n_4434)
);

AND2x4_ASAP7_75t_L g4435 ( 
.A(n_3791),
.B(n_2971),
.Y(n_4435)
);

AOI22xp5_ASAP7_75t_L g4436 ( 
.A1(n_3598),
.A2(n_2980),
.B1(n_2971),
.B2(n_3039),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_3545),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_3798),
.Y(n_4438)
);

BUFx3_ASAP7_75t_L g4439 ( 
.A(n_3801),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3546),
.Y(n_4440)
);

CKINVDCx5p33_ASAP7_75t_R g4441 ( 
.A(n_3679),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_3716),
.B(n_3632),
.Y(n_4442)
);

NOR2xp67_ASAP7_75t_L g4443 ( 
.A(n_3997),
.B(n_131),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_3808),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3556),
.Y(n_4445)
);

BUFx3_ASAP7_75t_L g4446 ( 
.A(n_3818),
.Y(n_4446)
);

INVx2_ASAP7_75t_SL g4447 ( 
.A(n_3840),
.Y(n_4447)
);

INVx2_ASAP7_75t_SL g4448 ( 
.A(n_3781),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_3775),
.B(n_131),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_3792),
.B(n_131),
.Y(n_4450)
);

BUFx3_ASAP7_75t_L g4451 ( 
.A(n_3769),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_3731),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_3735),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_3563),
.Y(n_4454)
);

NOR2xp33_ASAP7_75t_L g4455 ( 
.A(n_3871),
.B(n_132),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_3925),
.B(n_132),
.Y(n_4456)
);

INVx5_ASAP7_75t_L g4457 ( 
.A(n_3769),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_3573),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_SL g4459 ( 
.A(n_3517),
.B(n_3002),
.Y(n_4459)
);

AND2x2_ASAP7_75t_SL g4460 ( 
.A(n_3780),
.B(n_3014),
.Y(n_4460)
);

OAI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_3718),
.A2(n_3026),
.B1(n_3014),
.B2(n_3002),
.Y(n_4461)
);

INVx1_ASAP7_75t_SL g4462 ( 
.A(n_3932),
.Y(n_4462)
);

AOI22xp33_ASAP7_75t_L g4463 ( 
.A1(n_3796),
.A2(n_2980),
.B1(n_3039),
.B2(n_3026),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_3933),
.B(n_133),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_3748),
.B(n_133),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_3574),
.Y(n_4466)
);

OR2x2_ASAP7_75t_L g4467 ( 
.A(n_3939),
.B(n_133),
.Y(n_4467)
);

HB1xp67_ASAP7_75t_L g4468 ( 
.A(n_3879),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_3736),
.Y(n_4469)
);

AOI22xp5_ASAP7_75t_L g4470 ( 
.A1(n_3869),
.A2(n_3026),
.B1(n_136),
.B2(n_134),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_3783),
.B(n_134),
.Y(n_4471)
);

AND3x2_ASAP7_75t_SL g4472 ( 
.A(n_3829),
.B(n_134),
.C(n_135),
.Y(n_4472)
);

INVx5_ASAP7_75t_L g4473 ( 
.A(n_3617),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_3577),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3700),
.B(n_137),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_3578),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_3846),
.B(n_137),
.Y(n_4477)
);

BUFx2_ASAP7_75t_L g4478 ( 
.A(n_3962),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_3581),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_3584),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_3847),
.B(n_137),
.Y(n_4481)
);

NOR2xp33_ASAP7_75t_L g4482 ( 
.A(n_3921),
.B(n_138),
.Y(n_4482)
);

OR2x6_ASAP7_75t_L g4483 ( 
.A(n_3819),
.B(n_138),
.Y(n_4483)
);

INVx2_ASAP7_75t_L g4484 ( 
.A(n_3737),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_3851),
.B(n_138),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_3743),
.Y(n_4486)
);

INVxp67_ASAP7_75t_L g4487 ( 
.A(n_3888),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_3585),
.Y(n_4488)
);

BUFx3_ASAP7_75t_L g4489 ( 
.A(n_3898),
.Y(n_4489)
);

NOR2xp33_ASAP7_75t_L g4490 ( 
.A(n_3942),
.B(n_3949),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_3856),
.B(n_3857),
.Y(n_4491)
);

BUFx6f_ASAP7_75t_L g4492 ( 
.A(n_3646),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_3902),
.B(n_139),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_SL g4494 ( 
.A(n_3861),
.B(n_139),
.Y(n_4494)
);

AOI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_3778),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_4495)
);

OR2x6_ASAP7_75t_L g4496 ( 
.A(n_3824),
.B(n_140),
.Y(n_4496)
);

INVx3_ASAP7_75t_L g4497 ( 
.A(n_3980),
.Y(n_4497)
);

OR2x2_ASAP7_75t_L g4498 ( 
.A(n_3906),
.B(n_140),
.Y(n_4498)
);

AND2x6_ASAP7_75t_L g4499 ( 
.A(n_3744),
.B(n_141),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_3590),
.Y(n_4500)
);

BUFx3_ASAP7_75t_L g4501 ( 
.A(n_3907),
.Y(n_4501)
);

AOI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_3870),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_3591),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3858),
.B(n_143),
.Y(n_4504)
);

A2O1A1Ixp33_ASAP7_75t_L g4505 ( 
.A1(n_3708),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_3594),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_3859),
.B(n_144),
.Y(n_4507)
);

BUFx6f_ASAP7_75t_L g4508 ( 
.A(n_3506),
.Y(n_4508)
);

INVxp67_ASAP7_75t_L g4509 ( 
.A(n_3916),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_3822),
.B(n_145),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_3797),
.B(n_145),
.Y(n_4511)
);

BUFx6f_ASAP7_75t_L g4512 ( 
.A(n_3500),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_3802),
.B(n_146),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_3889),
.B(n_3855),
.Y(n_4514)
);

INVx1_ASAP7_75t_SL g4515 ( 
.A(n_3990),
.Y(n_4515)
);

BUFx6f_ASAP7_75t_L g4516 ( 
.A(n_3505),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_3764),
.B(n_146),
.Y(n_4517)
);

AO22x1_ASAP7_75t_L g4518 ( 
.A1(n_3924),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_3599),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_3600),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_3604),
.Y(n_4521)
);

AND2x4_ASAP7_75t_L g4522 ( 
.A(n_3909),
.B(n_147),
.Y(n_4522)
);

INVx2_ASAP7_75t_SL g4523 ( 
.A(n_3825),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_3968),
.Y(n_4524)
);

INVx2_ASAP7_75t_SL g4525 ( 
.A(n_3827),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3970),
.Y(n_4526)
);

INVx4_ASAP7_75t_L g4527 ( 
.A(n_3593),
.Y(n_4527)
);

AND2x6_ASAP7_75t_L g4528 ( 
.A(n_3706),
.B(n_147),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_3834),
.B(n_148),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_3872),
.B(n_148),
.Y(n_4530)
);

NAND3xp33_ASAP7_75t_L g4531 ( 
.A(n_3607),
.B(n_149),
.C(n_150),
.Y(n_4531)
);

OR2x2_ASAP7_75t_SL g4532 ( 
.A(n_3715),
.B(n_150),
.Y(n_4532)
);

BUFx2_ASAP7_75t_L g4533 ( 
.A(n_3491),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_3508),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_3513),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_SL g4536 ( 
.A(n_3905),
.B(n_149),
.Y(n_4536)
);

INVx2_ASAP7_75t_SL g4537 ( 
.A(n_3878),
.Y(n_4537)
);

INVx3_ASAP7_75t_L g4538 ( 
.A(n_3941),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_3509),
.B(n_150),
.Y(n_4539)
);

HB1xp67_ASAP7_75t_L g4540 ( 
.A(n_3883),
.Y(n_4540)
);

OAI221xp5_ASAP7_75t_L g4541 ( 
.A1(n_3989),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_4541)
);

INVxp67_ASAP7_75t_L g4542 ( 
.A(n_3576),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_3514),
.Y(n_4543)
);

CKINVDCx5p33_ASAP7_75t_R g4544 ( 
.A(n_3587),
.Y(n_4544)
);

NOR3xp33_ASAP7_75t_SL g4545 ( 
.A(n_3815),
.B(n_151),
.C(n_152),
.Y(n_4545)
);

INVx2_ASAP7_75t_SL g4546 ( 
.A(n_3597),
.Y(n_4546)
);

AND2x4_ASAP7_75t_L g4547 ( 
.A(n_3915),
.B(n_151),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_3516),
.Y(n_4548)
);

BUFx3_ASAP7_75t_L g4549 ( 
.A(n_3763),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_3786),
.Y(n_4550)
);

CKINVDCx8_ASAP7_75t_R g4551 ( 
.A(n_3833),
.Y(n_4551)
);

AND2x2_ASAP7_75t_SL g4552 ( 
.A(n_3830),
.B(n_153),
.Y(n_4552)
);

HB1xp67_ASAP7_75t_L g4553 ( 
.A(n_3480),
.Y(n_4553)
);

NOR2x2_ASAP7_75t_L g4554 ( 
.A(n_3842),
.B(n_153),
.Y(n_4554)
);

AOI22xp33_ASAP7_75t_L g4555 ( 
.A1(n_3948),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_4555)
);

NAND2x1p5_ASAP7_75t_L g4556 ( 
.A(n_3767),
.B(n_3601),
.Y(n_4556)
);

INVx4_ASAP7_75t_L g4557 ( 
.A(n_3984),
.Y(n_4557)
);

A2O1A1Ixp33_ASAP7_75t_L g4558 ( 
.A1(n_3639),
.A2(n_158),
.B(n_155),
.C(n_156),
.Y(n_4558)
);

AOI22xp5_ASAP7_75t_L g4559 ( 
.A1(n_3619),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_3477),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_3873),
.B(n_3876),
.Y(n_4561)
);

INVx2_ASAP7_75t_SL g4562 ( 
.A(n_3992),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_3441),
.Y(n_4563)
);

BUFx8_ASAP7_75t_L g4564 ( 
.A(n_4071),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4191),
.A2(n_3643),
.B(n_3963),
.Y(n_4565)
);

AO21x1_ASAP7_75t_L g4566 ( 
.A1(n_4347),
.A2(n_3908),
.B(n_3640),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4089),
.B(n_3624),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4025),
.Y(n_4568)
);

NOR2xp33_ASAP7_75t_L g4569 ( 
.A(n_4415),
.B(n_3476),
.Y(n_4569)
);

BUFx3_ASAP7_75t_L g4570 ( 
.A(n_4069),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4044),
.Y(n_4571)
);

A2O1A1Ixp33_ASAP7_75t_L g4572 ( 
.A1(n_4066),
.A2(n_3862),
.B(n_3874),
.C(n_3837),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4300),
.A2(n_3937),
.B(n_3918),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4006),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_4091),
.B(n_3911),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4065),
.Y(n_4576)
);

NOR2x1_ASAP7_75t_L g4577 ( 
.A(n_4068),
.B(n_3943),
.Y(n_4577)
);

NAND2xp5_ASAP7_75t_L g4578 ( 
.A(n_4092),
.B(n_3955),
.Y(n_4578)
);

AOI21xp5_ASAP7_75t_L g4579 ( 
.A1(n_4314),
.A2(n_3969),
.B(n_3950),
.Y(n_4579)
);

AOI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4552),
.A2(n_3987),
.B1(n_3957),
.B2(n_3891),
.Y(n_4580)
);

OAI21xp5_ASAP7_75t_L g4581 ( 
.A1(n_4558),
.A2(n_4310),
.B(n_4531),
.Y(n_4581)
);

BUFx3_ASAP7_75t_L g4582 ( 
.A(n_4070),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_SL g4583 ( 
.A(n_4210),
.B(n_3650),
.Y(n_4583)
);

HB1xp67_ASAP7_75t_L g4584 ( 
.A(n_4103),
.Y(n_4584)
);

O2A1O1Ixp33_ASAP7_75t_SL g4585 ( 
.A1(n_4002),
.A2(n_3765),
.B(n_3893),
.C(n_3496),
.Y(n_4585)
);

BUFx6f_ASAP7_75t_L g4586 ( 
.A(n_4021),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4096),
.B(n_3732),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4053),
.A2(n_4100),
.B(n_4255),
.Y(n_4588)
);

AOI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4175),
.A2(n_3658),
.B(n_3612),
.Y(n_4589)
);

AOI21xp5_ASAP7_75t_L g4590 ( 
.A1(n_4176),
.A2(n_3686),
.B(n_3665),
.Y(n_4590)
);

NOR2xp33_ASAP7_75t_L g4591 ( 
.A(n_4014),
.B(n_4327),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4234),
.B(n_3877),
.Y(n_4592)
);

INVx2_ASAP7_75t_L g4593 ( 
.A(n_4080),
.Y(n_4593)
);

BUFx2_ASAP7_75t_L g4594 ( 
.A(n_4302),
.Y(n_4594)
);

OAI22xp5_ASAP7_75t_L g4595 ( 
.A1(n_4532),
.A2(n_3845),
.B1(n_3884),
.B2(n_3493),
.Y(n_4595)
);

BUFx8_ASAP7_75t_SL g4596 ( 
.A(n_4035),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_4186),
.A2(n_3689),
.B(n_3687),
.Y(n_4597)
);

AOI21xp5_ASAP7_75t_L g4598 ( 
.A1(n_4207),
.A2(n_3707),
.B(n_3690),
.Y(n_4598)
);

OAI22xp5_ASAP7_75t_L g4599 ( 
.A1(n_4048),
.A2(n_4030),
.B1(n_4210),
.B2(n_4441),
.Y(n_4599)
);

AOI21xp5_ASAP7_75t_L g4600 ( 
.A1(n_4211),
.A2(n_3759),
.B(n_3738),
.Y(n_4600)
);

AOI22xp5_ASAP7_75t_L g4601 ( 
.A1(n_4514),
.A2(n_3811),
.B1(n_3823),
.B2(n_3507),
.Y(n_4601)
);

AOI21xp5_ASAP7_75t_L g4602 ( 
.A1(n_4111),
.A2(n_3502),
.B(n_3448),
.Y(n_4602)
);

OR2x6_ASAP7_75t_L g4603 ( 
.A(n_4162),
.B(n_3471),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4131),
.B(n_159),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4081),
.Y(n_4605)
);

AOI21xp5_ASAP7_75t_L g4606 ( 
.A1(n_4125),
.A2(n_3789),
.B(n_3740),
.Y(n_4606)
);

NOR2xp33_ASAP7_75t_SL g4607 ( 
.A(n_4115),
.B(n_160),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4010),
.B(n_160),
.Y(n_4608)
);

OR2x6_ASAP7_75t_SL g4609 ( 
.A(n_4085),
.B(n_161),
.Y(n_4609)
);

OAI21x1_ASAP7_75t_L g4610 ( 
.A1(n_4386),
.A2(n_983),
.B(n_975),
.Y(n_4610)
);

A2O1A1Ixp33_ASAP7_75t_L g4611 ( 
.A1(n_4545),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_4611)
);

AOI21xp5_ASAP7_75t_L g4612 ( 
.A1(n_4127),
.A2(n_162),
.B(n_163),
.Y(n_4612)
);

NOR2x1_ASAP7_75t_L g4613 ( 
.A(n_4135),
.B(n_162),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_SL g4614 ( 
.A(n_4210),
.B(n_163),
.Y(n_4614)
);

OAI22xp5_ASAP7_75t_L g4615 ( 
.A1(n_4019),
.A2(n_4162),
.B1(n_4496),
.B2(n_4483),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_4183),
.A2(n_164),
.B(n_165),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4016),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4017),
.Y(n_4618)
);

O2A1O1Ixp33_ASAP7_75t_L g4619 ( 
.A1(n_4036),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_SL g4620 ( 
.A(n_4060),
.B(n_165),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4007),
.B(n_167),
.Y(n_4621)
);

AOI21x1_ASAP7_75t_L g4622 ( 
.A1(n_4183),
.A2(n_167),
.B(n_168),
.Y(n_4622)
);

AOI21xp5_ASAP7_75t_L g4623 ( 
.A1(n_4147),
.A2(n_168),
.B(n_169),
.Y(n_4623)
);

A2O1A1Ixp33_ASAP7_75t_L g4624 ( 
.A1(n_4275),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_4624)
);

NOR2xp67_ASAP7_75t_L g4625 ( 
.A(n_4107),
.B(n_170),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4013),
.B(n_170),
.Y(n_4626)
);

INVx2_ASAP7_75t_L g4627 ( 
.A(n_4087),
.Y(n_4627)
);

OAI21xp5_ASAP7_75t_L g4628 ( 
.A1(n_4505),
.A2(n_171),
.B(n_172),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_SL g4629 ( 
.A(n_4060),
.B(n_171),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4020),
.B(n_172),
.Y(n_4630)
);

O2A1O1Ixp33_ASAP7_75t_L g4631 ( 
.A1(n_4491),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4528),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_4632)
);

AOI21x1_ASAP7_75t_L g4633 ( 
.A1(n_4283),
.A2(n_174),
.B(n_176),
.Y(n_4633)
);

AOI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_4156),
.A2(n_176),
.B(n_177),
.Y(n_4634)
);

AND2x2_ASAP7_75t_L g4635 ( 
.A(n_4345),
.B(n_4072),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4090),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4026),
.B(n_176),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4027),
.Y(n_4638)
);

AO32x1_ASAP7_75t_L g4639 ( 
.A1(n_4349),
.A2(n_180),
.A3(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4052),
.B(n_177),
.Y(n_4640)
);

AOI21x1_ASAP7_75t_L g4641 ( 
.A1(n_4379),
.A2(n_178),
.B(n_180),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4198),
.Y(n_4642)
);

INVx1_ASAP7_75t_SL g4643 ( 
.A(n_4021),
.Y(n_4643)
);

AOI21xp5_ASAP7_75t_L g4644 ( 
.A1(n_4258),
.A2(n_178),
.B(n_181),
.Y(n_4644)
);

BUFx6f_ASAP7_75t_L g4645 ( 
.A(n_4039),
.Y(n_4645)
);

AOI21xp33_ASAP7_75t_L g4646 ( 
.A1(n_4252),
.A2(n_181),
.B(n_182),
.Y(n_4646)
);

BUFx12f_ASAP7_75t_L g4647 ( 
.A(n_4157),
.Y(n_4647)
);

INVx3_ASAP7_75t_L g4648 ( 
.A(n_4410),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4067),
.B(n_182),
.Y(n_4649)
);

OAI21xp33_ASAP7_75t_L g4650 ( 
.A1(n_4490),
.A2(n_183),
.B(n_184),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4075),
.B(n_4076),
.Y(n_4651)
);

AOI21xp5_ASAP7_75t_L g4652 ( 
.A1(n_4355),
.A2(n_183),
.B(n_184),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4077),
.B(n_183),
.Y(n_4653)
);

OAI22xp5_ASAP7_75t_L g4654 ( 
.A1(n_4483),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4196),
.B(n_4395),
.Y(n_4655)
);

AOI21xp5_ASAP7_75t_L g4656 ( 
.A1(n_4367),
.A2(n_186),
.B(n_187),
.Y(n_4656)
);

NOR2xp33_ASAP7_75t_L g4657 ( 
.A(n_4106),
.B(n_186),
.Y(n_4657)
);

AOI221xp5_ASAP7_75t_L g4658 ( 
.A1(n_4482),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_4658)
);

A2O1A1Ixp33_ASAP7_75t_L g4659 ( 
.A1(n_4408),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_4659)
);

INVx11_ASAP7_75t_L g4660 ( 
.A(n_4232),
.Y(n_4660)
);

AOI21xp5_ASAP7_75t_L g4661 ( 
.A1(n_4459),
.A2(n_188),
.B(n_191),
.Y(n_4661)
);

BUFx2_ASAP7_75t_L g4662 ( 
.A(n_4103),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4079),
.B(n_191),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4086),
.B(n_192),
.Y(n_4664)
);

INVx4_ASAP7_75t_L g4665 ( 
.A(n_4015),
.Y(n_4665)
);

AOI22xp5_ASAP7_75t_L g4666 ( 
.A1(n_4528),
.A2(n_4499),
.B1(n_4195),
.B2(n_4037),
.Y(n_4666)
);

OAI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4496),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_4667)
);

OAI21xp5_ASAP7_75t_L g4668 ( 
.A1(n_4471),
.A2(n_4393),
.B(n_4443),
.Y(n_4668)
);

AOI21xp5_ASAP7_75t_L g4669 ( 
.A1(n_4202),
.A2(n_193),
.B(n_194),
.Y(n_4669)
);

AOI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4386),
.A2(n_193),
.B(n_194),
.Y(n_4670)
);

OR2x2_ASAP7_75t_L g4671 ( 
.A(n_4478),
.B(n_195),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4097),
.B(n_195),
.Y(n_4672)
);

INVx2_ASAP7_75t_SL g4673 ( 
.A(n_4029),
.Y(n_4673)
);

OAI21x1_ASAP7_75t_L g4674 ( 
.A1(n_4137),
.A2(n_983),
.B(n_975),
.Y(n_4674)
);

INVx3_ASAP7_75t_L g4675 ( 
.A(n_4232),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4105),
.B(n_195),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4108),
.B(n_196),
.Y(n_4677)
);

INVx2_ASAP7_75t_SL g4678 ( 
.A(n_4047),
.Y(n_4678)
);

OAI21x1_ASAP7_75t_L g4679 ( 
.A1(n_4139),
.A2(n_986),
.B(n_977),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4123),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4428),
.A2(n_196),
.B(n_197),
.Y(n_4681)
);

INVx1_ASAP7_75t_SL g4682 ( 
.A(n_4403),
.Y(n_4682)
);

AOI21xp5_ASAP7_75t_L g4683 ( 
.A1(n_4433),
.A2(n_4149),
.B(n_4143),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4387),
.A2(n_197),
.B(n_198),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_SL g4685 ( 
.A(n_4060),
.B(n_4256),
.Y(n_4685)
);

AOI21x1_ASAP7_75t_L g4686 ( 
.A1(n_4050),
.A2(n_197),
.B(n_198),
.Y(n_4686)
);

AOI21xp5_ASAP7_75t_L g4687 ( 
.A1(n_4344),
.A2(n_4049),
.B(n_4333),
.Y(n_4687)
);

AOI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4230),
.A2(n_198),
.B(n_199),
.Y(n_4688)
);

AOI21xp5_ASAP7_75t_L g4689 ( 
.A1(n_4250),
.A2(n_199),
.B(n_200),
.Y(n_4689)
);

AOI21xp5_ASAP7_75t_L g4690 ( 
.A1(n_4296),
.A2(n_4322),
.B(n_4317),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4124),
.B(n_200),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4153),
.B(n_200),
.Y(n_4692)
);

AOI21xp33_ASAP7_75t_L g4693 ( 
.A1(n_4323),
.A2(n_201),
.B(n_202),
.Y(n_4693)
);

O2A1O1Ixp33_ASAP7_75t_L g4694 ( 
.A1(n_4561),
.A2(n_204),
.B(n_201),
.C(n_202),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4167),
.B(n_4171),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4326),
.A2(n_204),
.B(n_205),
.Y(n_4696)
);

NOR2xp33_ASAP7_75t_L g4697 ( 
.A(n_4141),
.B(n_204),
.Y(n_4697)
);

BUFx6f_ASAP7_75t_L g4698 ( 
.A(n_4249),
.Y(n_4698)
);

AOI21x1_ASAP7_75t_L g4699 ( 
.A1(n_4291),
.A2(n_205),
.B(n_206),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_SL g4700 ( 
.A(n_4060),
.B(n_205),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_SL g4701 ( 
.A(n_4256),
.B(n_206),
.Y(n_4701)
);

O2A1O1Ixp33_ASAP7_75t_L g4702 ( 
.A1(n_4336),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4434),
.B(n_207),
.Y(n_4703)
);

BUFx2_ASAP7_75t_SL g4704 ( 
.A(n_4160),
.Y(n_4704)
);

NAND2x1p5_ASAP7_75t_L g4705 ( 
.A(n_3998),
.B(n_207),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4177),
.B(n_208),
.Y(n_4706)
);

O2A1O1Ixp33_ASAP7_75t_L g4707 ( 
.A1(n_4332),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_4707)
);

NOR2xp33_ASAP7_75t_L g4708 ( 
.A(n_4217),
.B(n_210),
.Y(n_4708)
);

O2A1O1Ixp33_ASAP7_75t_L g4709 ( 
.A1(n_4442),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_4709)
);

INVx3_ASAP7_75t_L g4710 ( 
.A(n_4232),
.Y(n_4710)
);

BUFx6f_ASAP7_75t_L g4711 ( 
.A(n_4249),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4405),
.A2(n_211),
.B(n_212),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4179),
.Y(n_4713)
);

AO22x1_ASAP7_75t_L g4714 ( 
.A1(n_4256),
.A2(n_214),
.B1(n_211),
.B2(n_213),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4188),
.B(n_213),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_L g4716 ( 
.A(n_4200),
.B(n_213),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4206),
.Y(n_4717)
);

OAI22xp5_ASAP7_75t_L g4718 ( 
.A1(n_4432),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_4718)
);

BUFx2_ASAP7_75t_L g4719 ( 
.A(n_4159),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_SL g4720 ( 
.A(n_4298),
.B(n_214),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4201),
.Y(n_4721)
);

AOI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4528),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_4722)
);

AOI21xp5_ASAP7_75t_L g4723 ( 
.A1(n_4461),
.A2(n_216),
.B(n_217),
.Y(n_4723)
);

INVxp67_ASAP7_75t_L g4724 ( 
.A(n_4237),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4204),
.B(n_218),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_4064),
.Y(n_4726)
);

AOI221xp5_ASAP7_75t_L g4727 ( 
.A1(n_4420),
.A2(n_221),
.B1(n_218),
.B2(n_220),
.C(n_222),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4205),
.B(n_218),
.Y(n_4728)
);

AOI21xp5_ASAP7_75t_L g4729 ( 
.A1(n_4274),
.A2(n_220),
.B(n_221),
.Y(n_4729)
);

AOI21xp5_ASAP7_75t_L g4730 ( 
.A1(n_4226),
.A2(n_220),
.B(n_221),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_4059),
.A2(n_4164),
.B(n_4114),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4216),
.B(n_222),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_SL g4733 ( 
.A(n_4394),
.B(n_222),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4218),
.B(n_223),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4220),
.B(n_223),
.Y(n_4735)
);

OR2x2_ASAP7_75t_L g4736 ( 
.A(n_4478),
.B(n_223),
.Y(n_4736)
);

NOR2xp33_ASAP7_75t_L g4737 ( 
.A(n_4222),
.B(n_224),
.Y(n_4737)
);

INVx2_ASAP7_75t_L g4738 ( 
.A(n_4213),
.Y(n_4738)
);

AO32x1_ASAP7_75t_L g4739 ( 
.A1(n_4003),
.A2(n_226),
.A3(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_4739)
);

AOI21x1_ASAP7_75t_L g4740 ( 
.A1(n_4008),
.A2(n_4012),
.B(n_4009),
.Y(n_4740)
);

OAI22xp5_ASAP7_75t_L g4741 ( 
.A1(n_4460),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_4741)
);

AOI21xp5_ASAP7_75t_L g4742 ( 
.A1(n_4005),
.A2(n_226),
.B(n_228),
.Y(n_4742)
);

BUFx2_ASAP7_75t_SL g4743 ( 
.A(n_4028),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4221),
.B(n_228),
.Y(n_4744)
);

AOI21xp5_ASAP7_75t_L g4745 ( 
.A1(n_4368),
.A2(n_4165),
.B(n_4034),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4223),
.B(n_229),
.Y(n_4746)
);

INVx3_ASAP7_75t_L g4747 ( 
.A(n_4054),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4227),
.B(n_230),
.Y(n_4748)
);

AOI22xp5_ASAP7_75t_L g4749 ( 
.A1(n_4499),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_4749)
);

NAND3x1_ASAP7_75t_L g4750 ( 
.A(n_4011),
.B(n_231),
.C(n_232),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4238),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_4246),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4253),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4240),
.Y(n_4754)
);

CKINVDCx11_ASAP7_75t_R g4755 ( 
.A(n_4315),
.Y(n_4755)
);

AO21x1_ASAP7_75t_L g4756 ( 
.A1(n_4288),
.A2(n_231),
.B(n_232),
.Y(n_4756)
);

AOI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4398),
.A2(n_233),
.B(n_234),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_SL g4758 ( 
.A(n_4117),
.B(n_4129),
.Y(n_4758)
);

NOR2xp67_ASAP7_75t_L g4759 ( 
.A(n_4132),
.B(n_233),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4245),
.B(n_233),
.Y(n_4760)
);

AOI21xp5_ASAP7_75t_L g4761 ( 
.A1(n_4435),
.A2(n_234),
.B(n_235),
.Y(n_4761)
);

NOR2xp67_ASAP7_75t_L g4762 ( 
.A(n_4121),
.B(n_234),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4259),
.B(n_235),
.Y(n_4763)
);

BUFx6f_ASAP7_75t_L g4764 ( 
.A(n_4182),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4266),
.B(n_235),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_SL g4766 ( 
.A(n_4138),
.B(n_236),
.Y(n_4766)
);

AO21x2_ASAP7_75t_L g4767 ( 
.A1(n_4022),
.A2(n_236),
.B(n_237),
.Y(n_4767)
);

BUFx6f_ASAP7_75t_L g4768 ( 
.A(n_4182),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4439),
.B(n_236),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4435),
.A2(n_237),
.B(n_238),
.Y(n_4770)
);

AOI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4329),
.A2(n_237),
.B(n_239),
.Y(n_4771)
);

BUFx12f_ASAP7_75t_L g4772 ( 
.A(n_4130),
.Y(n_4772)
);

O2A1O1Ixp33_ASAP7_75t_L g4773 ( 
.A1(n_4542),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4277),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_4134),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_4446),
.B(n_239),
.Y(n_4776)
);

AOI22xp5_ASAP7_75t_L g4777 ( 
.A1(n_4499),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4282),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4385),
.A2(n_240),
.B(n_242),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4284),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4297),
.B(n_242),
.Y(n_4781)
);

BUFx12f_ASAP7_75t_L g4782 ( 
.A(n_4101),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4267),
.Y(n_4783)
);

AOI21xp5_ASAP7_75t_L g4784 ( 
.A1(n_4382),
.A2(n_243),
.B(n_244),
.Y(n_4784)
);

BUFx6f_ASAP7_75t_L g4785 ( 
.A(n_4098),
.Y(n_4785)
);

INVxp67_ASAP7_75t_L g4786 ( 
.A(n_4088),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_SL g4787 ( 
.A(n_4055),
.B(n_243),
.Y(n_4787)
);

INVxp33_ASAP7_75t_SL g4788 ( 
.A(n_4161),
.Y(n_4788)
);

A2O1A1Ixp33_ASAP7_75t_L g4789 ( 
.A1(n_4180),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4299),
.B(n_244),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4306),
.B(n_245),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4038),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4145),
.B(n_245),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4382),
.A2(n_4354),
.B(n_4350),
.Y(n_4794)
);

INVxp67_ASAP7_75t_L g4795 ( 
.A(n_4163),
.Y(n_4795)
);

O2A1O1Ixp33_ASAP7_75t_SL g4796 ( 
.A1(n_4045),
.A2(n_4018),
.B(n_4494),
.C(n_4477),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_SL g4797 ( 
.A(n_4330),
.B(n_4148),
.Y(n_4797)
);

INVx11_ASAP7_75t_L g4798 ( 
.A(n_4287),
.Y(n_4798)
);

AOI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4546),
.A2(n_246),
.B(n_247),
.Y(n_4799)
);

AOI21xp5_ASAP7_75t_L g4800 ( 
.A1(n_4212),
.A2(n_246),
.B(n_247),
.Y(n_4800)
);

BUFx2_ASAP7_75t_L g4801 ( 
.A(n_4287),
.Y(n_4801)
);

INVx1_ASAP7_75t_SL g4802 ( 
.A(n_4078),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_SL g4803 ( 
.A(n_4290),
.B(n_248),
.Y(n_4803)
);

BUFx3_ASAP7_75t_L g4804 ( 
.A(n_4024),
.Y(n_4804)
);

AO21x1_ASAP7_75t_L g4805 ( 
.A1(n_4527),
.A2(n_248),
.B(n_249),
.Y(n_4805)
);

BUFx6f_ASAP7_75t_L g4806 ( 
.A(n_4098),
.Y(n_4806)
);

OA21x2_ASAP7_75t_L g4807 ( 
.A1(n_4004),
.A2(n_248),
.B(n_250),
.Y(n_4807)
);

AOI21xp33_ASAP7_75t_L g4808 ( 
.A1(n_4523),
.A2(n_250),
.B(n_251),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4404),
.B(n_4406),
.Y(n_4809)
);

AOI33xp33_ASAP7_75t_L g4810 ( 
.A1(n_4462),
.A2(n_252),
.A3(n_254),
.B1(n_250),
.B2(n_251),
.B3(n_253),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4319),
.Y(n_4811)
);

AOI21xp5_ASAP7_75t_L g4812 ( 
.A1(n_4212),
.A2(n_253),
.B(n_254),
.Y(n_4812)
);

CKINVDCx6p67_ASAP7_75t_R g4813 ( 
.A(n_4199),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_SL g4814 ( 
.A(n_4353),
.B(n_253),
.Y(n_4814)
);

AOI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4353),
.A2(n_254),
.B(n_255),
.Y(n_4815)
);

AOI21xp5_ASAP7_75t_L g4816 ( 
.A1(n_4375),
.A2(n_255),
.B(n_256),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4402),
.B(n_256),
.Y(n_4817)
);

OAI22xp5_ASAP7_75t_L g4818 ( 
.A1(n_4293),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_SL g4819 ( 
.A(n_4375),
.B(n_257),
.Y(n_4819)
);

AOI21xp5_ASAP7_75t_L g4820 ( 
.A1(n_4372),
.A2(n_257),
.B(n_258),
.Y(n_4820)
);

AND2x2_ASAP7_75t_L g4821 ( 
.A(n_4122),
.B(n_259),
.Y(n_4821)
);

AND2x2_ASAP7_75t_L g4822 ( 
.A(n_4364),
.B(n_260),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4417),
.B(n_4422),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4040),
.Y(n_4824)
);

NOR2xp33_ASAP7_75t_L g4825 ( 
.A(n_4378),
.B(n_260),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4251),
.Y(n_4826)
);

AND2x4_ASAP7_75t_L g4827 ( 
.A(n_4287),
.B(n_260),
.Y(n_4827)
);

BUFx2_ASAP7_75t_L g4828 ( 
.A(n_4348),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_L g4829 ( 
.A(n_4423),
.B(n_261),
.Y(n_4829)
);

OAI21xp5_ASAP7_75t_L g4830 ( 
.A1(n_4559),
.A2(n_261),
.B(n_262),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4424),
.B(n_261),
.Y(n_4831)
);

BUFx2_ASAP7_75t_L g4832 ( 
.A(n_4451),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4099),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4437),
.B(n_262),
.Y(n_4834)
);

O2A1O1Ixp33_ASAP7_75t_L g4835 ( 
.A1(n_4140),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4533),
.A2(n_4190),
.B1(n_4551),
.B2(n_4057),
.Y(n_4836)
);

OAI22xp5_ASAP7_75t_L g4837 ( 
.A1(n_4533),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_4837)
);

NOR2xp33_ASAP7_75t_L g4838 ( 
.A(n_4110),
.B(n_265),
.Y(n_4838)
);

O2A1O1Ixp33_ASAP7_75t_L g4839 ( 
.A1(n_4540),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_4839)
);

HB1xp67_ASAP7_75t_L g4840 ( 
.A(n_4219),
.Y(n_4840)
);

NOR2xp33_ASAP7_75t_L g4841 ( 
.A(n_4214),
.B(n_267),
.Y(n_4841)
);

INVxp33_ASAP7_75t_SL g4842 ( 
.A(n_4151),
.Y(n_4842)
);

HB1xp67_ASAP7_75t_L g4843 ( 
.A(n_4447),
.Y(n_4843)
);

AOI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_4396),
.A2(n_267),
.B(n_268),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4440),
.B(n_4445),
.Y(n_4845)
);

BUFx3_ASAP7_75t_L g4846 ( 
.A(n_4024),
.Y(n_4846)
);

NAND3xp33_ASAP7_75t_L g4847 ( 
.A(n_4455),
.B(n_269),
.C(n_270),
.Y(n_4847)
);

AOI21xp5_ASAP7_75t_L g4848 ( 
.A1(n_4396),
.A2(n_4411),
.B(n_4264),
.Y(n_4848)
);

CKINVDCx5p33_ASAP7_75t_R g4849 ( 
.A(n_4225),
.Y(n_4849)
);

A2O1A1Ixp33_ASAP7_75t_L g4850 ( 
.A1(n_4318),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4454),
.B(n_270),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4411),
.A2(n_271),
.B(n_272),
.Y(n_4852)
);

BUFx8_ASAP7_75t_L g4853 ( 
.A(n_4078),
.Y(n_4853)
);

HB1xp67_ASAP7_75t_L g4854 ( 
.A(n_4397),
.Y(n_4854)
);

OR2x6_ASAP7_75t_L g4855 ( 
.A(n_4294),
.B(n_271),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4338),
.Y(n_4856)
);

AO22x1_ASAP7_75t_L g4857 ( 
.A1(n_4239),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_4857)
);

O2A1O1Ixp33_ASAP7_75t_L g4858 ( 
.A1(n_4166),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_4858)
);

A2O1A1Ixp33_ASAP7_75t_L g4859 ( 
.A1(n_4493),
.A2(n_276),
.B(n_273),
.C(n_274),
.Y(n_4859)
);

OAI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_4553),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_4860)
);

O2A1O1Ixp33_ASAP7_75t_L g4861 ( 
.A1(n_4412),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_4861)
);

O2A1O1Ixp33_ASAP7_75t_L g4862 ( 
.A1(n_4416),
.A2(n_4247),
.B(n_4517),
.C(n_4549),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4458),
.B(n_279),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4466),
.B(n_279),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4251),
.Y(n_4865)
);

OAI21xp5_ASAP7_75t_L g4866 ( 
.A1(n_4470),
.A2(n_280),
.B(n_281),
.Y(n_4866)
);

NAND2x1p5_ASAP7_75t_L g4867 ( 
.A(n_4033),
.B(n_280),
.Y(n_4867)
);

AND2x4_ASAP7_75t_L g4868 ( 
.A(n_4095),
.B(n_280),
.Y(n_4868)
);

NAND2x1p5_ASAP7_75t_L g4869 ( 
.A(n_4033),
.B(n_281),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4474),
.B(n_282),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4476),
.B(n_282),
.Y(n_4871)
);

OAI22xp5_ASAP7_75t_L g4872 ( 
.A1(n_4280),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4309),
.Y(n_4873)
);

AO32x1_ASAP7_75t_L g4874 ( 
.A1(n_4557),
.A2(n_285),
.A3(n_283),
.B1(n_284),
.B2(n_286),
.Y(n_4874)
);

O2A1O1Ixp33_ASAP7_75t_L g4875 ( 
.A1(n_4465),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4312),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4479),
.B(n_285),
.Y(n_4877)
);

O2A1O1Ixp33_ASAP7_75t_L g4878 ( 
.A1(n_4511),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_L g4879 ( 
.A(n_4000),
.B(n_4544),
.Y(n_4879)
);

AND2x2_ASAP7_75t_L g4880 ( 
.A(n_4104),
.B(n_287),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4235),
.B(n_288),
.Y(n_4881)
);

OAI21xp33_ASAP7_75t_L g4882 ( 
.A1(n_4374),
.A2(n_4529),
.B(n_4513),
.Y(n_4882)
);

CKINVDCx6p67_ASAP7_75t_R g4883 ( 
.A(n_4119),
.Y(n_4883)
);

OAI22xp5_ASAP7_75t_L g4884 ( 
.A1(n_4292),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_4884)
);

AO21x1_ASAP7_75t_L g4885 ( 
.A1(n_4522),
.A2(n_289),
.B(n_290),
.Y(n_4885)
);

AOI21xp5_ASAP7_75t_L g4886 ( 
.A1(n_4308),
.A2(n_289),
.B(n_290),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4236),
.B(n_291),
.Y(n_4887)
);

AOI21x1_ASAP7_75t_L g4888 ( 
.A1(n_4093),
.A2(n_291),
.B(n_292),
.Y(n_4888)
);

A2O1A1Ixp33_ASAP7_75t_L g4889 ( 
.A1(n_4311),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_4889)
);

NOR2xp33_ASAP7_75t_L g4890 ( 
.A(n_4133),
.B(n_4056),
.Y(n_4890)
);

NOR2xp67_ASAP7_75t_SL g4891 ( 
.A(n_4320),
.B(n_292),
.Y(n_4891)
);

AOI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4341),
.A2(n_293),
.B(n_294),
.Y(n_4892)
);

AO22x1_ASAP7_75t_L g4893 ( 
.A1(n_4550),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4893)
);

AOI21xp5_ASAP7_75t_L g4894 ( 
.A1(n_4343),
.A2(n_295),
.B(n_296),
.Y(n_4894)
);

O2A1O1Ixp33_ASAP7_75t_SL g4895 ( 
.A1(n_4203),
.A2(n_297),
.B(n_295),
.C(n_296),
.Y(n_4895)
);

INVx4_ASAP7_75t_L g4896 ( 
.A(n_4320),
.Y(n_4896)
);

A2O1A1Ixp33_ASAP7_75t_L g4897 ( 
.A1(n_4328),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_4897)
);

AOI21xp5_ASAP7_75t_L g4898 ( 
.A1(n_4362),
.A2(n_298),
.B(n_300),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4480),
.B(n_300),
.Y(n_4899)
);

INVx4_ASAP7_75t_L g4900 ( 
.A(n_4320),
.Y(n_4900)
);

O2A1O1Ixp33_ASAP7_75t_L g4901 ( 
.A1(n_4481),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_L g4902 ( 
.A(n_4488),
.B(n_301),
.Y(n_4902)
);

AOI21xp33_ASAP7_75t_L g4903 ( 
.A1(n_4525),
.A2(n_4537),
.B(n_4562),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4500),
.B(n_301),
.Y(n_4904)
);

NAND2xp5_ASAP7_75t_L g4905 ( 
.A(n_4521),
.B(n_303),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_3999),
.B(n_303),
.Y(n_4906)
);

AOI21x1_ASAP7_75t_L g4907 ( 
.A1(n_4093),
.A2(n_304),
.B(n_305),
.Y(n_4907)
);

NOR3xp33_ASAP7_75t_L g4908 ( 
.A(n_4228),
.B(n_312),
.C(n_304),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4001),
.B(n_304),
.Y(n_4909)
);

INVx2_ASAP7_75t_L g4910 ( 
.A(n_4356),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4468),
.B(n_305),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4497),
.B(n_305),
.Y(n_4912)
);

AOI21xp5_ASAP7_75t_L g4913 ( 
.A1(n_4362),
.A2(n_306),
.B(n_307),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4335),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4361),
.Y(n_4915)
);

AOI21xp5_ASAP7_75t_L g4916 ( 
.A1(n_4334),
.A2(n_306),
.B(n_307),
.Y(n_4916)
);

OAI22xp5_ASAP7_75t_L g4917 ( 
.A1(n_4337),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4342),
.B(n_4358),
.Y(n_4918)
);

NOR2xp33_ASAP7_75t_L g4919 ( 
.A(n_4041),
.B(n_308),
.Y(n_4919)
);

CKINVDCx5p33_ASAP7_75t_R g4920 ( 
.A(n_4233),
.Y(n_4920)
);

INVx2_ASAP7_75t_L g4921 ( 
.A(n_4373),
.Y(n_4921)
);

BUFx6f_ASAP7_75t_L g4922 ( 
.A(n_4098),
.Y(n_4922)
);

AOI22xp5_ASAP7_75t_L g4923 ( 
.A1(n_4062),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_4923)
);

NOR2x1_ASAP7_75t_L g4924 ( 
.A(n_4421),
.B(n_309),
.Y(n_4924)
);

INVx1_ASAP7_75t_SL g4925 ( 
.A(n_4084),
.Y(n_4925)
);

NOR2xp67_ASAP7_75t_L g4926 ( 
.A(n_4209),
.B(n_310),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4369),
.B(n_311),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4538),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_4928)
);

BUFx6f_ASAP7_75t_L g4929 ( 
.A(n_4102),
.Y(n_4929)
);

A2O1A1Ixp33_ASAP7_75t_L g4930 ( 
.A1(n_4357),
.A2(n_314),
.B(n_311),
.C(n_313),
.Y(n_4930)
);

AOI22xp33_ASAP7_75t_L g4931 ( 
.A1(n_4489),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_4931)
);

OAI22xp5_ASAP7_75t_L g4932 ( 
.A1(n_4463),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_4932)
);

OAI21x1_ASAP7_75t_L g4933 ( 
.A1(n_4042),
.A2(n_982),
.B(n_973),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4370),
.B(n_315),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4371),
.B(n_316),
.Y(n_4935)
);

OAI21xp5_ASAP7_75t_L g4936 ( 
.A1(n_4279),
.A2(n_4555),
.B(n_4536),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4376),
.B(n_317),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4321),
.A2(n_317),
.B(n_318),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4381),
.Y(n_4939)
);

NOR2xp33_ASAP7_75t_L g4940 ( 
.A(n_4427),
.B(n_317),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4383),
.Y(n_4941)
);

NOR2xp33_ASAP7_75t_R g4942 ( 
.A(n_4181),
.B(n_318),
.Y(n_4942)
);

O2A1O1Ixp33_ASAP7_75t_L g4943 ( 
.A1(n_4485),
.A2(n_4504),
.B(n_4507),
.C(n_4524),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4031),
.B(n_4456),
.Y(n_4944)
);

NOR2xp33_ASAP7_75t_L g4945 ( 
.A(n_4083),
.B(n_4257),
.Y(n_4945)
);

AOI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4321),
.A2(n_319),
.B(n_320),
.Y(n_4946)
);

NOR2xp33_ASAP7_75t_L g4947 ( 
.A(n_4269),
.B(n_319),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4384),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4515),
.B(n_319),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_SL g4950 ( 
.A(n_4436),
.B(n_320),
.Y(n_4950)
);

NOR2xp33_ASAP7_75t_L g4951 ( 
.A(n_4158),
.B(n_321),
.Y(n_4951)
);

AOI22xp33_ASAP7_75t_L g4952 ( 
.A1(n_4501),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_4952)
);

O2A1O1Ixp33_ASAP7_75t_L g4953 ( 
.A1(n_4526),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_4953)
);

INVx3_ASAP7_75t_L g4954 ( 
.A(n_4023),
.Y(n_4954)
);

OAI21xp33_ASAP7_75t_L g4955 ( 
.A1(n_4449),
.A2(n_4450),
.B(n_4530),
.Y(n_4955)
);

AO22x1_ASAP7_75t_L g4956 ( 
.A1(n_4023),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4389),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_SL g4958 ( 
.A(n_4351),
.B(n_324),
.Y(n_4958)
);

AOI21x1_ASAP7_75t_L g4959 ( 
.A1(n_4352),
.A2(n_325),
.B(n_326),
.Y(n_4959)
);

NOR3xp33_ASAP7_75t_L g4960 ( 
.A(n_4448),
.B(n_333),
.C(n_325),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4400),
.Y(n_4961)
);

AOI21xp5_ASAP7_75t_L g4962 ( 
.A1(n_4095),
.A2(n_325),
.B(n_326),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4113),
.A2(n_326),
.B(n_327),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4487),
.B(n_327),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4429),
.Y(n_4965)
);

A2O1A1Ixp33_ASAP7_75t_L g4966 ( 
.A1(n_4391),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_4966)
);

O2A1O1Ixp33_ASAP7_75t_L g4967 ( 
.A1(n_4509),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_4967)
);

NOR2xp33_ASAP7_75t_L g4968 ( 
.A(n_4224),
.B(n_4243),
.Y(n_4968)
);

OR2x6_ASAP7_75t_SL g4969 ( 
.A(n_4263),
.B(n_4265),
.Y(n_4969)
);

AOI21x1_ASAP7_75t_L g4970 ( 
.A1(n_4352),
.A2(n_4113),
.B(n_4518),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4438),
.Y(n_4971)
);

O2A1O1Ixp33_ASAP7_75t_L g4972 ( 
.A1(n_4418),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4503),
.B(n_4506),
.Y(n_4973)
);

OAI22xp5_ASAP7_75t_L g4974 ( 
.A1(n_4294),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_4974)
);

OAI21xp33_ASAP7_75t_L g4975 ( 
.A1(n_4510),
.A2(n_4419),
.B(n_4475),
.Y(n_4975)
);

NOR2xp33_ASAP7_75t_L g4976 ( 
.A(n_4281),
.B(n_331),
.Y(n_4976)
);

OR2x6_ASAP7_75t_SL g4977 ( 
.A(n_4554),
.B(n_331),
.Y(n_4977)
);

AOI21x1_ASAP7_75t_L g4978 ( 
.A1(n_4360),
.A2(n_332),
.B(n_334),
.Y(n_4978)
);

INVx4_ASAP7_75t_L g4979 ( 
.A(n_4351),
.Y(n_4979)
);

INVx2_ASAP7_75t_L g4980 ( 
.A(n_4444),
.Y(n_4980)
);

OAI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4495),
.A2(n_335),
.B1(n_332),
.B2(n_334),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4094),
.Y(n_4982)
);

O2A1O1Ixp33_ASAP7_75t_L g4983 ( 
.A1(n_4254),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_4983)
);

AOI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_4563),
.A2(n_335),
.B(n_337),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4116),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4260),
.A2(n_337),
.B(n_338),
.Y(n_4986)
);

A2O1A1Ixp33_ASAP7_75t_L g4987 ( 
.A1(n_4325),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_4987)
);

A2O1A1Ixp33_ASAP7_75t_L g4988 ( 
.A1(n_4380),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_4988)
);

AOI22x1_ASAP7_75t_L g4989 ( 
.A1(n_4556),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4464),
.B(n_340),
.Y(n_4990)
);

AOI21xp5_ASAP7_75t_L g4991 ( 
.A1(n_4360),
.A2(n_341),
.B(n_342),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4120),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4126),
.Y(n_4993)
);

OAI22xp5_ASAP7_75t_SL g4994 ( 
.A1(n_4051),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_4994)
);

AOI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4289),
.A2(n_342),
.B(n_343),
.Y(n_4995)
);

AOI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4303),
.A2(n_344),
.B(n_345),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4519),
.B(n_345),
.Y(n_4997)
);

AOI21xp5_ASAP7_75t_L g4998 ( 
.A1(n_4304),
.A2(n_346),
.B(n_347),
.Y(n_4998)
);

AOI22xp33_ASAP7_75t_L g4999 ( 
.A1(n_4539),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_4999)
);

AOI33xp33_ASAP7_75t_L g5000 ( 
.A1(n_4430),
.A2(n_348),
.A3(n_350),
.B1(n_346),
.B2(n_347),
.B3(n_349),
.Y(n_5000)
);

O2A1O1Ixp33_ASAP7_75t_L g5001 ( 
.A1(n_4229),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_5001)
);

AOI21xp5_ASAP7_75t_L g5002 ( 
.A1(n_4305),
.A2(n_349),
.B(n_350),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4520),
.B(n_352),
.Y(n_5003)
);

OAI22xp5_ASAP7_75t_L g5004 ( 
.A1(n_4548),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_5004)
);

AOI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_4363),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_4128),
.Y(n_5006)
);

AOI21xp5_ASAP7_75t_L g5007 ( 
.A1(n_4316),
.A2(n_355),
.B(n_356),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_SL g5008 ( 
.A(n_4351),
.B(n_355),
.Y(n_5008)
);

AND2x6_ASAP7_75t_SL g5009 ( 
.A(n_4215),
.B(n_356),
.Y(n_5009)
);

AOI21xp5_ASAP7_75t_L g5010 ( 
.A1(n_4136),
.A2(n_357),
.B(n_358),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4146),
.Y(n_5011)
);

AOI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4154),
.A2(n_357),
.B(n_358),
.Y(n_5012)
);

BUFx8_ASAP7_75t_L g5013 ( 
.A(n_4058),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_L g5014 ( 
.A(n_4452),
.B(n_359),
.Y(n_5014)
);

INVx2_ASAP7_75t_SL g5015 ( 
.A(n_4192),
.Y(n_5015)
);

AOI22xp5_ASAP7_75t_L g5016 ( 
.A1(n_4560),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_5016)
);

INVx3_ASAP7_75t_L g5017 ( 
.A(n_4023),
.Y(n_5017)
);

BUFx4f_ASAP7_75t_L g5018 ( 
.A(n_4215),
.Y(n_5018)
);

AOI21xp5_ASAP7_75t_L g5019 ( 
.A1(n_4172),
.A2(n_360),
.B(n_361),
.Y(n_5019)
);

BUFx6f_ASAP7_75t_L g5020 ( 
.A(n_4102),
.Y(n_5020)
);

INVx2_ASAP7_75t_L g5021 ( 
.A(n_4174),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4185),
.Y(n_5022)
);

NOR2xp33_ASAP7_75t_L g5023 ( 
.A(n_4295),
.B(n_360),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4453),
.B(n_361),
.Y(n_5024)
);

AOI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4469),
.A2(n_362),
.B(n_363),
.Y(n_5025)
);

OA22x2_ASAP7_75t_L g5026 ( 
.A1(n_4109),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_5026)
);

AND2x6_ASAP7_75t_L g5027 ( 
.A(n_4063),
.B(n_364),
.Y(n_5027)
);

AOI22xp33_ASAP7_75t_L g5028 ( 
.A1(n_4541),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_5028)
);

AOI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4484),
.A2(n_365),
.B(n_366),
.Y(n_5029)
);

O2A1O1Ixp33_ASAP7_75t_L g5030 ( 
.A1(n_4261),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4486),
.A2(n_367),
.B(n_368),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_SL g5032 ( 
.A(n_4365),
.B(n_367),
.Y(n_5032)
);

INVx2_ASAP7_75t_SL g5033 ( 
.A(n_4032),
.Y(n_5033)
);

AOI21x1_ASAP7_75t_L g5034 ( 
.A1(n_4063),
.A2(n_368),
.B(n_369),
.Y(n_5034)
);

NOR2x1p5_ASAP7_75t_SL g5035 ( 
.A(n_4534),
.B(n_969),
.Y(n_5035)
);

AOI21xp5_ASAP7_75t_L g5036 ( 
.A1(n_4473),
.A2(n_369),
.B(n_370),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4473),
.A2(n_370),
.B(n_371),
.Y(n_5037)
);

O2A1O1Ixp33_ASAP7_75t_L g5038 ( 
.A1(n_4208),
.A2(n_372),
.B(n_370),
.C(n_371),
.Y(n_5038)
);

OAI21x1_ASAP7_75t_L g5039 ( 
.A1(n_4683),
.A2(n_4340),
.B(n_4286),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4588),
.A2(n_4473),
.B(n_4359),
.Y(n_5040)
);

HB1xp67_ASAP7_75t_L g5041 ( 
.A(n_4662),
.Y(n_5041)
);

AOI22xp5_ASAP7_75t_L g5042 ( 
.A1(n_4615),
.A2(n_4231),
.B1(n_4547),
.B2(n_4522),
.Y(n_5042)
);

AND2x4_ASAP7_75t_L g5043 ( 
.A(n_4594),
.B(n_4278),
.Y(n_5043)
);

AOI21xp5_ASAP7_75t_L g5044 ( 
.A1(n_4573),
.A2(n_4425),
.B(n_4390),
.Y(n_5044)
);

AO31x2_ASAP7_75t_L g5045 ( 
.A1(n_4566),
.A2(n_4399),
.A3(n_4426),
.B(n_4535),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4579),
.A2(n_4407),
.B(n_4365),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_SL g5047 ( 
.A(n_4645),
.B(n_4365),
.Y(n_5047)
);

OAI21x1_ASAP7_75t_L g5048 ( 
.A1(n_4565),
.A2(n_4346),
.B(n_4331),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4568),
.Y(n_5049)
);

BUFx6f_ASAP7_75t_L g5050 ( 
.A(n_4764),
.Y(n_5050)
);

NOR2xp33_ASAP7_75t_L g5051 ( 
.A(n_4643),
.B(n_4339),
.Y(n_5051)
);

A2O1A1Ixp33_ASAP7_75t_L g5052 ( 
.A1(n_4625),
.A2(n_4759),
.B(n_4926),
.C(n_4908),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4574),
.Y(n_5053)
);

OR2x6_ASAP7_75t_L g5054 ( 
.A(n_4719),
.B(n_4285),
.Y(n_5054)
);

OAI21x1_ASAP7_75t_L g5055 ( 
.A1(n_4740),
.A2(n_4388),
.B(n_4046),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4617),
.Y(n_5056)
);

OAI21x1_ASAP7_75t_SL g5057 ( 
.A1(n_4665),
.A2(n_4082),
.B(n_4061),
.Y(n_5057)
);

AOI21xp5_ASAP7_75t_L g5058 ( 
.A1(n_4685),
.A2(n_4457),
.B(n_4407),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4792),
.B(n_4543),
.Y(n_5059)
);

NOR2xp33_ASAP7_75t_L g5060 ( 
.A(n_4802),
.B(n_4170),
.Y(n_5060)
);

AND2x4_ASAP7_75t_L g5061 ( 
.A(n_4665),
.B(n_4407),
.Y(n_5061)
);

AOI21xp5_ASAP7_75t_L g5062 ( 
.A1(n_4687),
.A2(n_4457),
.B(n_4073),
.Y(n_5062)
);

OAI22xp5_ASAP7_75t_L g5063 ( 
.A1(n_4977),
.A2(n_4547),
.B1(n_4502),
.B2(n_4193),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4824),
.B(n_4173),
.Y(n_5064)
);

OAI22xp5_ASAP7_75t_L g5065 ( 
.A1(n_4666),
.A2(n_4472),
.B1(n_4498),
.B2(n_4467),
.Y(n_5065)
);

AOI21x1_ASAP7_75t_L g5066 ( 
.A1(n_4888),
.A2(n_4073),
.B(n_4168),
.Y(n_5066)
);

BUFx3_ASAP7_75t_L g5067 ( 
.A(n_4647),
.Y(n_5067)
);

INVx2_ASAP7_75t_SL g5068 ( 
.A(n_4853),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4973),
.B(n_4873),
.Y(n_5069)
);

AOI21x1_ASAP7_75t_SL g5070 ( 
.A1(n_4827),
.A2(n_4431),
.B(n_4150),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4618),
.Y(n_5071)
);

A2O1A1Ixp33_ASAP7_75t_L g5072 ( 
.A1(n_4611),
.A2(n_4144),
.B(n_4313),
.C(n_4043),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_4876),
.B(n_4413),
.Y(n_5073)
);

AOI211x1_ASAP7_75t_L g5074 ( 
.A1(n_4857),
.A2(n_4197),
.B(n_4074),
.C(n_4194),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_L g5075 ( 
.A(n_4914),
.B(n_4377),
.Y(n_5075)
);

AOI21x1_ASAP7_75t_L g5076 ( 
.A1(n_4907),
.A2(n_4169),
.B(n_4168),
.Y(n_5076)
);

OAI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_4847),
.A2(n_4142),
.B(n_4262),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_4939),
.B(n_4169),
.Y(n_5078)
);

A2O1A1Ixp33_ASAP7_75t_L g5079 ( 
.A1(n_4924),
.A2(n_4043),
.B(n_4118),
.C(n_4178),
.Y(n_5079)
);

AOI21xp33_ASAP7_75t_L g5080 ( 
.A1(n_4862),
.A2(n_4301),
.B(n_4270),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4638),
.Y(n_5081)
);

O2A1O1Ixp5_ASAP7_75t_L g5082 ( 
.A1(n_4956),
.A2(n_4118),
.B(n_4272),
.C(n_4268),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4680),
.Y(n_5083)
);

INVx2_ASAP7_75t_SL g5084 ( 
.A(n_4853),
.Y(n_5084)
);

A2O1A1Ixp33_ASAP7_75t_L g5085 ( 
.A1(n_4607),
.A2(n_4187),
.B(n_4189),
.C(n_4178),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4948),
.B(n_4187),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_4713),
.B(n_4189),
.Y(n_5087)
);

AND2x2_ASAP7_75t_L g5088 ( 
.A(n_4635),
.B(n_4244),
.Y(n_5088)
);

INVx2_ASAP7_75t_L g5089 ( 
.A(n_4571),
.Y(n_5089)
);

BUFx2_ASAP7_75t_L g5090 ( 
.A(n_4764),
.Y(n_5090)
);

INVx1_ASAP7_75t_SL g5091 ( 
.A(n_4704),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4721),
.B(n_4244),
.Y(n_5092)
);

AOI21x1_ASAP7_75t_L g5093 ( 
.A1(n_4970),
.A2(n_4155),
.B(n_4152),
.Y(n_5093)
);

AND2x2_ASAP7_75t_L g5094 ( 
.A(n_4944),
.B(n_4271),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_4751),
.Y(n_5095)
);

A2O1A1Ixp33_ASAP7_75t_L g5096 ( 
.A1(n_5000),
.A2(n_4271),
.B(n_4155),
.C(n_4152),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_L g5097 ( 
.A(n_4754),
.B(n_4276),
.Y(n_5097)
);

OR2x2_ASAP7_75t_L g5098 ( 
.A(n_4584),
.B(n_4324),
.Y(n_5098)
);

BUFx2_ASAP7_75t_L g5099 ( 
.A(n_4764),
.Y(n_5099)
);

A2O1A1Ixp33_ASAP7_75t_L g5100 ( 
.A1(n_4810),
.A2(n_4241),
.B(n_4242),
.C(n_4324),
.Y(n_5100)
);

AOI21x1_ASAP7_75t_SL g5101 ( 
.A1(n_4827),
.A2(n_4248),
.B(n_4457),
.Y(n_5101)
);

AOI21x1_ASAP7_75t_SL g5102 ( 
.A1(n_4868),
.A2(n_372),
.B(n_373),
.Y(n_5102)
);

AOI21xp5_ASAP7_75t_SL g5103 ( 
.A1(n_4599),
.A2(n_4733),
.B(n_4741),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4774),
.B(n_4492),
.Y(n_5104)
);

AND2x2_ASAP7_75t_L g5105 ( 
.A(n_4655),
.B(n_4307),
.Y(n_5105)
);

NOR2xp67_ASAP7_75t_SL g5106 ( 
.A(n_4743),
.B(n_4307),
.Y(n_5106)
);

INVx2_ASAP7_75t_L g5107 ( 
.A(n_4576),
.Y(n_5107)
);

OAI21x1_ASAP7_75t_L g5108 ( 
.A1(n_4690),
.A2(n_4273),
.B(n_4112),
.Y(n_5108)
);

INVx3_ASAP7_75t_L g5109 ( 
.A(n_4645),
.Y(n_5109)
);

AOI21x1_ASAP7_75t_L g5110 ( 
.A1(n_4959),
.A2(n_4112),
.B(n_4102),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_4778),
.B(n_4492),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4780),
.Y(n_5112)
);

AOI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_4797),
.A2(n_4590),
.B(n_4589),
.Y(n_5113)
);

OAI21x1_ASAP7_75t_L g5114 ( 
.A1(n_4606),
.A2(n_4184),
.B(n_4112),
.Y(n_5114)
);

OAI21x1_ASAP7_75t_L g5115 ( 
.A1(n_4731),
.A2(n_4577),
.B(n_4848),
.Y(n_5115)
);

NAND2x1p5_ASAP7_75t_L g5116 ( 
.A(n_5018),
.B(n_4366),
.Y(n_5116)
);

INVx1_ASAP7_75t_SL g5117 ( 
.A(n_4883),
.Y(n_5117)
);

OA22x2_ASAP7_75t_L g5118 ( 
.A1(n_4855),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_5118)
);

OAI22xp5_ASAP7_75t_L g5119 ( 
.A1(n_4855),
.A2(n_4508),
.B1(n_4492),
.B2(n_4512),
.Y(n_5119)
);

NAND2xp5_ASAP7_75t_L g5120 ( 
.A(n_4840),
.B(n_4366),
.Y(n_5120)
);

HB1xp67_ASAP7_75t_L g5121 ( 
.A(n_4843),
.Y(n_5121)
);

AO21x1_ASAP7_75t_L g5122 ( 
.A1(n_4758),
.A2(n_373),
.B(n_374),
.Y(n_5122)
);

OAI21x1_ASAP7_75t_L g5123 ( 
.A1(n_4597),
.A2(n_4184),
.B(n_4392),
.Y(n_5123)
);

OAI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_4789),
.A2(n_374),
.B(n_375),
.Y(n_5124)
);

OAI21x1_ASAP7_75t_L g5125 ( 
.A1(n_4598),
.A2(n_4184),
.B(n_4392),
.Y(n_5125)
);

OAI21x1_ASAP7_75t_L g5126 ( 
.A1(n_4600),
.A2(n_4409),
.B(n_4401),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_4809),
.B(n_4401),
.Y(n_5127)
);

INVx2_ASAP7_75t_L g5128 ( 
.A(n_4593),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_4745),
.A2(n_4414),
.B(n_4409),
.Y(n_5129)
);

OAI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4633),
.A2(n_4414),
.B(n_4508),
.Y(n_5130)
);

OA21x2_ASAP7_75t_L g5131 ( 
.A1(n_4794),
.A2(n_4508),
.B(n_4512),
.Y(n_5131)
);

NOR2xp67_ASAP7_75t_L g5132 ( 
.A(n_4648),
.B(n_376),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_4823),
.B(n_376),
.Y(n_5133)
);

OAI21x1_ASAP7_75t_L g5134 ( 
.A1(n_4641),
.A2(n_4516),
.B(n_4512),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_4845),
.B(n_376),
.Y(n_5135)
);

NOR2xp33_ASAP7_75t_L g5136 ( 
.A(n_4925),
.B(n_377),
.Y(n_5136)
);

A2O1A1Ixp33_ASAP7_75t_L g5137 ( 
.A1(n_4650),
.A2(n_4516),
.B(n_380),
.C(n_378),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4918),
.Y(n_5138)
);

OAI22xp5_ASAP7_75t_L g5139 ( 
.A1(n_4580),
.A2(n_4516),
.B1(n_380),
.B2(n_378),
.Y(n_5139)
);

OAI22xp5_ASAP7_75t_L g5140 ( 
.A1(n_4750),
.A2(n_381),
.B1(n_378),
.B2(n_379),
.Y(n_5140)
);

OAI21x1_ASAP7_75t_L g5141 ( 
.A1(n_4933),
.A2(n_971),
.B(n_970),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_SL g5142 ( 
.A(n_4645),
.B(n_4768),
.Y(n_5142)
);

OR2x2_ASAP7_75t_L g5143 ( 
.A(n_4786),
.B(n_379),
.Y(n_5143)
);

NAND2x1p5_ASAP7_75t_L g5144 ( 
.A(n_4570),
.B(n_381),
.Y(n_5144)
);

OAI21x1_ASAP7_75t_L g5145 ( 
.A1(n_4610),
.A2(n_972),
.B(n_971),
.Y(n_5145)
);

OAI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4659),
.A2(n_382),
.B(n_383),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_4651),
.Y(n_5147)
);

AO31x2_ASAP7_75t_L g5148 ( 
.A1(n_4836),
.A2(n_384),
.A3(n_382),
.B(n_383),
.Y(n_5148)
);

INVx1_ASAP7_75t_L g5149 ( 
.A(n_4695),
.Y(n_5149)
);

INVx6_ASAP7_75t_L g5150 ( 
.A(n_5013),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_L g5151 ( 
.A(n_4957),
.B(n_382),
.Y(n_5151)
);

OAI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4749),
.A2(n_384),
.B(n_385),
.Y(n_5152)
);

HB1xp67_ASAP7_75t_L g5153 ( 
.A(n_4854),
.Y(n_5153)
);

OR2x6_ASAP7_75t_L g5154 ( 
.A(n_4801),
.B(n_384),
.Y(n_5154)
);

OAI21x1_ASAP7_75t_SL g5155 ( 
.A1(n_4885),
.A2(n_4756),
.B(n_4805),
.Y(n_5155)
);

BUFx3_ASAP7_75t_L g5156 ( 
.A(n_5013),
.Y(n_5156)
);

AND3x4_ASAP7_75t_L g5157 ( 
.A(n_4582),
.B(n_385),
.C(n_386),
.Y(n_5157)
);

OAI21x1_ASAP7_75t_L g5158 ( 
.A1(n_4674),
.A2(n_973),
.B(n_972),
.Y(n_5158)
);

AOI21xp5_ASAP7_75t_L g5159 ( 
.A1(n_4583),
.A2(n_386),
.B(n_387),
.Y(n_5159)
);

AOI21xp5_ASAP7_75t_L g5160 ( 
.A1(n_4581),
.A2(n_386),
.B(n_387),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_4961),
.B(n_388),
.Y(n_5161)
);

AOI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_4620),
.A2(n_388),
.B(n_389),
.Y(n_5162)
);

AND2x2_ASAP7_75t_L g5163 ( 
.A(n_4604),
.B(n_388),
.Y(n_5163)
);

OAI21x1_ASAP7_75t_L g5164 ( 
.A1(n_4679),
.A2(n_976),
.B(n_974),
.Y(n_5164)
);

OAI21x1_ASAP7_75t_L g5165 ( 
.A1(n_4699),
.A2(n_977),
.B(n_974),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_L g5166 ( 
.A(n_4965),
.B(n_389),
.Y(n_5166)
);

OAI21x1_ASAP7_75t_L g5167 ( 
.A1(n_4954),
.A2(n_979),
.B(n_978),
.Y(n_5167)
);

O2A1O1Ixp5_ASAP7_75t_L g5168 ( 
.A1(n_4714),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_5168)
);

AOI221xp5_ASAP7_75t_SL g5169 ( 
.A1(n_4994),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.C(n_393),
.Y(n_5169)
);

BUFx3_ASAP7_75t_L g5170 ( 
.A(n_4596),
.Y(n_5170)
);

AOI21xp33_ASAP7_75t_L g5171 ( 
.A1(n_4943),
.A2(n_390),
.B(n_391),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_5033),
.B(n_392),
.Y(n_5172)
);

AOI21x1_ASAP7_75t_L g5173 ( 
.A1(n_4622),
.A2(n_393),
.B(n_394),
.Y(n_5173)
);

AOI21x1_ASAP7_75t_L g5174 ( 
.A1(n_4978),
.A2(n_393),
.B(n_394),
.Y(n_5174)
);

AO21x1_ASAP7_75t_L g5175 ( 
.A1(n_4868),
.A2(n_394),
.B(n_395),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4971),
.B(n_395),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_L g5177 ( 
.A(n_4985),
.B(n_395),
.Y(n_5177)
);

INVx1_ASAP7_75t_SL g5178 ( 
.A(n_4804),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4993),
.Y(n_5179)
);

OAI21x1_ASAP7_75t_L g5180 ( 
.A1(n_4954),
.A2(n_980),
.B(n_979),
.Y(n_5180)
);

NOR2xp33_ASAP7_75t_L g5181 ( 
.A(n_4724),
.B(n_396),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_5011),
.B(n_396),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5022),
.Y(n_5183)
);

OAI21xp5_ASAP7_75t_L g5184 ( 
.A1(n_4777),
.A2(n_397),
.B(n_398),
.Y(n_5184)
);

AOI21xp5_ASAP7_75t_L g5185 ( 
.A1(n_4629),
.A2(n_397),
.B(n_398),
.Y(n_5185)
);

AND2x4_ASAP7_75t_L g5186 ( 
.A(n_4698),
.B(n_398),
.Y(n_5186)
);

OAI21x1_ASAP7_75t_L g5187 ( 
.A1(n_5017),
.A2(n_981),
.B(n_980),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_4826),
.B(n_399),
.Y(n_5188)
);

NAND2x1p5_ASAP7_75t_L g5189 ( 
.A(n_4747),
.B(n_399),
.Y(n_5189)
);

OAI21x1_ASAP7_75t_L g5190 ( 
.A1(n_5017),
.A2(n_984),
.B(n_981),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4865),
.Y(n_5191)
);

OAI21xp5_ASAP7_75t_L g5192 ( 
.A1(n_4632),
.A2(n_399),
.B(n_400),
.Y(n_5192)
);

AO22x1_ASAP7_75t_L g5193 ( 
.A1(n_4788),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_5193)
);

HB1xp67_ASAP7_75t_L g5194 ( 
.A(n_4832),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4605),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_SL g5196 ( 
.A(n_4768),
.B(n_400),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_4627),
.B(n_401),
.Y(n_5197)
);

OAI21x1_ASAP7_75t_L g5198 ( 
.A1(n_4723),
.A2(n_985),
.B(n_984),
.Y(n_5198)
);

OAI21x1_ASAP7_75t_SL g5199 ( 
.A1(n_4668),
.A2(n_401),
.B(n_402),
.Y(n_5199)
);

AOI21xp5_ASAP7_75t_L g5200 ( 
.A1(n_4700),
.A2(n_402),
.B(n_404),
.Y(n_5200)
);

OAI21x1_ASAP7_75t_SL g5201 ( 
.A1(n_4613),
.A2(n_404),
.B(n_405),
.Y(n_5201)
);

OAI21x1_ASAP7_75t_L g5202 ( 
.A1(n_4602),
.A2(n_988),
.B(n_987),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_4636),
.B(n_404),
.Y(n_5203)
);

INVx3_ASAP7_75t_L g5204 ( 
.A(n_4768),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_4642),
.B(n_405),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_4717),
.B(n_406),
.Y(n_5206)
);

BUFx6f_ASAP7_75t_L g5207 ( 
.A(n_4586),
.Y(n_5207)
);

INVxp67_ASAP7_75t_L g5208 ( 
.A(n_4698),
.Y(n_5208)
);

NAND2xp5_ASAP7_75t_L g5209 ( 
.A(n_4738),
.B(n_406),
.Y(n_5209)
);

OAI21x1_ASAP7_75t_L g5210 ( 
.A1(n_4686),
.A2(n_988),
.B(n_987),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_4585),
.A2(n_407),
.B(n_408),
.Y(n_5211)
);

OR2x2_ASAP7_75t_L g5212 ( 
.A(n_4671),
.B(n_408),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_SL g5213 ( 
.A(n_4698),
.B(n_408),
.Y(n_5213)
);

NAND2x1p5_ASAP7_75t_L g5214 ( 
.A(n_4648),
.B(n_409),
.Y(n_5214)
);

AOI21xp5_ASAP7_75t_L g5215 ( 
.A1(n_4572),
.A2(n_409),
.B(n_410),
.Y(n_5215)
);

HB1xp67_ASAP7_75t_L g5216 ( 
.A(n_4736),
.Y(n_5216)
);

INVx4_ASAP7_75t_L g5217 ( 
.A(n_4755),
.Y(n_5217)
);

INVx1_ASAP7_75t_SL g5218 ( 
.A(n_4846),
.Y(n_5218)
);

AOI21x1_ASAP7_75t_L g5219 ( 
.A1(n_4762),
.A2(n_5034),
.B(n_4891),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_L g5220 ( 
.A(n_4752),
.B(n_410),
.Y(n_5220)
);

INVx2_ASAP7_75t_SL g5221 ( 
.A(n_4586),
.Y(n_5221)
);

AOI21xp5_ASAP7_75t_L g5222 ( 
.A1(n_4950),
.A2(n_410),
.B(n_411),
.Y(n_5222)
);

AOI21xp33_ASAP7_75t_L g5223 ( 
.A1(n_4967),
.A2(n_411),
.B(n_412),
.Y(n_5223)
);

INVx2_ASAP7_75t_L g5224 ( 
.A(n_4753),
.Y(n_5224)
);

AOI22xp33_ASAP7_75t_L g5225 ( 
.A1(n_5027),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_5225)
);

BUFx12f_ASAP7_75t_L g5226 ( 
.A(n_4564),
.Y(n_5226)
);

CKINVDCx20_ASAP7_75t_R g5227 ( 
.A(n_4564),
.Y(n_5227)
);

AND2x2_ASAP7_75t_L g5228 ( 
.A(n_4621),
.B(n_413),
.Y(n_5228)
);

OAI21x1_ASAP7_75t_L g5229 ( 
.A1(n_4684),
.A2(n_991),
.B(n_990),
.Y(n_5229)
);

AOI21xp5_ASAP7_75t_L g5230 ( 
.A1(n_4595),
.A2(n_414),
.B(n_415),
.Y(n_5230)
);

BUFx2_ASAP7_75t_L g5231 ( 
.A(n_4711),
.Y(n_5231)
);

INVx5_ASAP7_75t_L g5232 ( 
.A(n_5027),
.Y(n_5232)
);

OAI21xp5_ASAP7_75t_L g5233 ( 
.A1(n_4722),
.A2(n_414),
.B(n_415),
.Y(n_5233)
);

OAI21x1_ASAP7_75t_L g5234 ( 
.A1(n_4675),
.A2(n_4710),
.B(n_4661),
.Y(n_5234)
);

OAI21xp5_ASAP7_75t_L g5235 ( 
.A1(n_4624),
.A2(n_414),
.B(n_415),
.Y(n_5235)
);

NAND2xp33_ASAP7_75t_L g5236 ( 
.A(n_5027),
.B(n_416),
.Y(n_5236)
);

OAI21x1_ASAP7_75t_L g5237 ( 
.A1(n_4675),
.A2(n_991),
.B(n_990),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_4783),
.Y(n_5238)
);

A2O1A1Ixp33_ASAP7_75t_L g5239 ( 
.A1(n_5001),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4811),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_4856),
.Y(n_5241)
);

AND2x4_ASAP7_75t_L g5242 ( 
.A(n_4711),
.B(n_417),
.Y(n_5242)
);

AOI21xp5_ASAP7_75t_L g5243 ( 
.A1(n_4796),
.A2(n_417),
.B(n_418),
.Y(n_5243)
);

BUFx12f_ASAP7_75t_L g5244 ( 
.A(n_4726),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_4910),
.Y(n_5245)
);

OAI22x1_ASAP7_75t_L g5246 ( 
.A1(n_4682),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_4915),
.Y(n_5247)
);

BUFx12f_ASAP7_75t_L g5248 ( 
.A(n_4920),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_4631),
.A2(n_419),
.B(n_420),
.Y(n_5249)
);

OAI21x1_ASAP7_75t_L g5250 ( 
.A1(n_4710),
.A2(n_994),
.B(n_993),
.Y(n_5250)
);

OAI21x1_ASAP7_75t_L g5251 ( 
.A1(n_4712),
.A2(n_994),
.B(n_993),
.Y(n_5251)
);

AOI21x1_ASAP7_75t_L g5252 ( 
.A1(n_4720),
.A2(n_421),
.B(n_422),
.Y(n_5252)
);

OR2x2_ASAP7_75t_L g5253 ( 
.A(n_4921),
.B(n_421),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_4941),
.B(n_422),
.Y(n_5254)
);

INVx1_ASAP7_75t_SL g5255 ( 
.A(n_4586),
.Y(n_5255)
);

BUFx6f_ASAP7_75t_L g5256 ( 
.A(n_4711),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_4730),
.A2(n_996),
.B(n_995),
.Y(n_5257)
);

AND2x4_ASAP7_75t_L g5258 ( 
.A(n_4828),
.B(n_422),
.Y(n_5258)
);

CKINVDCx5p33_ASAP7_75t_R g5259 ( 
.A(n_4772),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_4980),
.B(n_423),
.Y(n_5260)
);

AOI21xp5_ASAP7_75t_L g5261 ( 
.A1(n_4814),
.A2(n_424),
.B(n_425),
.Y(n_5261)
);

BUFx6f_ASAP7_75t_L g5262 ( 
.A(n_4896),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_L g5263 ( 
.A(n_4982),
.B(n_424),
.Y(n_5263)
);

AND2x4_ASAP7_75t_L g5264 ( 
.A(n_4795),
.B(n_4673),
.Y(n_5264)
);

NOR3xp33_ASAP7_75t_L g5265 ( 
.A(n_4882),
.B(n_424),
.C(n_425),
.Y(n_5265)
);

OAI21xp5_ASAP7_75t_L g5266 ( 
.A1(n_4694),
.A2(n_425),
.B(n_426),
.Y(n_5266)
);

AND3x4_ASAP7_75t_L g5267 ( 
.A(n_4969),
.B(n_426),
.C(n_427),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_4992),
.B(n_426),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_5006),
.B(n_427),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_5021),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_4817),
.B(n_428),
.Y(n_5271)
);

AOI21x1_ASAP7_75t_L g5272 ( 
.A1(n_4893),
.A2(n_428),
.B(n_429),
.Y(n_5272)
);

OAI21x1_ASAP7_75t_SL g5273 ( 
.A1(n_4896),
.A2(n_429),
.B(n_430),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_4822),
.B(n_429),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_4591),
.B(n_430),
.Y(n_5275)
);

OAI21x1_ASAP7_75t_L g5276 ( 
.A1(n_4886),
.A2(n_996),
.B(n_995),
.Y(n_5276)
);

NAND2x1p5_ASAP7_75t_L g5277 ( 
.A(n_4900),
.B(n_430),
.Y(n_5277)
);

BUFx12f_ASAP7_75t_L g5278 ( 
.A(n_4782),
.Y(n_5278)
);

OAI21x1_ASAP7_75t_L g5279 ( 
.A1(n_4819),
.A2(n_998),
.B(n_997),
.Y(n_5279)
);

OAI21xp5_ASAP7_75t_L g5280 ( 
.A1(n_4707),
.A2(n_431),
.B(n_433),
.Y(n_5280)
);

AOI21xp5_ASAP7_75t_L g5281 ( 
.A1(n_4693),
.A2(n_431),
.B(n_433),
.Y(n_5281)
);

AOI21xp5_ASAP7_75t_L g5282 ( 
.A1(n_4988),
.A2(n_434),
.B(n_435),
.Y(n_5282)
);

INVx6_ASAP7_75t_L g5283 ( 
.A(n_4900),
.Y(n_5283)
);

OAI21x1_ASAP7_75t_L g5284 ( 
.A1(n_4669),
.A2(n_1000),
.B(n_999),
.Y(n_5284)
);

INVxp67_ASAP7_75t_SL g5285 ( 
.A(n_4785),
.Y(n_5285)
);

AO31x2_ASAP7_75t_L g5286 ( 
.A1(n_4818),
.A2(n_438),
.A3(n_436),
.B(n_437),
.Y(n_5286)
);

OAI21x1_ASAP7_75t_L g5287 ( 
.A1(n_4644),
.A2(n_1000),
.B(n_999),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4936),
.A2(n_437),
.B(n_439),
.Y(n_5288)
);

NAND2x1_ASAP7_75t_L g5289 ( 
.A(n_5027),
.B(n_437),
.Y(n_5289)
);

NOR2x1_ASAP7_75t_SL g5290 ( 
.A(n_4603),
.B(n_439),
.Y(n_5290)
);

OAI22xp5_ASAP7_75t_L g5291 ( 
.A1(n_4609),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_5291)
);

NAND2xp5_ASAP7_75t_L g5292 ( 
.A(n_4880),
.B(n_440),
.Y(n_5292)
);

OAI22xp5_ASAP7_75t_L g5293 ( 
.A1(n_4601),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_5293)
);

AO31x2_ASAP7_75t_L g5294 ( 
.A1(n_4850),
.A2(n_444),
.A3(n_442),
.B(n_443),
.Y(n_5294)
);

NAND2x1p5_ASAP7_75t_L g5295 ( 
.A(n_4979),
.B(n_444),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4911),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_4630),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_4567),
.A2(n_444),
.B(n_445),
.Y(n_5298)
);

OAI21x1_ASAP7_75t_L g5299 ( 
.A1(n_4986),
.A2(n_1002),
.B(n_1001),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4575),
.A2(n_445),
.B(n_446),
.Y(n_5300)
);

OAI21x1_ASAP7_75t_L g5301 ( 
.A1(n_4670),
.A2(n_1003),
.B(n_1002),
.Y(n_5301)
);

A2O1A1Ixp33_ASAP7_75t_L g5302 ( 
.A1(n_4983),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_5302)
);

OAI21xp5_ASAP7_75t_L g5303 ( 
.A1(n_4654),
.A2(n_447),
.B(n_448),
.Y(n_5303)
);

INVx1_ASAP7_75t_SL g5304 ( 
.A(n_4678),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_4703),
.B(n_448),
.Y(n_5305)
);

OAI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_4667),
.A2(n_448),
.B(n_449),
.Y(n_5306)
);

OAI21x1_ASAP7_75t_L g5307 ( 
.A1(n_4757),
.A2(n_1005),
.B(n_1004),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_4821),
.B(n_449),
.Y(n_5308)
);

AOI21xp5_ASAP7_75t_L g5309 ( 
.A1(n_4578),
.A2(n_449),
.B(n_450),
.Y(n_5309)
);

INVx6_ASAP7_75t_L g5310 ( 
.A(n_4979),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_L g5311 ( 
.A(n_4769),
.B(n_450),
.Y(n_5311)
);

AND2x2_ASAP7_75t_L g5312 ( 
.A(n_4881),
.B(n_450),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_4776),
.B(n_451),
.Y(n_5313)
);

O2A1O1Ixp5_ASAP7_75t_L g5314 ( 
.A1(n_4614),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_5314)
);

OR2x2_ASAP7_75t_L g5315 ( 
.A(n_4949),
.B(n_452),
.Y(n_5315)
);

A2O1A1Ixp33_ASAP7_75t_L g5316 ( 
.A1(n_5030),
.A2(n_455),
.B(n_453),
.C(n_454),
.Y(n_5316)
);

A2O1A1Ixp33_ASAP7_75t_L g5317 ( 
.A1(n_4858),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_5317)
);

NAND2xp33_ASAP7_75t_L g5318 ( 
.A(n_4942),
.B(n_454),
.Y(n_5318)
);

OAI21xp5_ASAP7_75t_L g5319 ( 
.A1(n_4709),
.A2(n_455),
.B(n_456),
.Y(n_5319)
);

BUFx2_ASAP7_75t_L g5320 ( 
.A(n_5015),
.Y(n_5320)
);

A2O1A1Ixp33_ASAP7_75t_L g5321 ( 
.A1(n_5038),
.A2(n_458),
.B(n_456),
.C(n_457),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_4637),
.Y(n_5322)
);

OAI21x1_ASAP7_75t_SL g5323 ( 
.A1(n_4616),
.A2(n_457),
.B(n_458),
.Y(n_5323)
);

AOI21xp5_ASAP7_75t_L g5324 ( 
.A1(n_4955),
.A2(n_458),
.B(n_459),
.Y(n_5324)
);

AOI21xp5_ASAP7_75t_SL g5325 ( 
.A1(n_4930),
.A2(n_459),
.B(n_460),
.Y(n_5325)
);

NAND2x1p5_ASAP7_75t_L g5326 ( 
.A(n_4697),
.B(n_459),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_L g5327 ( 
.A(n_4608),
.B(n_4626),
.Y(n_5327)
);

OAI21x1_ASAP7_75t_SL g5328 ( 
.A1(n_4702),
.A2(n_460),
.B(n_461),
.Y(n_5328)
);

NOR2x1_ASAP7_75t_SL g5329 ( 
.A(n_4603),
.B(n_460),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_4951),
.B(n_461),
.Y(n_5330)
);

BUFx2_ASAP7_75t_L g5331 ( 
.A(n_4785),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_4587),
.B(n_4990),
.Y(n_5332)
);

AO31x2_ASAP7_75t_L g5333 ( 
.A1(n_4987),
.A2(n_4833),
.A3(n_4860),
.B(n_4932),
.Y(n_5333)
);

BUFx2_ASAP7_75t_L g5334 ( 
.A(n_4785),
.Y(n_5334)
);

AND2x4_ASAP7_75t_L g5335 ( 
.A(n_4887),
.B(n_461),
.Y(n_5335)
);

AOI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_4701),
.A2(n_462),
.B(n_463),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_4640),
.Y(n_5337)
);

OAI21x1_ASAP7_75t_L g5338 ( 
.A1(n_4989),
.A2(n_1007),
.B(n_1005),
.Y(n_5338)
);

AOI31xp33_ASAP7_75t_L g5339 ( 
.A1(n_4705),
.A2(n_464),
.A3(n_462),
.B(n_463),
.Y(n_5339)
);

NAND3xp33_ASAP7_75t_L g5340 ( 
.A(n_4940),
.B(n_462),
.C(n_463),
.Y(n_5340)
);

OAI21x1_ASAP7_75t_L g5341 ( 
.A1(n_4761),
.A2(n_4770),
.B(n_4729),
.Y(n_5341)
);

INVxp67_ASAP7_75t_SL g5342 ( 
.A(n_4806),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_4649),
.B(n_464),
.Y(n_5343)
);

AND2x2_ASAP7_75t_L g5344 ( 
.A(n_4968),
.B(n_464),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_4653),
.B(n_465),
.Y(n_5345)
);

AOI21x1_ASAP7_75t_L g5346 ( 
.A1(n_4803),
.A2(n_4766),
.B(n_4958),
.Y(n_5346)
);

AOI21xp33_ASAP7_75t_L g5347 ( 
.A1(n_4619),
.A2(n_465),
.B(n_466),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_4663),
.B(n_465),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_4775),
.Y(n_5349)
);

NAND2xp5_ASAP7_75t_L g5350 ( 
.A(n_4664),
.B(n_466),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4672),
.Y(n_5351)
);

AND2x4_ASAP7_75t_L g5352 ( 
.A(n_4890),
.B(n_467),
.Y(n_5352)
);

AOI21xp33_ASAP7_75t_L g5353 ( 
.A1(n_4839),
.A2(n_467),
.B(n_468),
.Y(n_5353)
);

AND2x4_ASAP7_75t_L g5354 ( 
.A(n_4806),
.B(n_468),
.Y(n_5354)
);

OAI21xp5_ASAP7_75t_L g5355 ( 
.A1(n_4960),
.A2(n_468),
.B(n_469),
.Y(n_5355)
);

INVx6_ASAP7_75t_SL g5356 ( 
.A(n_5054),
.Y(n_5356)
);

NAND2xp5_ASAP7_75t_L g5357 ( 
.A(n_5138),
.B(n_5147),
.Y(n_5357)
);

INVx4_ASAP7_75t_L g5358 ( 
.A(n_5150),
.Y(n_5358)
);

NAND2x1p5_ASAP7_75t_L g5359 ( 
.A(n_5156),
.B(n_5008),
.Y(n_5359)
);

BUFx2_ASAP7_75t_SL g5360 ( 
.A(n_5227),
.Y(n_5360)
);

BUFx3_ASAP7_75t_L g5361 ( 
.A(n_5150),
.Y(n_5361)
);

AOI22xp5_ASAP7_75t_L g5362 ( 
.A1(n_5236),
.A2(n_4975),
.B1(n_4919),
.B2(n_4974),
.Y(n_5362)
);

BUFx10_ASAP7_75t_L g5363 ( 
.A(n_5068),
.Y(n_5363)
);

INVx1_ASAP7_75t_SL g5364 ( 
.A(n_5091),
.Y(n_5364)
);

INVx3_ASAP7_75t_L g5365 ( 
.A(n_5061),
.Y(n_5365)
);

INVx2_ASAP7_75t_L g5366 ( 
.A(n_5049),
.Y(n_5366)
);

INVx3_ASAP7_75t_L g5367 ( 
.A(n_5226),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_5149),
.B(n_4825),
.Y(n_5368)
);

NAND2x1p5_ASAP7_75t_L g5369 ( 
.A(n_5106),
.B(n_5032),
.Y(n_5369)
);

NAND2xp5_ASAP7_75t_L g5370 ( 
.A(n_5216),
.B(n_4708),
.Y(n_5370)
);

INVx2_ASAP7_75t_L g5371 ( 
.A(n_5089),
.Y(n_5371)
);

BUFx3_ASAP7_75t_L g5372 ( 
.A(n_5067),
.Y(n_5372)
);

BUFx6f_ASAP7_75t_L g5373 ( 
.A(n_5262),
.Y(n_5373)
);

BUFx3_ASAP7_75t_L g5374 ( 
.A(n_5084),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_5053),
.Y(n_5375)
);

CKINVDCx8_ASAP7_75t_R g5376 ( 
.A(n_5259),
.Y(n_5376)
);

NAND2x1p5_ASAP7_75t_L g5377 ( 
.A(n_5170),
.B(n_5023),
.Y(n_5377)
);

BUFx3_ASAP7_75t_L g5378 ( 
.A(n_5264),
.Y(n_5378)
);

NAND2x1p5_ASAP7_75t_L g5379 ( 
.A(n_5117),
.B(n_4787),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_5056),
.Y(n_5380)
);

NAND2xp5_ASAP7_75t_L g5381 ( 
.A(n_5153),
.B(n_5297),
.Y(n_5381)
);

AND2x4_ASAP7_75t_L g5382 ( 
.A(n_5232),
.B(n_4806),
.Y(n_5382)
);

BUFx8_ASAP7_75t_L g5383 ( 
.A(n_5278),
.Y(n_5383)
);

NAND2x1p5_ASAP7_75t_L g5384 ( 
.A(n_5232),
.B(n_4813),
.Y(n_5384)
);

BUFx2_ASAP7_75t_L g5385 ( 
.A(n_5262),
.Y(n_5385)
);

INVx3_ASAP7_75t_L g5386 ( 
.A(n_5283),
.Y(n_5386)
);

INVx2_ASAP7_75t_L g5387 ( 
.A(n_5107),
.Y(n_5387)
);

INVx5_ASAP7_75t_L g5388 ( 
.A(n_5283),
.Y(n_5388)
);

INVx2_ASAP7_75t_SL g5389 ( 
.A(n_5304),
.Y(n_5389)
);

BUFx4f_ASAP7_75t_SL g5390 ( 
.A(n_5244),
.Y(n_5390)
);

NAND2x1p5_ASAP7_75t_L g5391 ( 
.A(n_5232),
.B(n_4947),
.Y(n_5391)
);

NOR2xp33_ASAP7_75t_SL g5392 ( 
.A(n_5157),
.B(n_4842),
.Y(n_5392)
);

INVx2_ASAP7_75t_L g5393 ( 
.A(n_5128),
.Y(n_5393)
);

BUFx12f_ASAP7_75t_L g5394 ( 
.A(n_5349),
.Y(n_5394)
);

AOI22xp33_ASAP7_75t_SL g5395 ( 
.A1(n_5057),
.A2(n_5026),
.B1(n_4867),
.B2(n_4869),
.Y(n_5395)
);

INVx3_ASAP7_75t_L g5396 ( 
.A(n_5310),
.Y(n_5396)
);

BUFx4f_ASAP7_75t_L g5397 ( 
.A(n_5267),
.Y(n_5397)
);

BUFx12f_ASAP7_75t_L g5398 ( 
.A(n_5217),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5071),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_5081),
.Y(n_5400)
);

BUFx8_ASAP7_75t_L g5401 ( 
.A(n_5248),
.Y(n_5401)
);

NAND2x1p5_ASAP7_75t_L g5402 ( 
.A(n_5289),
.B(n_4838),
.Y(n_5402)
);

BUFx6f_ASAP7_75t_L g5403 ( 
.A(n_5050),
.Y(n_5403)
);

INVx3_ASAP7_75t_SL g5404 ( 
.A(n_5178),
.Y(n_5404)
);

CKINVDCx11_ASAP7_75t_R g5405 ( 
.A(n_5218),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5083),
.Y(n_5406)
);

AOI22xp5_ASAP7_75t_L g5407 ( 
.A1(n_5318),
.A2(n_4657),
.B1(n_4872),
.B2(n_4841),
.Y(n_5407)
);

INVx2_ASAP7_75t_SL g5408 ( 
.A(n_5310),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5095),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5112),
.Y(n_5410)
);

NAND2x1p5_ASAP7_75t_L g5411 ( 
.A(n_5047),
.B(n_4660),
.Y(n_5411)
);

INVx3_ASAP7_75t_L g5412 ( 
.A(n_5050),
.Y(n_5412)
);

BUFx3_ASAP7_75t_L g5413 ( 
.A(n_5320),
.Y(n_5413)
);

INVx2_ASAP7_75t_L g5414 ( 
.A(n_5195),
.Y(n_5414)
);

CKINVDCx20_ASAP7_75t_R g5415 ( 
.A(n_5194),
.Y(n_5415)
);

BUFx8_ASAP7_75t_SL g5416 ( 
.A(n_5054),
.Y(n_5416)
);

BUFx12f_ASAP7_75t_L g5417 ( 
.A(n_5144),
.Y(n_5417)
);

BUFx5_ASAP7_75t_L g5418 ( 
.A(n_5354),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5179),
.Y(n_5419)
);

INVx1_ASAP7_75t_SL g5420 ( 
.A(n_5088),
.Y(n_5420)
);

HB1xp67_ASAP7_75t_L g5421 ( 
.A(n_5041),
.Y(n_5421)
);

BUFx6f_ASAP7_75t_L g5422 ( 
.A(n_5207),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5183),
.Y(n_5423)
);

INVx3_ASAP7_75t_L g5424 ( 
.A(n_5043),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5121),
.Y(n_5425)
);

HB1xp67_ASAP7_75t_L g5426 ( 
.A(n_5105),
.Y(n_5426)
);

AND2x2_ASAP7_75t_L g5427 ( 
.A(n_5094),
.B(n_4945),
.Y(n_5427)
);

INVx2_ASAP7_75t_L g5428 ( 
.A(n_5224),
.Y(n_5428)
);

CKINVDCx20_ASAP7_75t_R g5429 ( 
.A(n_5051),
.Y(n_5429)
);

INVx2_ASAP7_75t_SL g5430 ( 
.A(n_5207),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5322),
.B(n_4737),
.Y(n_5431)
);

NOR2xp33_ASAP7_75t_L g5432 ( 
.A(n_5136),
.B(n_5009),
.Y(n_5432)
);

INVx1_ASAP7_75t_SL g5433 ( 
.A(n_5090),
.Y(n_5433)
);

BUFx12f_ASAP7_75t_L g5434 ( 
.A(n_5214),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_5238),
.Y(n_5435)
);

INVx3_ASAP7_75t_L g5436 ( 
.A(n_5256),
.Y(n_5436)
);

INVx5_ASAP7_75t_L g5437 ( 
.A(n_5154),
.Y(n_5437)
);

INVx3_ASAP7_75t_L g5438 ( 
.A(n_5256),
.Y(n_5438)
);

NAND2x1p5_ASAP7_75t_L g5439 ( 
.A(n_5132),
.B(n_4798),
.Y(n_5439)
);

BUFx2_ASAP7_75t_L g5440 ( 
.A(n_5099),
.Y(n_5440)
);

HB1xp67_ASAP7_75t_L g5441 ( 
.A(n_5270),
.Y(n_5441)
);

INVx1_ASAP7_75t_SL g5442 ( 
.A(n_5255),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5069),
.Y(n_5443)
);

INVx1_ASAP7_75t_SL g5444 ( 
.A(n_5172),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_5240),
.Y(n_5445)
);

CKINVDCx20_ASAP7_75t_R g5446 ( 
.A(n_5163),
.Y(n_5446)
);

OR2x6_ASAP7_75t_L g5447 ( 
.A(n_5154),
.B(n_5103),
.Y(n_5447)
);

INVx3_ASAP7_75t_L g5448 ( 
.A(n_5109),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5073),
.Y(n_5449)
);

INVx3_ASAP7_75t_L g5450 ( 
.A(n_5204),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5120),
.B(n_4879),
.Y(n_5451)
);

CKINVDCx16_ASAP7_75t_R g5452 ( 
.A(n_5335),
.Y(n_5452)
);

INVx2_ASAP7_75t_SL g5453 ( 
.A(n_5231),
.Y(n_5453)
);

AOI22xp33_ASAP7_75t_L g5454 ( 
.A1(n_5265),
.A2(n_4830),
.B1(n_4718),
.B2(n_4628),
.Y(n_5454)
);

CKINVDCx16_ASAP7_75t_R g5455 ( 
.A(n_5352),
.Y(n_5455)
);

INVx6_ASAP7_75t_SL g5456 ( 
.A(n_5258),
.Y(n_5456)
);

INVx1_ASAP7_75t_SL g5457 ( 
.A(n_5142),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_5075),
.Y(n_5458)
);

BUFx6f_ASAP7_75t_SL g5459 ( 
.A(n_5186),
.Y(n_5459)
);

BUFx6f_ASAP7_75t_L g5460 ( 
.A(n_5116),
.Y(n_5460)
);

NAND2xp5_ASAP7_75t_L g5461 ( 
.A(n_5337),
.B(n_4793),
.Y(n_5461)
);

BUFx12f_ASAP7_75t_L g5462 ( 
.A(n_5189),
.Y(n_5462)
);

AND2x2_ASAP7_75t_L g5463 ( 
.A(n_5098),
.B(n_4903),
.Y(n_5463)
);

BUFx6f_ASAP7_75t_L g5464 ( 
.A(n_5221),
.Y(n_5464)
);

AND2x4_ASAP7_75t_L g5465 ( 
.A(n_5208),
.B(n_4922),
.Y(n_5465)
);

INVx3_ASAP7_75t_L g5466 ( 
.A(n_5277),
.Y(n_5466)
);

INVx3_ASAP7_75t_L g5467 ( 
.A(n_5295),
.Y(n_5467)
);

NOR2x1_ASAP7_75t_R g5468 ( 
.A(n_5228),
.B(n_4849),
.Y(n_5468)
);

NAND2x1p5_ASAP7_75t_L g5469 ( 
.A(n_5242),
.B(n_4922),
.Y(n_5469)
);

BUFx2_ASAP7_75t_L g5470 ( 
.A(n_5285),
.Y(n_5470)
);

AND2x4_ASAP7_75t_L g5471 ( 
.A(n_5342),
.B(n_4922),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5241),
.Y(n_5472)
);

NAND2x1p5_ASAP7_75t_L g5473 ( 
.A(n_5196),
.B(n_4929),
.Y(n_5473)
);

INVx1_ASAP7_75t_SL g5474 ( 
.A(n_5308),
.Y(n_5474)
);

OAI22xp33_ASAP7_75t_L g5475 ( 
.A1(n_5042),
.A2(n_4923),
.B1(n_4681),
.B2(n_4816),
.Y(n_5475)
);

INVx6_ASAP7_75t_SL g5476 ( 
.A(n_5101),
.Y(n_5476)
);

BUFx3_ASAP7_75t_L g5477 ( 
.A(n_5060),
.Y(n_5477)
);

BUFx3_ASAP7_75t_L g5478 ( 
.A(n_5127),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5245),
.Y(n_5479)
);

AND2x2_ASAP7_75t_L g5480 ( 
.A(n_5191),
.B(n_4976),
.Y(n_5480)
);

INVx5_ASAP7_75t_L g5481 ( 
.A(n_5331),
.Y(n_5481)
);

BUFx6f_ASAP7_75t_L g5482 ( 
.A(n_5334),
.Y(n_5482)
);

INVx4_ASAP7_75t_L g5483 ( 
.A(n_5118),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5247),
.Y(n_5484)
);

BUFx3_ASAP7_75t_L g5485 ( 
.A(n_5326),
.Y(n_5485)
);

BUFx5_ASAP7_75t_L g5486 ( 
.A(n_5351),
.Y(n_5486)
);

BUFx4_ASAP7_75t_SL g5487 ( 
.A(n_5143),
.Y(n_5487)
);

INVx3_ASAP7_75t_L g5488 ( 
.A(n_5093),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_5059),
.Y(n_5489)
);

AND2x2_ASAP7_75t_L g5490 ( 
.A(n_5296),
.B(n_4807),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_5104),
.Y(n_5491)
);

BUFx3_ASAP7_75t_L g5492 ( 
.A(n_5312),
.Y(n_5492)
);

NAND2x1p5_ASAP7_75t_L g5493 ( 
.A(n_5213),
.B(n_4929),
.Y(n_5493)
);

NAND2x1p5_ASAP7_75t_L g5494 ( 
.A(n_5167),
.B(n_4929),
.Y(n_5494)
);

INVx2_ASAP7_75t_SL g5495 ( 
.A(n_5086),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_5111),
.Y(n_5496)
);

INVx2_ASAP7_75t_L g5497 ( 
.A(n_5078),
.Y(n_5497)
);

INVx2_ASAP7_75t_SL g5498 ( 
.A(n_5087),
.Y(n_5498)
);

BUFx6f_ASAP7_75t_L g5499 ( 
.A(n_5126),
.Y(n_5499)
);

CKINVDCx5p33_ASAP7_75t_R g5500 ( 
.A(n_5344),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5064),
.B(n_4964),
.Y(n_5501)
);

BUFx3_ASAP7_75t_L g5502 ( 
.A(n_5181),
.Y(n_5502)
);

INVx3_ASAP7_75t_L g5503 ( 
.A(n_5253),
.Y(n_5503)
);

INVx2_ASAP7_75t_L g5504 ( 
.A(n_5092),
.Y(n_5504)
);

INVx1_ASAP7_75t_SL g5505 ( 
.A(n_5212),
.Y(n_5505)
);

BUFx6f_ASAP7_75t_L g5506 ( 
.A(n_5108),
.Y(n_5506)
);

BUFx4_ASAP7_75t_SL g5507 ( 
.A(n_5340),
.Y(n_5507)
);

NAND2x1p5_ASAP7_75t_L g5508 ( 
.A(n_5180),
.B(n_5020),
.Y(n_5508)
);

BUFx6f_ASAP7_75t_L g5509 ( 
.A(n_5123),
.Y(n_5509)
);

BUFx3_ASAP7_75t_L g5510 ( 
.A(n_5305),
.Y(n_5510)
);

INVx1_ASAP7_75t_SL g5511 ( 
.A(n_5311),
.Y(n_5511)
);

BUFx2_ASAP7_75t_SL g5512 ( 
.A(n_5175),
.Y(n_5512)
);

BUFx2_ASAP7_75t_SL g5513 ( 
.A(n_5122),
.Y(n_5513)
);

INVxp67_ASAP7_75t_SL g5514 ( 
.A(n_5131),
.Y(n_5514)
);

INVx4_ASAP7_75t_L g5515 ( 
.A(n_5315),
.Y(n_5515)
);

BUFx3_ASAP7_75t_L g5516 ( 
.A(n_5313),
.Y(n_5516)
);

CKINVDCx16_ASAP7_75t_R g5517 ( 
.A(n_5291),
.Y(n_5517)
);

AND2x2_ASAP7_75t_L g5518 ( 
.A(n_5332),
.B(n_4807),
.Y(n_5518)
);

BUFx6f_ASAP7_75t_L g5519 ( 
.A(n_5125),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5131),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5097),
.Y(n_5521)
);

INVx8_ASAP7_75t_L g5522 ( 
.A(n_5339),
.Y(n_5522)
);

CKINVDCx16_ASAP7_75t_R g5523 ( 
.A(n_5065),
.Y(n_5523)
);

BUFx12f_ASAP7_75t_L g5524 ( 
.A(n_5290),
.Y(n_5524)
);

INVx2_ASAP7_75t_SL g5525 ( 
.A(n_5246),
.Y(n_5525)
);

BUFx6f_ASAP7_75t_L g5526 ( 
.A(n_5114),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_5055),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_5327),
.B(n_4829),
.Y(n_5528)
);

INVx4_ASAP7_75t_L g5529 ( 
.A(n_5329),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_5151),
.Y(n_5530)
);

OAI22xp5_ASAP7_75t_L g5531 ( 
.A1(n_5052),
.A2(n_4952),
.B1(n_4931),
.B2(n_4999),
.Y(n_5531)
);

INVx6_ASAP7_75t_SL g5532 ( 
.A(n_5070),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5161),
.Y(n_5533)
);

NAND2x1p5_ASAP7_75t_L g5534 ( 
.A(n_5187),
.B(n_5020),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5166),
.Y(n_5535)
);

BUFx3_ASAP7_75t_L g5536 ( 
.A(n_5292),
.Y(n_5536)
);

INVx5_ASAP7_75t_L g5537 ( 
.A(n_5193),
.Y(n_5537)
);

INVxp67_ASAP7_75t_SL g5538 ( 
.A(n_5110),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_5048),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_L g5540 ( 
.A(n_5080),
.B(n_4831),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5176),
.Y(n_5541)
);

BUFx6f_ASAP7_75t_SL g5542 ( 
.A(n_5273),
.Y(n_5542)
);

NAND2xp5_ASAP7_75t_L g5543 ( 
.A(n_5275),
.B(n_4834),
.Y(n_5543)
);

BUFx12f_ASAP7_75t_L g5544 ( 
.A(n_5225),
.Y(n_5544)
);

AOI22xp33_ASAP7_75t_L g5545 ( 
.A1(n_5544),
.A2(n_5155),
.B1(n_5140),
.B2(n_5215),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5375),
.Y(n_5546)
);

BUFx6f_ASAP7_75t_L g5547 ( 
.A(n_5373),
.Y(n_5547)
);

A2O1A1Ixp33_ASAP7_75t_L g5548 ( 
.A1(n_5522),
.A2(n_5085),
.B(n_5082),
.C(n_5243),
.Y(n_5548)
);

INVx3_ASAP7_75t_L g5549 ( 
.A(n_5358),
.Y(n_5549)
);

OR2x6_ASAP7_75t_L g5550 ( 
.A(n_5447),
.B(n_5119),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5380),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5399),
.Y(n_5552)
);

INVx3_ASAP7_75t_L g5553 ( 
.A(n_5374),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5400),
.Y(n_5554)
);

AO32x2_ASAP7_75t_L g5555 ( 
.A1(n_5389),
.A2(n_5063),
.A3(n_5139),
.B1(n_5293),
.B2(n_4837),
.Y(n_5555)
);

OAI21x1_ASAP7_75t_L g5556 ( 
.A1(n_5488),
.A2(n_5066),
.B(n_5076),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5406),
.Y(n_5557)
);

INVxp67_ASAP7_75t_L g5558 ( 
.A(n_5468),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5409),
.Y(n_5559)
);

NOR2xp33_ASAP7_75t_L g5560 ( 
.A(n_5404),
.B(n_5330),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5410),
.Y(n_5561)
);

NAND2xp5_ASAP7_75t_L g5562 ( 
.A(n_5518),
.B(n_5115),
.Y(n_5562)
);

INVx6_ASAP7_75t_L g5563 ( 
.A(n_5363),
.Y(n_5563)
);

NAND2xp5_ASAP7_75t_L g5564 ( 
.A(n_5443),
.B(n_5521),
.Y(n_5564)
);

O2A1O1Ixp33_ASAP7_75t_SL g5565 ( 
.A1(n_5525),
.A2(n_5079),
.B(n_5137),
.C(n_5096),
.Y(n_5565)
);

OAI21x1_ASAP7_75t_L g5566 ( 
.A1(n_5538),
.A2(n_5113),
.B(n_5134),
.Y(n_5566)
);

OAI21x1_ASAP7_75t_L g5567 ( 
.A1(n_5520),
.A2(n_5384),
.B(n_5514),
.Y(n_5567)
);

AND2x4_ASAP7_75t_L g5568 ( 
.A(n_5470),
.B(n_5234),
.Y(n_5568)
);

AO21x2_ASAP7_75t_L g5569 ( 
.A1(n_5527),
.A2(n_5381),
.B(n_5539),
.Y(n_5569)
);

OAI21xp5_ASAP7_75t_L g5570 ( 
.A1(n_5397),
.A2(n_5168),
.B(n_5169),
.Y(n_5570)
);

AOI22xp33_ASAP7_75t_L g5571 ( 
.A1(n_5483),
.A2(n_5347),
.B1(n_5199),
.B2(n_5328),
.Y(n_5571)
);

OAI222xp33_ASAP7_75t_L g5572 ( 
.A1(n_5447),
.A2(n_5040),
.B1(n_5272),
.B2(n_5219),
.C1(n_5230),
.C2(n_5288),
.Y(n_5572)
);

OAI22xp5_ASAP7_75t_L g5573 ( 
.A1(n_5523),
.A2(n_5517),
.B1(n_5437),
.B2(n_5522),
.Y(n_5573)
);

NOR2xp33_ASAP7_75t_L g5574 ( 
.A(n_5360),
.B(n_5271),
.Y(n_5574)
);

AOI22xp33_ASAP7_75t_L g5575 ( 
.A1(n_5512),
.A2(n_5353),
.B1(n_5223),
.B2(n_5266),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_5490),
.B(n_5148),
.Y(n_5576)
);

BUFx3_ASAP7_75t_L g5577 ( 
.A(n_5372),
.Y(n_5577)
);

OAI21x1_ASAP7_75t_L g5578 ( 
.A1(n_5402),
.A2(n_5130),
.B(n_5062),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_L g5579 ( 
.A(n_5489),
.B(n_5148),
.Y(n_5579)
);

OAI21x1_ASAP7_75t_L g5580 ( 
.A1(n_5365),
.A2(n_5044),
.B(n_5058),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5419),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5441),
.Y(n_5582)
);

NAND2xp5_ASAP7_75t_L g5583 ( 
.A(n_5449),
.B(n_5074),
.Y(n_5583)
);

OAI21x1_ASAP7_75t_L g5584 ( 
.A1(n_5386),
.A2(n_5046),
.B(n_5173),
.Y(n_5584)
);

BUFx2_ASAP7_75t_L g5585 ( 
.A(n_5415),
.Y(n_5585)
);

INVx2_ASAP7_75t_L g5586 ( 
.A(n_5486),
.Y(n_5586)
);

OAI21x1_ASAP7_75t_L g5587 ( 
.A1(n_5396),
.A2(n_5174),
.B(n_5102),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_L g5588 ( 
.A(n_5458),
.B(n_5133),
.Y(n_5588)
);

AOI22xp33_ASAP7_75t_SL g5589 ( 
.A1(n_5513),
.A2(n_5201),
.B1(n_5355),
.B2(n_5323),
.Y(n_5589)
);

INVx2_ASAP7_75t_L g5590 ( 
.A(n_5486),
.Y(n_5590)
);

INVxp67_ASAP7_75t_L g5591 ( 
.A(n_5492),
.Y(n_5591)
);

OA21x2_ASAP7_75t_L g5592 ( 
.A1(n_5540),
.A2(n_5129),
.B(n_5039),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5425),
.B(n_5421),
.Y(n_5593)
);

AOI22xp5_ASAP7_75t_L g5594 ( 
.A1(n_5362),
.A2(n_5407),
.B1(n_5542),
.B2(n_5529),
.Y(n_5594)
);

INVxp33_ASAP7_75t_L g5595 ( 
.A(n_5405),
.Y(n_5595)
);

OAI21x1_ASAP7_75t_L g5596 ( 
.A1(n_5439),
.A2(n_5346),
.B(n_5252),
.Y(n_5596)
);

INVx3_ASAP7_75t_L g5597 ( 
.A(n_5361),
.Y(n_5597)
);

OAI21xp5_ASAP7_75t_L g5598 ( 
.A1(n_5392),
.A2(n_5211),
.B(n_5160),
.Y(n_5598)
);

BUFx2_ASAP7_75t_SL g5599 ( 
.A(n_5388),
.Y(n_5599)
);

AOI21xp5_ASAP7_75t_L g5600 ( 
.A1(n_5408),
.A2(n_5072),
.B(n_5325),
.Y(n_5600)
);

AO21x2_ASAP7_75t_L g5601 ( 
.A1(n_5370),
.A2(n_5171),
.B(n_5324),
.Y(n_5601)
);

OAI22xp5_ASAP7_75t_L g5602 ( 
.A1(n_5437),
.A2(n_5100),
.B1(n_5302),
.B2(n_5239),
.Y(n_5602)
);

OAI21x1_ASAP7_75t_L g5603 ( 
.A1(n_5411),
.A2(n_5391),
.B(n_5494),
.Y(n_5603)
);

AOI221xp5_ASAP7_75t_L g5604 ( 
.A1(n_5530),
.A2(n_5309),
.B1(n_5300),
.B2(n_5298),
.C(n_5343),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5423),
.Y(n_5605)
);

OAI21x1_ASAP7_75t_L g5606 ( 
.A1(n_5508),
.A2(n_5190),
.B(n_5338),
.Y(n_5606)
);

OAI21xp33_ASAP7_75t_SL g5607 ( 
.A1(n_5420),
.A2(n_5250),
.B(n_5237),
.Y(n_5607)
);

O2A1O1Ixp33_ASAP7_75t_SL g5608 ( 
.A1(n_5364),
.A2(n_5316),
.B(n_5321),
.C(n_5317),
.Y(n_5608)
);

OAI21x1_ASAP7_75t_L g5609 ( 
.A1(n_5534),
.A2(n_5202),
.B(n_5165),
.Y(n_5609)
);

INVx2_ASAP7_75t_L g5610 ( 
.A(n_5486),
.Y(n_5610)
);

INVx2_ASAP7_75t_L g5611 ( 
.A(n_5366),
.Y(n_5611)
);

INVx2_ASAP7_75t_SL g5612 ( 
.A(n_5378),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_L g5613 ( 
.A(n_5533),
.B(n_5135),
.Y(n_5613)
);

BUFx3_ASAP7_75t_L g5614 ( 
.A(n_5383),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5445),
.Y(n_5615)
);

INVx2_ASAP7_75t_L g5616 ( 
.A(n_5371),
.Y(n_5616)
);

AOI21xp5_ASAP7_75t_L g5617 ( 
.A1(n_5385),
.A2(n_5280),
.B(n_5249),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_5426),
.B(n_5045),
.Y(n_5618)
);

INVx3_ASAP7_75t_L g5619 ( 
.A(n_5416),
.Y(n_5619)
);

AND2x2_ASAP7_75t_L g5620 ( 
.A(n_5463),
.B(n_5045),
.Y(n_5620)
);

INVx2_ASAP7_75t_L g5621 ( 
.A(n_5387),
.Y(n_5621)
);

AOI22xp33_ASAP7_75t_L g5622 ( 
.A1(n_5537),
.A2(n_5319),
.B1(n_5306),
.B2(n_5303),
.Y(n_5622)
);

NAND3xp33_ASAP7_75t_L g5623 ( 
.A(n_5537),
.B(n_5395),
.C(n_5535),
.Y(n_5623)
);

OAI21xp5_ASAP7_75t_L g5624 ( 
.A1(n_5432),
.A2(n_5314),
.B(n_5159),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_5357),
.Y(n_5625)
);

AND2x2_ASAP7_75t_L g5626 ( 
.A(n_5424),
.B(n_5077),
.Y(n_5626)
);

OAI222xp33_ASAP7_75t_L g5627 ( 
.A1(n_5452),
.A2(n_5274),
.B1(n_5005),
.B2(n_4812),
.C1(n_4800),
.C2(n_5336),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_5541),
.B(n_4767),
.Y(n_5628)
);

INVx1_ASAP7_75t_SL g5629 ( 
.A(n_5413),
.Y(n_5629)
);

BUFx3_ASAP7_75t_L g5630 ( 
.A(n_5401),
.Y(n_5630)
);

OA21x2_ASAP7_75t_L g5631 ( 
.A1(n_5440),
.A2(n_5182),
.B(n_5177),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_5393),
.Y(n_5632)
);

OAI21x1_ASAP7_75t_L g5633 ( 
.A1(n_5379),
.A2(n_5210),
.B(n_5145),
.Y(n_5633)
);

AO21x2_ASAP7_75t_L g5634 ( 
.A1(n_5461),
.A2(n_5203),
.B(n_5197),
.Y(n_5634)
);

NOR2xp33_ASAP7_75t_L g5635 ( 
.A(n_5398),
.B(n_5345),
.Y(n_5635)
);

OAI21x1_ASAP7_75t_L g5636 ( 
.A1(n_5359),
.A2(n_5141),
.B(n_5341),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5472),
.Y(n_5637)
);

CKINVDCx5p33_ASAP7_75t_R g5638 ( 
.A(n_5376),
.Y(n_5638)
);

INVx2_ASAP7_75t_L g5639 ( 
.A(n_5414),
.Y(n_5639)
);

INVx2_ASAP7_75t_L g5640 ( 
.A(n_5428),
.Y(n_5640)
);

OAI21x1_ASAP7_75t_L g5641 ( 
.A1(n_5369),
.A2(n_5164),
.B(n_5158),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5479),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_5484),
.Y(n_5643)
);

OAI22xp5_ASAP7_75t_L g5644 ( 
.A1(n_5455),
.A2(n_5206),
.B1(n_5209),
.B2(n_5205),
.Y(n_5644)
);

AO31x2_ASAP7_75t_L g5645 ( 
.A1(n_5501),
.A2(n_5220),
.A3(n_5260),
.B(n_5254),
.Y(n_5645)
);

OAI21x1_ASAP7_75t_L g5646 ( 
.A1(n_5473),
.A2(n_5493),
.B(n_5448),
.Y(n_5646)
);

OA21x2_ASAP7_75t_L g5647 ( 
.A1(n_5435),
.A2(n_5268),
.B(n_5263),
.Y(n_5647)
);

NAND2xp5_ASAP7_75t_L g5648 ( 
.A(n_5497),
.B(n_5188),
.Y(n_5648)
);

AND2x4_ASAP7_75t_L g5649 ( 
.A(n_5388),
.B(n_5035),
.Y(n_5649)
);

OAI21x1_ASAP7_75t_L g5650 ( 
.A1(n_5450),
.A2(n_5279),
.B(n_5269),
.Y(n_5650)
);

OAI21x1_ASAP7_75t_L g5651 ( 
.A1(n_5466),
.A2(n_5301),
.B(n_5287),
.Y(n_5651)
);

BUFx12f_ASAP7_75t_L g5652 ( 
.A(n_5462),
.Y(n_5652)
);

AO21x2_ASAP7_75t_L g5653 ( 
.A1(n_5431),
.A2(n_4646),
.B(n_5152),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5504),
.Y(n_5654)
);

NOR2xp33_ASAP7_75t_L g5655 ( 
.A(n_5367),
.B(n_5348),
.Y(n_5655)
);

INVx2_ASAP7_75t_L g5656 ( 
.A(n_5491),
.Y(n_5656)
);

OAI21x1_ASAP7_75t_L g5657 ( 
.A1(n_5467),
.A2(n_5229),
.B(n_5257),
.Y(n_5657)
);

OAI21x1_ASAP7_75t_L g5658 ( 
.A1(n_5412),
.A2(n_5276),
.B(n_5198),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5496),
.Y(n_5659)
);

BUFx8_ASAP7_75t_L g5660 ( 
.A(n_5394),
.Y(n_5660)
);

NAND2xp5_ASAP7_75t_L g5661 ( 
.A(n_5495),
.B(n_5350),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5498),
.Y(n_5662)
);

OAI21xp5_ASAP7_75t_L g5663 ( 
.A1(n_5454),
.A2(n_5146),
.B(n_5124),
.Y(n_5663)
);

NAND2xp5_ASAP7_75t_L g5664 ( 
.A(n_5480),
.B(n_5286),
.Y(n_5664)
);

AND2x4_ASAP7_75t_L g5665 ( 
.A(n_5478),
.B(n_5020),
.Y(n_5665)
);

NAND2xp5_ASAP7_75t_SL g5666 ( 
.A(n_5373),
.B(n_5235),
.Y(n_5666)
);

OAI21xp33_ASAP7_75t_SL g5667 ( 
.A1(n_5474),
.A2(n_5192),
.B(n_5184),
.Y(n_5667)
);

BUFx6f_ASAP7_75t_L g5668 ( 
.A(n_5403),
.Y(n_5668)
);

BUFx3_ASAP7_75t_L g5669 ( 
.A(n_5390),
.Y(n_5669)
);

AO32x2_ASAP7_75t_L g5670 ( 
.A1(n_5453),
.A2(n_5004),
.A3(n_4917),
.B1(n_4884),
.B2(n_4981),
.Y(n_5670)
);

AND2x2_ASAP7_75t_L g5671 ( 
.A(n_5427),
.B(n_4569),
.Y(n_5671)
);

BUFx3_ASAP7_75t_L g5672 ( 
.A(n_5417),
.Y(n_5672)
);

INVx3_ASAP7_75t_L g5673 ( 
.A(n_5524),
.Y(n_5673)
);

OAI21x1_ASAP7_75t_L g5674 ( 
.A1(n_5436),
.A2(n_5284),
.B(n_5185),
.Y(n_5674)
);

NAND2x1p5_ASAP7_75t_L g5675 ( 
.A(n_5485),
.B(n_5460),
.Y(n_5675)
);

OAI22xp5_ASAP7_75t_L g5676 ( 
.A1(n_5446),
.A2(n_5233),
.B1(n_4912),
.B2(n_4859),
.Y(n_5676)
);

AOI22xp33_ASAP7_75t_SL g5677 ( 
.A1(n_5573),
.A2(n_5459),
.B1(n_5477),
.B2(n_5434),
.Y(n_5677)
);

BUFx6f_ASAP7_75t_L g5678 ( 
.A(n_5614),
.Y(n_5678)
);

OA21x2_ASAP7_75t_L g5679 ( 
.A1(n_5567),
.A2(n_5368),
.B(n_5528),
.Y(n_5679)
);

BUFx2_ASAP7_75t_L g5680 ( 
.A(n_5577),
.Y(n_5680)
);

INVxp67_ASAP7_75t_L g5681 ( 
.A(n_5585),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5582),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5615),
.Y(n_5683)
);

OAI21x1_ASAP7_75t_L g5684 ( 
.A1(n_5556),
.A2(n_5377),
.B(n_5438),
.Y(n_5684)
);

NAND2x1p5_ASAP7_75t_L g5685 ( 
.A(n_5672),
.B(n_5673),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5546),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5551),
.Y(n_5687)
);

AOI22xp33_ASAP7_75t_L g5688 ( 
.A1(n_5570),
.A2(n_5502),
.B1(n_5532),
.B2(n_5515),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_5552),
.Y(n_5689)
);

AOI22xp33_ASAP7_75t_L g5690 ( 
.A1(n_5663),
.A2(n_5510),
.B1(n_5516),
.B2(n_5536),
.Y(n_5690)
);

AOI22xp33_ASAP7_75t_L g5691 ( 
.A1(n_5623),
.A2(n_5531),
.B1(n_5475),
.B2(n_5511),
.Y(n_5691)
);

OAI21x1_ASAP7_75t_L g5692 ( 
.A1(n_5580),
.A2(n_5503),
.B(n_5469),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_5611),
.Y(n_5693)
);

INVxp67_ASAP7_75t_L g5694 ( 
.A(n_5585),
.Y(n_5694)
);

CKINVDCx5p33_ASAP7_75t_R g5695 ( 
.A(n_5630),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_5554),
.Y(n_5696)
);

INVx4_ASAP7_75t_L g5697 ( 
.A(n_5652),
.Y(n_5697)
);

BUFx2_ASAP7_75t_R g5698 ( 
.A(n_5669),
.Y(n_5698)
);

AND2x2_ASAP7_75t_L g5699 ( 
.A(n_5626),
.B(n_5433),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5620),
.B(n_5618),
.Y(n_5700)
);

NAND2xp5_ASAP7_75t_L g5701 ( 
.A(n_5576),
.B(n_5442),
.Y(n_5701)
);

INVx1_ASAP7_75t_SL g5702 ( 
.A(n_5629),
.Y(n_5702)
);

INVx3_ASAP7_75t_L g5703 ( 
.A(n_5563),
.Y(n_5703)
);

INVxp67_ASAP7_75t_L g5704 ( 
.A(n_5560),
.Y(n_5704)
);

HB1xp67_ASAP7_75t_L g5705 ( 
.A(n_5612),
.Y(n_5705)
);

AOI21x1_ASAP7_75t_L g5706 ( 
.A1(n_5550),
.A2(n_5543),
.B(n_5382),
.Y(n_5706)
);

CKINVDCx11_ASAP7_75t_R g5707 ( 
.A(n_5547),
.Y(n_5707)
);

OAI21x1_ASAP7_75t_L g5708 ( 
.A1(n_5566),
.A2(n_5578),
.B(n_5603),
.Y(n_5708)
);

CKINVDCx11_ASAP7_75t_R g5709 ( 
.A(n_5547),
.Y(n_5709)
);

INVx2_ASAP7_75t_L g5710 ( 
.A(n_5616),
.Y(n_5710)
);

AOI22xp5_ASAP7_75t_L g5711 ( 
.A1(n_5667),
.A2(n_5505),
.B1(n_5444),
.B2(n_5500),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5621),
.Y(n_5712)
);

AOI22xp33_ASAP7_75t_SL g5713 ( 
.A1(n_5599),
.A2(n_5429),
.B1(n_5418),
.B2(n_5481),
.Y(n_5713)
);

NAND2xp5_ASAP7_75t_L g5714 ( 
.A(n_5664),
.B(n_5482),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_5557),
.Y(n_5715)
);

NAND2x1p5_ASAP7_75t_L g5716 ( 
.A(n_5549),
.B(n_5460),
.Y(n_5716)
);

OA21x2_ASAP7_75t_L g5717 ( 
.A1(n_5562),
.A2(n_5451),
.B(n_5457),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5559),
.Y(n_5718)
);

CKINVDCx11_ASAP7_75t_R g5719 ( 
.A(n_5660),
.Y(n_5719)
);

HB1xp67_ASAP7_75t_L g5720 ( 
.A(n_5553),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5561),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_5581),
.Y(n_5722)
);

OA21x2_ASAP7_75t_L g5723 ( 
.A1(n_5583),
.A2(n_5471),
.B(n_5465),
.Y(n_5723)
);

NOR2xp33_ASAP7_75t_L g5724 ( 
.A(n_5595),
.B(n_5356),
.Y(n_5724)
);

OAI21xp33_ASAP7_75t_SL g5725 ( 
.A1(n_5550),
.A2(n_5476),
.B(n_5430),
.Y(n_5725)
);

OAI21x1_ASAP7_75t_L g5726 ( 
.A1(n_5646),
.A2(n_5200),
.B(n_5162),
.Y(n_5726)
);

INVx2_ASAP7_75t_L g5727 ( 
.A(n_5632),
.Y(n_5727)
);

BUFx10_ASAP7_75t_L g5728 ( 
.A(n_5563),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5605),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_5637),
.Y(n_5730)
);

INVx3_ASAP7_75t_L g5731 ( 
.A(n_5619),
.Y(n_5731)
);

AND2x2_ASAP7_75t_L g5732 ( 
.A(n_5662),
.B(n_5482),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5642),
.Y(n_5733)
);

HB1xp67_ASAP7_75t_L g5734 ( 
.A(n_5656),
.Y(n_5734)
);

BUFx2_ASAP7_75t_L g5735 ( 
.A(n_5597),
.Y(n_5735)
);

INVx1_ASAP7_75t_SL g5736 ( 
.A(n_5599),
.Y(n_5736)
);

INVx3_ASAP7_75t_L g5737 ( 
.A(n_5675),
.Y(n_5737)
);

AND2x4_ASAP7_75t_L g5738 ( 
.A(n_5568),
.B(n_5481),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5643),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5654),
.Y(n_5740)
);

BUFx2_ASAP7_75t_R g5741 ( 
.A(n_5638),
.Y(n_5741)
);

HB1xp67_ASAP7_75t_L g5742 ( 
.A(n_5659),
.Y(n_5742)
);

OAI21x1_ASAP7_75t_L g5743 ( 
.A1(n_5584),
.A2(n_5261),
.B(n_5251),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5564),
.Y(n_5744)
);

INVx3_ASAP7_75t_L g5745 ( 
.A(n_5668),
.Y(n_5745)
);

BUFx2_ASAP7_75t_L g5746 ( 
.A(n_5591),
.Y(n_5746)
);

INVx8_ASAP7_75t_L g5747 ( 
.A(n_5668),
.Y(n_5747)
);

INVx3_ASAP7_75t_L g5748 ( 
.A(n_5665),
.Y(n_5748)
);

INVx2_ASAP7_75t_SL g5749 ( 
.A(n_5671),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5625),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5639),
.Y(n_5751)
);

INVx2_ASAP7_75t_L g5752 ( 
.A(n_5640),
.Y(n_5752)
);

OAI21x1_ASAP7_75t_L g5753 ( 
.A1(n_5579),
.A2(n_5307),
.B(n_4815),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5647),
.Y(n_5754)
);

INVx2_ASAP7_75t_L g5755 ( 
.A(n_5647),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_5593),
.Y(n_5756)
);

BUFx3_ASAP7_75t_L g5757 ( 
.A(n_5635),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_5574),
.Y(n_5758)
);

INVx2_ASAP7_75t_L g5759 ( 
.A(n_5568),
.Y(n_5759)
);

AND2x2_ASAP7_75t_L g5760 ( 
.A(n_5594),
.B(n_5569),
.Y(n_5760)
);

BUFx2_ASAP7_75t_L g5761 ( 
.A(n_5607),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5631),
.Y(n_5762)
);

BUFx3_ASAP7_75t_L g5763 ( 
.A(n_5655),
.Y(n_5763)
);

BUFx6f_ASAP7_75t_L g5764 ( 
.A(n_5649),
.Y(n_5764)
);

AOI21x1_ASAP7_75t_L g5765 ( 
.A1(n_5596),
.A2(n_4677),
.B(n_4676),
.Y(n_5765)
);

INVx2_ASAP7_75t_SL g5766 ( 
.A(n_5661),
.Y(n_5766)
);

BUFx2_ASAP7_75t_L g5767 ( 
.A(n_5558),
.Y(n_5767)
);

INVx3_ASAP7_75t_L g5768 ( 
.A(n_5649),
.Y(n_5768)
);

NAND2x1p5_ASAP7_75t_L g5769 ( 
.A(n_5666),
.B(n_5403),
.Y(n_5769)
);

BUFx6f_ASAP7_75t_L g5770 ( 
.A(n_5651),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5628),
.Y(n_5771)
);

AND2x4_ASAP7_75t_L g5772 ( 
.A(n_5586),
.B(n_5590),
.Y(n_5772)
);

HB1xp67_ASAP7_75t_L g5773 ( 
.A(n_5631),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5588),
.Y(n_5774)
);

AOI22xp33_ASAP7_75t_L g5775 ( 
.A1(n_5598),
.A2(n_5602),
.B1(n_5545),
.B2(n_5622),
.Y(n_5775)
);

CKINVDCx11_ASAP7_75t_R g5776 ( 
.A(n_5644),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5648),
.Y(n_5777)
);

BUFx3_ASAP7_75t_L g5778 ( 
.A(n_5613),
.Y(n_5778)
);

OAI21xp5_ASAP7_75t_L g5779 ( 
.A1(n_5548),
.A2(n_4991),
.B(n_4835),
.Y(n_5779)
);

HB1xp67_ASAP7_75t_L g5780 ( 
.A(n_5634),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_5645),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5645),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5592),
.Y(n_5783)
);

AOI22xp33_ASAP7_75t_SL g5784 ( 
.A1(n_5676),
.A2(n_5600),
.B1(n_5601),
.B2(n_5617),
.Y(n_5784)
);

AOI22xp33_ASAP7_75t_L g5785 ( 
.A1(n_5653),
.A2(n_5418),
.B1(n_5456),
.B2(n_4592),
.Y(n_5785)
);

AOI22xp33_ASAP7_75t_L g5786 ( 
.A1(n_5589),
.A2(n_5418),
.B1(n_4779),
.B2(n_4808),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5592),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5636),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_5610),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5650),
.Y(n_5790)
);

AO21x2_ASAP7_75t_L g5791 ( 
.A1(n_5565),
.A2(n_4692),
.B(n_4691),
.Y(n_5791)
);

AND2x4_ASAP7_75t_L g5792 ( 
.A(n_5657),
.B(n_5464),
.Y(n_5792)
);

NAND2xp5_ASAP7_75t_L g5793 ( 
.A(n_5575),
.B(n_5464),
.Y(n_5793)
);

BUFx3_ASAP7_75t_L g5794 ( 
.A(n_5587),
.Y(n_5794)
);

CKINVDCx11_ASAP7_75t_R g5795 ( 
.A(n_5624),
.Y(n_5795)
);

HB1xp67_ASAP7_75t_L g5796 ( 
.A(n_5633),
.Y(n_5796)
);

AO21x2_ASAP7_75t_L g5797 ( 
.A1(n_5572),
.A2(n_4715),
.B(n_4706),
.Y(n_5797)
);

INVx6_ASAP7_75t_L g5798 ( 
.A(n_5555),
.Y(n_5798)
);

INVx8_ASAP7_75t_L g5799 ( 
.A(n_5555),
.Y(n_5799)
);

AND2x2_ASAP7_75t_L g5800 ( 
.A(n_5670),
.B(n_5506),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5606),
.Y(n_5801)
);

INVx2_ASAP7_75t_L g5802 ( 
.A(n_5658),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5609),
.Y(n_5803)
);

INVx4_ASAP7_75t_L g5804 ( 
.A(n_5670),
.Y(n_5804)
);

CKINVDCx11_ASAP7_75t_R g5805 ( 
.A(n_5627),
.Y(n_5805)
);

OA21x2_ASAP7_75t_L g5806 ( 
.A1(n_5641),
.A2(n_4725),
.B(n_4716),
.Y(n_5806)
);

BUFx3_ASAP7_75t_L g5807 ( 
.A(n_5719),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5683),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5680),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5680),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5740),
.Y(n_5811)
);

INVx3_ASAP7_75t_L g5812 ( 
.A(n_5685),
.Y(n_5812)
);

OR2x6_ASAP7_75t_L g5813 ( 
.A(n_5747),
.B(n_5674),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_5734),
.Y(n_5814)
);

INVx3_ASAP7_75t_L g5815 ( 
.A(n_5728),
.Y(n_5815)
);

AND2x6_ASAP7_75t_L g5816 ( 
.A(n_5736),
.B(n_5506),
.Y(n_5816)
);

AND2x4_ASAP7_75t_L g5817 ( 
.A(n_5735),
.B(n_5422),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5750),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5742),
.Y(n_5819)
);

BUFx2_ASAP7_75t_L g5820 ( 
.A(n_5725),
.Y(n_5820)
);

OA21x2_ASAP7_75t_L g5821 ( 
.A1(n_5761),
.A2(n_5571),
.B(n_5604),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5686),
.Y(n_5822)
);

HB1xp67_ASAP7_75t_L g5823 ( 
.A(n_5735),
.Y(n_5823)
);

AOI22xp33_ASAP7_75t_L g5824 ( 
.A1(n_5805),
.A2(n_5799),
.B1(n_5795),
.B2(n_5798),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5687),
.Y(n_5825)
);

OAI21x1_ASAP7_75t_L g5826 ( 
.A1(n_5706),
.A2(n_5037),
.B(n_5036),
.Y(n_5826)
);

INVx2_ASAP7_75t_L g5827 ( 
.A(n_5746),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5689),
.Y(n_5828)
);

INVx2_ASAP7_75t_L g5829 ( 
.A(n_5746),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5696),
.Y(n_5830)
);

INVx2_ASAP7_75t_L g5831 ( 
.A(n_5754),
.Y(n_5831)
);

O2A1O1Ixp33_ASAP7_75t_L g5832 ( 
.A1(n_5775),
.A2(n_5608),
.B(n_4966),
.C(n_4889),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5755),
.Y(n_5833)
);

INVx3_ASAP7_75t_L g5834 ( 
.A(n_5678),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5715),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5718),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5721),
.Y(n_5837)
);

INVx2_ASAP7_75t_L g5838 ( 
.A(n_5693),
.Y(n_5838)
);

OAI21x1_ASAP7_75t_L g5839 ( 
.A1(n_5706),
.A2(n_4852),
.B(n_4844),
.Y(n_5839)
);

HB1xp67_ASAP7_75t_L g5840 ( 
.A(n_5705),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5722),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_5729),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5730),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5733),
.Y(n_5844)
);

OAI21x1_ASAP7_75t_L g5845 ( 
.A1(n_5717),
.A2(n_5762),
.B(n_5768),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5710),
.Y(n_5846)
);

INVx2_ASAP7_75t_L g5847 ( 
.A(n_5712),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5739),
.Y(n_5848)
);

OAI21x1_ASAP7_75t_L g5849 ( 
.A1(n_5717),
.A2(n_4623),
.B(n_5299),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5727),
.Y(n_5850)
);

OR2x2_ASAP7_75t_L g5851 ( 
.A(n_5771),
.B(n_5499),
.Y(n_5851)
);

AOI22xp33_ASAP7_75t_L g5852 ( 
.A1(n_5799),
.A2(n_5499),
.B1(n_5519),
.B2(n_5509),
.Y(n_5852)
);

INVx2_ASAP7_75t_L g5853 ( 
.A(n_5751),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5744),
.Y(n_5854)
);

CKINVDCx5p33_ASAP7_75t_R g5855 ( 
.A(n_5695),
.Y(n_5855)
);

INVx2_ASAP7_75t_L g5856 ( 
.A(n_5752),
.Y(n_5856)
);

BUFx6f_ASAP7_75t_L g5857 ( 
.A(n_5678),
.Y(n_5857)
);

BUFx12f_ASAP7_75t_L g5858 ( 
.A(n_5697),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5773),
.Y(n_5859)
);

INVx3_ASAP7_75t_L g5860 ( 
.A(n_5731),
.Y(n_5860)
);

O2A1O1Ixp33_ASAP7_75t_L g5861 ( 
.A1(n_5767),
.A2(n_4897),
.B(n_4861),
.C(n_4878),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5781),
.Y(n_5862)
);

INVx3_ASAP7_75t_L g5863 ( 
.A(n_5707),
.Y(n_5863)
);

HB1xp67_ASAP7_75t_L g5864 ( 
.A(n_5681),
.Y(n_5864)
);

AND2x4_ASAP7_75t_L g5865 ( 
.A(n_5703),
.B(n_5422),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5782),
.Y(n_5866)
);

AOI22xp33_ASAP7_75t_L g5867 ( 
.A1(n_5798),
.A2(n_5509),
.B1(n_5519),
.B2(n_5526),
.Y(n_5867)
);

BUFx6f_ASAP7_75t_L g5868 ( 
.A(n_5709),
.Y(n_5868)
);

BUFx2_ASAP7_75t_L g5869 ( 
.A(n_5767),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5682),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5701),
.Y(n_5871)
);

BUFx6f_ASAP7_75t_L g5872 ( 
.A(n_5747),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5777),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5756),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5780),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5789),
.Y(n_5876)
);

OR2x2_ASAP7_75t_L g5877 ( 
.A(n_5774),
.B(n_5526),
.Y(n_5877)
);

INVxp67_ASAP7_75t_L g5878 ( 
.A(n_5720),
.Y(n_5878)
);

BUFx6f_ASAP7_75t_L g5879 ( 
.A(n_5716),
.Y(n_5879)
);

INVxp67_ASAP7_75t_L g5880 ( 
.A(n_5698),
.Y(n_5880)
);

INVx2_ASAP7_75t_L g5881 ( 
.A(n_5749),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5803),
.Y(n_5882)
);

INVx2_ASAP7_75t_L g5883 ( 
.A(n_5802),
.Y(n_5883)
);

AND2x2_ASAP7_75t_L g5884 ( 
.A(n_5700),
.B(n_5286),
.Y(n_5884)
);

AND2x2_ASAP7_75t_L g5885 ( 
.A(n_5723),
.B(n_5487),
.Y(n_5885)
);

OAI21xp5_ASAP7_75t_L g5886 ( 
.A1(n_5784),
.A2(n_4963),
.B(n_4962),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5694),
.Y(n_5887)
);

BUFx2_ASAP7_75t_SL g5888 ( 
.A(n_5737),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_5796),
.Y(n_5889)
);

NOR3xp33_ASAP7_75t_L g5890 ( 
.A(n_5804),
.B(n_4901),
.C(n_4875),
.Y(n_5890)
);

HB1xp67_ASAP7_75t_L g5891 ( 
.A(n_5702),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5714),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5793),
.Y(n_5893)
);

AO22x1_ASAP7_75t_L g5894 ( 
.A1(n_5761),
.A2(n_5507),
.B1(n_4866),
.B2(n_4732),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5766),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5788),
.Y(n_5896)
);

INVx2_ASAP7_75t_L g5897 ( 
.A(n_5801),
.Y(n_5897)
);

CKINVDCx6p67_ASAP7_75t_R g5898 ( 
.A(n_5776),
.Y(n_5898)
);

BUFx3_ASAP7_75t_L g5899 ( 
.A(n_5757),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5783),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5679),
.Y(n_5901)
);

AND2x4_ASAP7_75t_L g5902 ( 
.A(n_5724),
.B(n_4728),
.Y(n_5902)
);

OR2x6_ASAP7_75t_L g5903 ( 
.A(n_5769),
.B(n_4938),
.Y(n_5903)
);

OR2x2_ASAP7_75t_L g5904 ( 
.A(n_5778),
.B(n_4997),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_5787),
.Y(n_5905)
);

AND2x6_ASAP7_75t_L g5906 ( 
.A(n_5711),
.B(n_5016),
.Y(n_5906)
);

BUFx2_ASAP7_75t_L g5907 ( 
.A(n_5723),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5790),
.Y(n_5908)
);

BUFx2_ASAP7_75t_L g5909 ( 
.A(n_5679),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5699),
.Y(n_5910)
);

AND2x4_ASAP7_75t_L g5911 ( 
.A(n_5758),
.B(n_4734),
.Y(n_5911)
);

AOI22xp33_ASAP7_75t_L g5912 ( 
.A1(n_5797),
.A2(n_4799),
.B1(n_4820),
.B2(n_5281),
.Y(n_5912)
);

NAND2xp5_ASAP7_75t_L g5913 ( 
.A(n_5800),
.B(n_5333),
.Y(n_5913)
);

BUFx2_ASAP7_75t_L g5914 ( 
.A(n_5738),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5772),
.Y(n_5915)
);

OA21x2_ASAP7_75t_L g5916 ( 
.A1(n_5684),
.A2(n_4744),
.B(n_4735),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5794),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5772),
.Y(n_5918)
);

INVx2_ASAP7_75t_L g5919 ( 
.A(n_5759),
.Y(n_5919)
);

OA21x2_ASAP7_75t_L g5920 ( 
.A1(n_5760),
.A2(n_4748),
.B(n_4746),
.Y(n_5920)
);

NAND2xp5_ASAP7_75t_L g5921 ( 
.A(n_5869),
.B(n_5691),
.Y(n_5921)
);

NAND2xp5_ASAP7_75t_L g5922 ( 
.A(n_5869),
.B(n_5785),
.Y(n_5922)
);

OR2x6_ASAP7_75t_L g5923 ( 
.A(n_5888),
.B(n_5726),
.Y(n_5923)
);

HB1xp67_ASAP7_75t_L g5924 ( 
.A(n_5840),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5900),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5864),
.Y(n_5926)
);

INVx2_ASAP7_75t_L g5927 ( 
.A(n_5899),
.Y(n_5927)
);

AO21x2_ASAP7_75t_L g5928 ( 
.A1(n_5875),
.A2(n_5708),
.B(n_5765),
.Y(n_5928)
);

OR2x2_ASAP7_75t_L g5929 ( 
.A(n_5827),
.B(n_5806),
.Y(n_5929)
);

OAI21x1_ASAP7_75t_L g5930 ( 
.A1(n_5845),
.A2(n_5692),
.B(n_5690),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5905),
.Y(n_5931)
);

BUFx2_ASAP7_75t_L g5932 ( 
.A(n_5885),
.Y(n_5932)
);

BUFx2_ASAP7_75t_L g5933 ( 
.A(n_5907),
.Y(n_5933)
);

OR2x2_ASAP7_75t_L g5934 ( 
.A(n_5829),
.B(n_5806),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5891),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5887),
.Y(n_5936)
);

INVx1_ASAP7_75t_L g5937 ( 
.A(n_5809),
.Y(n_5937)
);

AO21x2_ASAP7_75t_L g5938 ( 
.A1(n_5889),
.A2(n_5765),
.B(n_5791),
.Y(n_5938)
);

INVx1_ASAP7_75t_L g5939 ( 
.A(n_5810),
.Y(n_5939)
);

OR2x2_ASAP7_75t_L g5940 ( 
.A(n_5814),
.B(n_5764),
.Y(n_5940)
);

INVx2_ASAP7_75t_L g5941 ( 
.A(n_5819),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5873),
.Y(n_5942)
);

INVx2_ASAP7_75t_L g5943 ( 
.A(n_5823),
.Y(n_5943)
);

INVx2_ASAP7_75t_L g5944 ( 
.A(n_5831),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5854),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5833),
.Y(n_5946)
);

HB1xp67_ASAP7_75t_L g5947 ( 
.A(n_5859),
.Y(n_5947)
);

OR2x6_ASAP7_75t_L g5948 ( 
.A(n_5888),
.B(n_5764),
.Y(n_5948)
);

INVx2_ASAP7_75t_L g5949 ( 
.A(n_5907),
.Y(n_5949)
);

NOR2x1_ASAP7_75t_L g5950 ( 
.A(n_5820),
.B(n_5763),
.Y(n_5950)
);

OAI21xp5_ASAP7_75t_L g5951 ( 
.A1(n_5821),
.A2(n_5677),
.B(n_5688),
.Y(n_5951)
);

NAND2xp5_ASAP7_75t_L g5952 ( 
.A(n_5920),
.B(n_5704),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5818),
.Y(n_5953)
);

AND2x2_ASAP7_75t_L g5954 ( 
.A(n_5914),
.B(n_5738),
.Y(n_5954)
);

OR2x6_ASAP7_75t_L g5955 ( 
.A(n_5858),
.B(n_5807),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5838),
.Y(n_5956)
);

OA21x2_ASAP7_75t_L g5957 ( 
.A1(n_5824),
.A2(n_5743),
.B(n_5792),
.Y(n_5957)
);

NAND2xp5_ASAP7_75t_L g5958 ( 
.A(n_5920),
.B(n_5753),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5846),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5874),
.Y(n_5960)
);

INVx3_ASAP7_75t_L g5961 ( 
.A(n_5812),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5808),
.Y(n_5962)
);

AOI22xp33_ASAP7_75t_L g5963 ( 
.A1(n_5906),
.A2(n_5779),
.B1(n_5786),
.B2(n_5770),
.Y(n_5963)
);

AOI221xp5_ASAP7_75t_L g5964 ( 
.A1(n_5894),
.A2(n_5770),
.B1(n_4727),
.B2(n_4658),
.C(n_4972),
.Y(n_5964)
);

INVx2_ASAP7_75t_L g5965 ( 
.A(n_5847),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5811),
.Y(n_5966)
);

INVx3_ASAP7_75t_SL g5967 ( 
.A(n_5868),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5822),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5825),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5828),
.Y(n_5970)
);

HB1xp67_ASAP7_75t_L g5971 ( 
.A(n_5878),
.Y(n_5971)
);

AND2x2_ASAP7_75t_L g5972 ( 
.A(n_5914),
.B(n_5732),
.Y(n_5972)
);

INVx2_ASAP7_75t_L g5973 ( 
.A(n_5850),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5853),
.Y(n_5974)
);

OR2x2_ASAP7_75t_L g5975 ( 
.A(n_5913),
.B(n_5748),
.Y(n_5975)
);

BUFx2_ASAP7_75t_L g5976 ( 
.A(n_5898),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5830),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5835),
.Y(n_5978)
);

INVx2_ASAP7_75t_L g5979 ( 
.A(n_5856),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5836),
.Y(n_5980)
);

INVx2_ASAP7_75t_L g5981 ( 
.A(n_5870),
.Y(n_5981)
);

AND2x2_ASAP7_75t_L g5982 ( 
.A(n_5893),
.B(n_5713),
.Y(n_5982)
);

AOI21xp5_ASAP7_75t_L g5983 ( 
.A1(n_5820),
.A2(n_5745),
.B(n_4895),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5837),
.Y(n_5984)
);

INVx3_ASAP7_75t_L g5985 ( 
.A(n_5857),
.Y(n_5985)
);

OR2x2_ASAP7_75t_L g5986 ( 
.A(n_5884),
.B(n_4760),
.Y(n_5986)
);

OAI21xp5_ASAP7_75t_L g5987 ( 
.A1(n_5821),
.A2(n_4946),
.B(n_5282),
.Y(n_5987)
);

OR2x2_ASAP7_75t_L g5988 ( 
.A(n_5871),
.B(n_4763),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5841),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5842),
.Y(n_5990)
);

AND2x4_ASAP7_75t_L g5991 ( 
.A(n_5815),
.B(n_5003),
.Y(n_5991)
);

INVx3_ASAP7_75t_L g5992 ( 
.A(n_5857),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5843),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5844),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5848),
.Y(n_5995)
);

HB1xp67_ASAP7_75t_L g5996 ( 
.A(n_5882),
.Y(n_5996)
);

AND2x2_ASAP7_75t_L g5997 ( 
.A(n_5860),
.B(n_5741),
.Y(n_5997)
);

INVx2_ASAP7_75t_L g5998 ( 
.A(n_5876),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5896),
.Y(n_5999)
);

BUFx3_ASAP7_75t_L g6000 ( 
.A(n_5868),
.Y(n_6000)
);

INVx3_ASAP7_75t_L g6001 ( 
.A(n_5863),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5879),
.B(n_5817),
.Y(n_6002)
);

AOI21xp5_ASAP7_75t_L g6003 ( 
.A1(n_5880),
.A2(n_4874),
.B(n_4863),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5910),
.Y(n_6004)
);

AO21x2_ASAP7_75t_L g6005 ( 
.A1(n_5917),
.A2(n_4781),
.B(n_4765),
.Y(n_6005)
);

AO21x2_ASAP7_75t_L g6006 ( 
.A1(n_5901),
.A2(n_4791),
.B(n_4790),
.Y(n_6006)
);

AO21x2_ASAP7_75t_L g6007 ( 
.A1(n_5862),
.A2(n_4864),
.B(n_4851),
.Y(n_6007)
);

AND2x4_ASAP7_75t_L g6008 ( 
.A(n_5834),
.B(n_5014),
.Y(n_6008)
);

INVx2_ASAP7_75t_L g6009 ( 
.A(n_5897),
.Y(n_6009)
);

INVx2_ASAP7_75t_L g6010 ( 
.A(n_5883),
.Y(n_6010)
);

AND2x2_ASAP7_75t_L g6011 ( 
.A(n_5879),
.B(n_5294),
.Y(n_6011)
);

AND2x2_ASAP7_75t_L g6012 ( 
.A(n_5852),
.B(n_5294),
.Y(n_6012)
);

INVx2_ASAP7_75t_L g6013 ( 
.A(n_5919),
.Y(n_6013)
);

HB1xp67_ASAP7_75t_L g6014 ( 
.A(n_5908),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5867),
.B(n_5333),
.Y(n_6015)
);

OR2x2_ASAP7_75t_L g6016 ( 
.A(n_5877),
.B(n_5024),
.Y(n_6016)
);

BUFx2_ASAP7_75t_L g6017 ( 
.A(n_5813),
.Y(n_6017)
);

AO21x2_ASAP7_75t_L g6018 ( 
.A1(n_5866),
.A2(n_4871),
.B(n_4870),
.Y(n_6018)
);

NAND2xp5_ASAP7_75t_L g6019 ( 
.A(n_5906),
.B(n_4877),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5851),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5892),
.Y(n_6021)
);

AOI221xp5_ASAP7_75t_L g6022 ( 
.A1(n_5832),
.A2(n_4773),
.B1(n_4953),
.B2(n_5222),
.C(n_4742),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5895),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_5906),
.B(n_4899),
.Y(n_6024)
);

INVx2_ASAP7_75t_L g6025 ( 
.A(n_5881),
.Y(n_6025)
);

INVx2_ASAP7_75t_L g6026 ( 
.A(n_5915),
.Y(n_6026)
);

NAND2xp5_ASAP7_75t_L g6027 ( 
.A(n_5890),
.B(n_4902),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5904),
.Y(n_6028)
);

OR2x2_ASAP7_75t_L g6029 ( 
.A(n_5909),
.B(n_4904),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5909),
.Y(n_6030)
);

HB1xp67_ASAP7_75t_L g6031 ( 
.A(n_5916),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5918),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5916),
.Y(n_6033)
);

INVx2_ASAP7_75t_L g6034 ( 
.A(n_5849),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5911),
.Y(n_6035)
);

BUFx2_ASAP7_75t_L g6036 ( 
.A(n_5813),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5903),
.Y(n_6037)
);

NAND2xp5_ASAP7_75t_L g6038 ( 
.A(n_5912),
.B(n_4905),
.Y(n_6038)
);

BUFx3_ASAP7_75t_L g6039 ( 
.A(n_5855),
.Y(n_6039)
);

AND2x4_ASAP7_75t_L g6040 ( 
.A(n_5872),
.B(n_4927),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5865),
.B(n_4934),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5903),
.Y(n_6042)
);

BUFx6f_ASAP7_75t_L g6043 ( 
.A(n_5872),
.Y(n_6043)
);

AND2x2_ASAP7_75t_L g6044 ( 
.A(n_5902),
.B(n_4935),
.Y(n_6044)
);

OA21x2_ASAP7_75t_L g6045 ( 
.A1(n_5826),
.A2(n_5839),
.B(n_5886),
.Y(n_6045)
);

NAND2xp5_ASAP7_75t_L g6046 ( 
.A(n_5816),
.B(n_4937),
.Y(n_6046)
);

INVx2_ASAP7_75t_L g6047 ( 
.A(n_5816),
.Y(n_6047)
);

INVx1_ASAP7_75t_L g6048 ( 
.A(n_5816),
.Y(n_6048)
);

INVx1_ASAP7_75t_L g6049 ( 
.A(n_5861),
.Y(n_6049)
);

AO21x2_ASAP7_75t_L g6050 ( 
.A1(n_5875),
.A2(n_4909),
.B(n_4906),
.Y(n_6050)
);

INVx2_ASAP7_75t_L g6051 ( 
.A(n_5899),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5864),
.Y(n_6052)
);

BUFx3_ASAP7_75t_L g6053 ( 
.A(n_5807),
.Y(n_6053)
);

INVx2_ASAP7_75t_L g6054 ( 
.A(n_5899),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5864),
.Y(n_6055)
);

INVx2_ASAP7_75t_L g6056 ( 
.A(n_5899),
.Y(n_6056)
);

HB1xp67_ASAP7_75t_L g6057 ( 
.A(n_5840),
.Y(n_6057)
);

NAND2xp33_ASAP7_75t_SL g6058 ( 
.A(n_5820),
.B(n_4928),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_5900),
.Y(n_6059)
);

INVx3_ASAP7_75t_L g6060 ( 
.A(n_5899),
.Y(n_6060)
);

AOI21xp5_ASAP7_75t_L g6061 ( 
.A1(n_5885),
.A2(n_4874),
.B(n_4639),
.Y(n_6061)
);

OAI21x1_ASAP7_75t_L g6062 ( 
.A1(n_5845),
.A2(n_4913),
.B(n_4898),
.Y(n_6062)
);

AND2x4_ASAP7_75t_L g6063 ( 
.A(n_5885),
.B(n_4612),
.Y(n_6063)
);

AND2x2_ASAP7_75t_L g6064 ( 
.A(n_5885),
.B(n_4916),
.Y(n_6064)
);

INVx2_ASAP7_75t_L g6065 ( 
.A(n_5899),
.Y(n_6065)
);

AND2x2_ASAP7_75t_L g6066 ( 
.A(n_5885),
.B(n_4892),
.Y(n_6066)
);

OA21x2_ASAP7_75t_L g6067 ( 
.A1(n_5824),
.A2(n_4634),
.B(n_4784),
.Y(n_6067)
);

INVxp67_ASAP7_75t_SL g6068 ( 
.A(n_6060),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_5924),
.Y(n_6069)
);

AND2x2_ASAP7_75t_L g6070 ( 
.A(n_5932),
.B(n_4894),
.Y(n_6070)
);

NOR2xp33_ASAP7_75t_L g6071 ( 
.A(n_5976),
.B(n_469),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5933),
.Y(n_6072)
);

INVxp67_ASAP7_75t_L g6073 ( 
.A(n_5976),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5933),
.Y(n_6074)
);

INVxp67_ASAP7_75t_SL g6075 ( 
.A(n_6053),
.Y(n_6075)
);

OR2x2_ASAP7_75t_L g6076 ( 
.A(n_5935),
.B(n_470),
.Y(n_6076)
);

INVx2_ASAP7_75t_L g6077 ( 
.A(n_5927),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_6057),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5971),
.Y(n_6079)
);

NAND2xp5_ASAP7_75t_L g6080 ( 
.A(n_6028),
.B(n_4995),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_6030),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_5932),
.B(n_4996),
.Y(n_6082)
);

INVx2_ASAP7_75t_L g6083 ( 
.A(n_6051),
.Y(n_6083)
);

AOI221xp5_ASAP7_75t_L g6084 ( 
.A1(n_6049),
.A2(n_5007),
.B1(n_5002),
.B2(n_4998),
.C(n_4771),
.Y(n_6084)
);

INVx2_ASAP7_75t_SL g6085 ( 
.A(n_5948),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5948),
.B(n_4688),
.Y(n_6086)
);

OAI221xp5_ASAP7_75t_L g6087 ( 
.A1(n_5951),
.A2(n_5028),
.B1(n_4984),
.B2(n_5029),
.C(n_5025),
.Y(n_6087)
);

INVxp67_ASAP7_75t_L g6088 ( 
.A(n_6054),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5947),
.Y(n_6089)
);

BUFx2_ASAP7_75t_L g6090 ( 
.A(n_5997),
.Y(n_6090)
);

AND2x2_ASAP7_75t_L g6091 ( 
.A(n_5961),
.B(n_4689),
.Y(n_6091)
);

NAND2xp5_ASAP7_75t_L g6092 ( 
.A(n_5926),
.B(n_4696),
.Y(n_6092)
);

AND2x2_ASAP7_75t_L g6093 ( 
.A(n_5954),
.B(n_5031),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_6052),
.Y(n_6094)
);

INVx2_ASAP7_75t_L g6095 ( 
.A(n_6056),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_L g6096 ( 
.A(n_6055),
.B(n_6050),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5949),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5943),
.Y(n_6098)
);

OR2x2_ASAP7_75t_SL g6099 ( 
.A(n_5957),
.B(n_4639),
.Y(n_6099)
);

NAND2x1p5_ASAP7_75t_L g6100 ( 
.A(n_6001),
.B(n_4656),
.Y(n_6100)
);

NAND2xp5_ASAP7_75t_L g6101 ( 
.A(n_6021),
.B(n_4652),
.Y(n_6101)
);

INVx2_ASAP7_75t_L g6102 ( 
.A(n_6065),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_6002),
.B(n_470),
.Y(n_6103)
);

INVx3_ASAP7_75t_L g6104 ( 
.A(n_6043),
.Y(n_6104)
);

NAND2xp5_ASAP7_75t_L g6105 ( 
.A(n_6005),
.B(n_5010),
.Y(n_6105)
);

INVx2_ASAP7_75t_L g6106 ( 
.A(n_6025),
.Y(n_6106)
);

OR2x2_ASAP7_75t_L g6107 ( 
.A(n_5952),
.B(n_470),
.Y(n_6107)
);

INVx2_ASAP7_75t_L g6108 ( 
.A(n_5944),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5996),
.Y(n_6109)
);

INVxp67_ASAP7_75t_L g6110 ( 
.A(n_6000),
.Y(n_6110)
);

AO31x2_ASAP7_75t_L g6111 ( 
.A1(n_6017),
.A2(n_6036),
.A3(n_5921),
.B(n_5922),
.Y(n_6111)
);

HB1xp67_ASAP7_75t_L g6112 ( 
.A(n_5937),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5936),
.Y(n_6113)
);

AND2x2_ASAP7_75t_L g6114 ( 
.A(n_5972),
.B(n_5982),
.Y(n_6114)
);

HB1xp67_ASAP7_75t_L g6115 ( 
.A(n_5939),
.Y(n_6115)
);

HB1xp67_ASAP7_75t_L g6116 ( 
.A(n_5941),
.Y(n_6116)
);

AND2x2_ASAP7_75t_L g6117 ( 
.A(n_5985),
.B(n_471),
.Y(n_6117)
);

INVxp67_ASAP7_75t_SL g6118 ( 
.A(n_6043),
.Y(n_6118)
);

AND2x2_ASAP7_75t_L g6119 ( 
.A(n_5992),
.B(n_471),
.Y(n_6119)
);

OR2x2_ASAP7_75t_L g6120 ( 
.A(n_6029),
.B(n_471),
.Y(n_6120)
);

AND2x4_ASAP7_75t_L g6121 ( 
.A(n_6037),
.B(n_5012),
.Y(n_6121)
);

HB1xp67_ASAP7_75t_L g6122 ( 
.A(n_5925),
.Y(n_6122)
);

INVx2_ASAP7_75t_L g6123 ( 
.A(n_5946),
.Y(n_6123)
);

OR2x2_ASAP7_75t_L g6124 ( 
.A(n_5986),
.B(n_472),
.Y(n_6124)
);

AND2x2_ASAP7_75t_L g6125 ( 
.A(n_6042),
.B(n_472),
.Y(n_6125)
);

INVx2_ASAP7_75t_L g6126 ( 
.A(n_5956),
.Y(n_6126)
);

INVx2_ASAP7_75t_L g6127 ( 
.A(n_5959),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_6016),
.Y(n_6128)
);

INVx1_ASAP7_75t_SL g6129 ( 
.A(n_5967),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5925),
.Y(n_6130)
);

AND2x2_ASAP7_75t_L g6131 ( 
.A(n_6063),
.B(n_472),
.Y(n_6131)
);

AND2x2_ASAP7_75t_L g6132 ( 
.A(n_6063),
.B(n_473),
.Y(n_6132)
);

INVx3_ASAP7_75t_L g6133 ( 
.A(n_5955),
.Y(n_6133)
);

OR2x2_ASAP7_75t_L g6134 ( 
.A(n_6004),
.B(n_473),
.Y(n_6134)
);

AOI22xp33_ASAP7_75t_L g6135 ( 
.A1(n_6058),
.A2(n_5019),
.B1(n_4739),
.B2(n_476),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_5942),
.Y(n_6136)
);

HB1xp67_ASAP7_75t_L g6137 ( 
.A(n_5931),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_5945),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_L g6139 ( 
.A(n_6007),
.B(n_474),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5960),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5953),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_5950),
.B(n_474),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5962),
.Y(n_6143)
);

INVx2_ASAP7_75t_L g6144 ( 
.A(n_5965),
.Y(n_6144)
);

NAND2xp5_ASAP7_75t_L g6145 ( 
.A(n_6018),
.B(n_475),
.Y(n_6145)
);

NAND2xp5_ASAP7_75t_L g6146 ( 
.A(n_6006),
.B(n_475),
.Y(n_6146)
);

NAND2xp5_ASAP7_75t_L g6147 ( 
.A(n_6038),
.B(n_476),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5966),
.Y(n_6148)
);

AND2x4_ASAP7_75t_L g6149 ( 
.A(n_5955),
.B(n_476),
.Y(n_6149)
);

OR2x2_ASAP7_75t_L g6150 ( 
.A(n_6023),
.B(n_477),
.Y(n_6150)
);

INVx2_ASAP7_75t_SL g6151 ( 
.A(n_6039),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_5973),
.Y(n_6152)
);

OR2x2_ASAP7_75t_L g6153 ( 
.A(n_6026),
.B(n_477),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_6064),
.B(n_477),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_5974),
.Y(n_6155)
);

INVx2_ASAP7_75t_L g6156 ( 
.A(n_5979),
.Y(n_6156)
);

HB1xp67_ASAP7_75t_L g6157 ( 
.A(n_5931),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5968),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_5969),
.Y(n_6159)
);

AND2x4_ASAP7_75t_L g6160 ( 
.A(n_6035),
.B(n_478),
.Y(n_6160)
);

OR2x2_ASAP7_75t_L g6161 ( 
.A(n_6032),
.B(n_478),
.Y(n_6161)
);

AND2x2_ASAP7_75t_L g6162 ( 
.A(n_6066),
.B(n_478),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_5970),
.Y(n_6163)
);

INVx2_ASAP7_75t_L g6164 ( 
.A(n_5981),
.Y(n_6164)
);

AND2x2_ASAP7_75t_L g6165 ( 
.A(n_6015),
.B(n_479),
.Y(n_6165)
);

INVx2_ASAP7_75t_L g6166 ( 
.A(n_6013),
.Y(n_6166)
);

INVxp67_ASAP7_75t_L g6167 ( 
.A(n_6040),
.Y(n_6167)
);

BUFx3_ASAP7_75t_L g6168 ( 
.A(n_6040),
.Y(n_6168)
);

AND2x2_ASAP7_75t_L g6169 ( 
.A(n_6017),
.B(n_479),
.Y(n_6169)
);

OR2x2_ASAP7_75t_L g6170 ( 
.A(n_5977),
.B(n_479),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_5978),
.Y(n_6171)
);

OR2x2_ASAP7_75t_L g6172 ( 
.A(n_5980),
.B(n_5984),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_6059),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_6036),
.B(n_480),
.Y(n_6174)
);

INVx2_ASAP7_75t_L g6175 ( 
.A(n_5998),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_5963),
.B(n_480),
.Y(n_6176)
);

INVx2_ASAP7_75t_L g6177 ( 
.A(n_6009),
.Y(n_6177)
);

HB1xp67_ASAP7_75t_L g6178 ( 
.A(n_6059),
.Y(n_6178)
);

HB1xp67_ASAP7_75t_L g6179 ( 
.A(n_6033),
.Y(n_6179)
);

BUFx2_ASAP7_75t_L g6180 ( 
.A(n_5923),
.Y(n_6180)
);

INVx1_ASAP7_75t_L g6181 ( 
.A(n_5989),
.Y(n_6181)
);

INVx2_ASAP7_75t_L g6182 ( 
.A(n_6010),
.Y(n_6182)
);

HB1xp67_ASAP7_75t_L g6183 ( 
.A(n_6031),
.Y(n_6183)
);

INVx2_ASAP7_75t_L g6184 ( 
.A(n_6020),
.Y(n_6184)
);

INVx2_ASAP7_75t_SL g6185 ( 
.A(n_5940),
.Y(n_6185)
);

OR2x2_ASAP7_75t_L g6186 ( 
.A(n_5990),
.B(n_480),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_6019),
.B(n_481),
.Y(n_6187)
);

INVx1_ASAP7_75t_L g6188 ( 
.A(n_5993),
.Y(n_6188)
);

INVx2_ASAP7_75t_L g6189 ( 
.A(n_6011),
.Y(n_6189)
);

HB1xp67_ASAP7_75t_L g6190 ( 
.A(n_6014),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5994),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_5995),
.Y(n_6192)
);

NAND2xp5_ASAP7_75t_L g6193 ( 
.A(n_6024),
.B(n_481),
.Y(n_6193)
);

HB1xp67_ASAP7_75t_L g6194 ( 
.A(n_5999),
.Y(n_6194)
);

OAI22xp5_ASAP7_75t_L g6195 ( 
.A1(n_5923),
.A2(n_5975),
.B1(n_5983),
.B2(n_6048),
.Y(n_6195)
);

INVx2_ASAP7_75t_L g6196 ( 
.A(n_6034),
.Y(n_6196)
);

NAND2xp5_ASAP7_75t_L g6197 ( 
.A(n_6003),
.B(n_6067),
.Y(n_6197)
);

NAND2xp5_ASAP7_75t_L g6198 ( 
.A(n_6067),
.B(n_481),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_5929),
.Y(n_6199)
);

OR2x2_ASAP7_75t_L g6200 ( 
.A(n_5988),
.B(n_482),
.Y(n_6200)
);

AND3x1_ASAP7_75t_L g6201 ( 
.A(n_6047),
.B(n_4739),
.C(n_483),
.Y(n_6201)
);

AND2x2_ASAP7_75t_L g6202 ( 
.A(n_5957),
.B(n_6048),
.Y(n_6202)
);

BUFx2_ASAP7_75t_L g6203 ( 
.A(n_6045),
.Y(n_6203)
);

INVx2_ASAP7_75t_L g6204 ( 
.A(n_5934),
.Y(n_6204)
);

NOR2xp33_ASAP7_75t_SL g6205 ( 
.A(n_5991),
.B(n_483),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_6044),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_6027),
.B(n_483),
.Y(n_6207)
);

INVx2_ASAP7_75t_L g6208 ( 
.A(n_5991),
.Y(n_6208)
);

AND2x2_ASAP7_75t_L g6209 ( 
.A(n_6045),
.B(n_484),
.Y(n_6209)
);

BUFx3_ASAP7_75t_L g6210 ( 
.A(n_6008),
.Y(n_6210)
);

AND2x2_ASAP7_75t_L g6211 ( 
.A(n_5930),
.B(n_484),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_6046),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_6008),
.Y(n_6213)
);

BUFx3_ASAP7_75t_L g6214 ( 
.A(n_6041),
.Y(n_6214)
);

AND2x2_ASAP7_75t_L g6215 ( 
.A(n_6012),
.B(n_485),
.Y(n_6215)
);

AND2x4_ASAP7_75t_L g6216 ( 
.A(n_6062),
.B(n_485),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_5938),
.B(n_485),
.Y(n_6217)
);

OR2x2_ASAP7_75t_L g6218 ( 
.A(n_5958),
.B(n_486),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_5928),
.Y(n_6219)
);

INVx2_ASAP7_75t_L g6220 ( 
.A(n_5987),
.Y(n_6220)
);

AND2x2_ASAP7_75t_L g6221 ( 
.A(n_5964),
.B(n_486),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_6061),
.Y(n_6222)
);

HB1xp67_ASAP7_75t_L g6223 ( 
.A(n_6022),
.Y(n_6223)
);

AND2x4_ASAP7_75t_L g6224 ( 
.A(n_5976),
.B(n_486),
.Y(n_6224)
);

INVxp67_ASAP7_75t_SL g6225 ( 
.A(n_6060),
.Y(n_6225)
);

INVx1_ASAP7_75t_L g6226 ( 
.A(n_5924),
.Y(n_6226)
);

INVx2_ASAP7_75t_SL g6227 ( 
.A(n_6053),
.Y(n_6227)
);

INVx2_ASAP7_75t_L g6228 ( 
.A(n_6060),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_6060),
.Y(n_6229)
);

AND2x2_ASAP7_75t_L g6230 ( 
.A(n_5932),
.B(n_487),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5924),
.Y(n_6231)
);

BUFx3_ASAP7_75t_L g6232 ( 
.A(n_6053),
.Y(n_6232)
);

AND2x2_ASAP7_75t_L g6233 ( 
.A(n_5932),
.B(n_488),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_6072),
.Y(n_6234)
);

AND2x2_ASAP7_75t_L g6235 ( 
.A(n_6075),
.B(n_488),
.Y(n_6235)
);

INVx2_ASAP7_75t_SL g6236 ( 
.A(n_6232),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_6072),
.Y(n_6237)
);

NAND2xp5_ASAP7_75t_L g6238 ( 
.A(n_6073),
.B(n_488),
.Y(n_6238)
);

INVx2_ASAP7_75t_L g6239 ( 
.A(n_6077),
.Y(n_6239)
);

NAND2xp5_ASAP7_75t_L g6240 ( 
.A(n_6222),
.B(n_489),
.Y(n_6240)
);

AND2x2_ASAP7_75t_L g6241 ( 
.A(n_6068),
.B(n_489),
.Y(n_6241)
);

NAND2xp5_ASAP7_75t_L g6242 ( 
.A(n_6169),
.B(n_489),
.Y(n_6242)
);

BUFx6f_ASAP7_75t_L g6243 ( 
.A(n_6133),
.Y(n_6243)
);

NAND2x1p5_ASAP7_75t_L g6244 ( 
.A(n_6149),
.B(n_1008),
.Y(n_6244)
);

INVx2_ASAP7_75t_L g6245 ( 
.A(n_6083),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_6074),
.Y(n_6246)
);

AND2x4_ASAP7_75t_L g6247 ( 
.A(n_6133),
.B(n_490),
.Y(n_6247)
);

AND2x2_ASAP7_75t_L g6248 ( 
.A(n_6225),
.B(n_491),
.Y(n_6248)
);

BUFx6f_ASAP7_75t_L g6249 ( 
.A(n_6151),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_6074),
.Y(n_6250)
);

HB1xp67_ASAP7_75t_L g6251 ( 
.A(n_6183),
.Y(n_6251)
);

HB1xp67_ASAP7_75t_L g6252 ( 
.A(n_6179),
.Y(n_6252)
);

AND2x4_ASAP7_75t_L g6253 ( 
.A(n_6227),
.B(n_491),
.Y(n_6253)
);

AND2x4_ASAP7_75t_L g6254 ( 
.A(n_6129),
.B(n_492),
.Y(n_6254)
);

AOI22xp33_ASAP7_75t_L g6255 ( 
.A1(n_6090),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_6255)
);

INVx1_ASAP7_75t_SL g6256 ( 
.A(n_6149),
.Y(n_6256)
);

HB1xp67_ASAP7_75t_L g6257 ( 
.A(n_6079),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6118),
.B(n_492),
.Y(n_6258)
);

OR2x2_ASAP7_75t_L g6259 ( 
.A(n_6069),
.B(n_494),
.Y(n_6259)
);

AND2x2_ASAP7_75t_L g6260 ( 
.A(n_6228),
.B(n_494),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_6095),
.Y(n_6261)
);

AND2x2_ASAP7_75t_L g6262 ( 
.A(n_6229),
.B(n_495),
.Y(n_6262)
);

AND2x2_ASAP7_75t_L g6263 ( 
.A(n_6110),
.B(n_495),
.Y(n_6263)
);

AND2x2_ASAP7_75t_L g6264 ( 
.A(n_6104),
.B(n_495),
.Y(n_6264)
);

BUFx5_ASAP7_75t_L g6265 ( 
.A(n_6224),
.Y(n_6265)
);

INVx2_ASAP7_75t_L g6266 ( 
.A(n_6102),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_6190),
.Y(n_6267)
);

AND2x2_ASAP7_75t_L g6268 ( 
.A(n_6104),
.B(n_496),
.Y(n_6268)
);

AND2x2_ASAP7_75t_L g6269 ( 
.A(n_6088),
.B(n_496),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_6230),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_6233),
.Y(n_6271)
);

AND2x2_ASAP7_75t_L g6272 ( 
.A(n_6085),
.B(n_497),
.Y(n_6272)
);

AND2x2_ASAP7_75t_L g6273 ( 
.A(n_6168),
.B(n_497),
.Y(n_6273)
);

INVx2_ASAP7_75t_L g6274 ( 
.A(n_6224),
.Y(n_6274)
);

INVx2_ASAP7_75t_L g6275 ( 
.A(n_6184),
.Y(n_6275)
);

INVx2_ASAP7_75t_L g6276 ( 
.A(n_6199),
.Y(n_6276)
);

NOR2x1_ASAP7_75t_SL g6277 ( 
.A(n_6195),
.B(n_498),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_6174),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_6204),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_6078),
.Y(n_6280)
);

AND2x2_ASAP7_75t_L g6281 ( 
.A(n_6185),
.B(n_497),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_6226),
.Y(n_6282)
);

AND2x2_ASAP7_75t_L g6283 ( 
.A(n_6114),
.B(n_6176),
.Y(n_6283)
);

BUFx3_ASAP7_75t_L g6284 ( 
.A(n_6117),
.Y(n_6284)
);

OR2x2_ASAP7_75t_L g6285 ( 
.A(n_6231),
.B(n_498),
.Y(n_6285)
);

HB1xp67_ASAP7_75t_L g6286 ( 
.A(n_6097),
.Y(n_6286)
);

NOR2xp33_ASAP7_75t_L g6287 ( 
.A(n_6071),
.B(n_498),
.Y(n_6287)
);

INVx3_ASAP7_75t_L g6288 ( 
.A(n_6210),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6112),
.Y(n_6289)
);

BUFx2_ASAP7_75t_L g6290 ( 
.A(n_6180),
.Y(n_6290)
);

AND2x4_ASAP7_75t_L g6291 ( 
.A(n_6167),
.B(n_499),
.Y(n_6291)
);

INVx3_ASAP7_75t_SL g6292 ( 
.A(n_6160),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_6115),
.Y(n_6293)
);

HB1xp67_ASAP7_75t_L g6294 ( 
.A(n_6098),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_6214),
.B(n_499),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_6089),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6122),
.Y(n_6297)
);

HB1xp67_ASAP7_75t_L g6298 ( 
.A(n_6116),
.Y(n_6298)
);

INVx5_ASAP7_75t_L g6299 ( 
.A(n_6209),
.Y(n_6299)
);

INVx2_ASAP7_75t_L g6300 ( 
.A(n_6106),
.Y(n_6300)
);

INVx2_ASAP7_75t_L g6301 ( 
.A(n_6108),
.Y(n_6301)
);

INVx2_ASAP7_75t_L g6302 ( 
.A(n_6123),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_6137),
.Y(n_6303)
);

AND2x2_ASAP7_75t_L g6304 ( 
.A(n_6082),
.B(n_499),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_6126),
.Y(n_6305)
);

BUFx3_ASAP7_75t_L g6306 ( 
.A(n_6119),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_6157),
.Y(n_6307)
);

INVx3_ASAP7_75t_L g6308 ( 
.A(n_6160),
.Y(n_6308)
);

BUFx2_ASAP7_75t_L g6309 ( 
.A(n_6211),
.Y(n_6309)
);

AND2x4_ASAP7_75t_L g6310 ( 
.A(n_6208),
.B(n_500),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_6178),
.Y(n_6311)
);

BUFx2_ASAP7_75t_L g6312 ( 
.A(n_6203),
.Y(n_6312)
);

CKINVDCx5p33_ASAP7_75t_R g6313 ( 
.A(n_6221),
.Y(n_6313)
);

INVx2_ASAP7_75t_L g6314 ( 
.A(n_6127),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6194),
.Y(n_6315)
);

OR2x2_ASAP7_75t_L g6316 ( 
.A(n_6107),
.B(n_500),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_6109),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6131),
.Y(n_6318)
);

INVx4_ASAP7_75t_L g6319 ( 
.A(n_6103),
.Y(n_6319)
);

HB1xp67_ASAP7_75t_L g6320 ( 
.A(n_6081),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_6132),
.Y(n_6321)
);

AND2x2_ASAP7_75t_L g6322 ( 
.A(n_6070),
.B(n_501),
.Y(n_6322)
);

HB1xp67_ASAP7_75t_L g6323 ( 
.A(n_6094),
.Y(n_6323)
);

BUFx2_ASAP7_75t_L g6324 ( 
.A(n_6111),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6153),
.Y(n_6325)
);

AND2x2_ASAP7_75t_L g6326 ( 
.A(n_6213),
.B(n_6154),
.Y(n_6326)
);

AND2x2_ASAP7_75t_L g6327 ( 
.A(n_6162),
.B(n_501),
.Y(n_6327)
);

INVxp67_ASAP7_75t_SL g6328 ( 
.A(n_6142),
.Y(n_6328)
);

INVx2_ASAP7_75t_L g6329 ( 
.A(n_6144),
.Y(n_6329)
);

AND2x2_ASAP7_75t_L g6330 ( 
.A(n_6093),
.B(n_501),
.Y(n_6330)
);

OR2x2_ASAP7_75t_L g6331 ( 
.A(n_6212),
.B(n_502),
.Y(n_6331)
);

AND2x2_ASAP7_75t_L g6332 ( 
.A(n_6165),
.B(n_502),
.Y(n_6332)
);

AND2x2_ASAP7_75t_L g6333 ( 
.A(n_6091),
.B(n_502),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_6161),
.Y(n_6334)
);

AND2x4_ASAP7_75t_L g6335 ( 
.A(n_6086),
.B(n_503),
.Y(n_6335)
);

INVx3_ASAP7_75t_L g6336 ( 
.A(n_6152),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_6155),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_6206),
.Y(n_6338)
);

AND2x2_ASAP7_75t_L g6339 ( 
.A(n_6215),
.B(n_503),
.Y(n_6339)
);

INVx2_ASAP7_75t_L g6340 ( 
.A(n_6156),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6128),
.Y(n_6341)
);

BUFx3_ASAP7_75t_L g6342 ( 
.A(n_6125),
.Y(n_6342)
);

AND2x2_ASAP7_75t_L g6343 ( 
.A(n_6189),
.B(n_504),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_6101),
.Y(n_6344)
);

OR2x2_ASAP7_75t_L g6345 ( 
.A(n_6218),
.B(n_504),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_6220),
.B(n_504),
.Y(n_6346)
);

AND2x4_ASAP7_75t_L g6347 ( 
.A(n_6121),
.B(n_6216),
.Y(n_6347)
);

AND2x2_ASAP7_75t_L g6348 ( 
.A(n_6202),
.B(n_505),
.Y(n_6348)
);

AND2x2_ASAP7_75t_L g6349 ( 
.A(n_6223),
.B(n_505),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_6164),
.Y(n_6350)
);

BUFx3_ASAP7_75t_L g6351 ( 
.A(n_6100),
.Y(n_6351)
);

AND2x2_ASAP7_75t_L g6352 ( 
.A(n_6217),
.B(n_505),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_6166),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6124),
.B(n_506),
.Y(n_6354)
);

INVxp67_ASAP7_75t_L g6355 ( 
.A(n_6205),
.Y(n_6355)
);

BUFx2_ASAP7_75t_L g6356 ( 
.A(n_6111),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_6177),
.Y(n_6357)
);

AND2x2_ASAP7_75t_L g6358 ( 
.A(n_6120),
.B(n_506),
.Y(n_6358)
);

BUFx2_ASAP7_75t_L g6359 ( 
.A(n_6111),
.Y(n_6359)
);

OR2x2_ASAP7_75t_L g6360 ( 
.A(n_6198),
.B(n_506),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_6182),
.Y(n_6361)
);

NAND2xp5_ASAP7_75t_L g6362 ( 
.A(n_6197),
.B(n_507),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6121),
.B(n_507),
.Y(n_6363)
);

OR2x2_ASAP7_75t_L g6364 ( 
.A(n_6139),
.B(n_507),
.Y(n_6364)
);

INVx3_ASAP7_75t_L g6365 ( 
.A(n_6175),
.Y(n_6365)
);

INVx2_ASAP7_75t_L g6366 ( 
.A(n_6196),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_6092),
.Y(n_6367)
);

NAND2xp5_ASAP7_75t_L g6368 ( 
.A(n_6146),
.B(n_6145),
.Y(n_6368)
);

INVxp67_ASAP7_75t_SL g6369 ( 
.A(n_6147),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_6080),
.Y(n_6370)
);

CKINVDCx5p33_ASAP7_75t_R g6371 ( 
.A(n_6207),
.Y(n_6371)
);

OR2x2_ASAP7_75t_L g6372 ( 
.A(n_6105),
.B(n_508),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_6200),
.B(n_6150),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_6076),
.Y(n_6374)
);

INVx2_ASAP7_75t_L g6375 ( 
.A(n_6216),
.Y(n_6375)
);

OR2x2_ASAP7_75t_L g6376 ( 
.A(n_6187),
.B(n_508),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_6172),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6134),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_6130),
.Y(n_6379)
);

HB1xp67_ASAP7_75t_L g6380 ( 
.A(n_6113),
.Y(n_6380)
);

INVx1_ASAP7_75t_SL g6381 ( 
.A(n_6170),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_6186),
.B(n_508),
.Y(n_6382)
);

AND2x2_ASAP7_75t_L g6383 ( 
.A(n_6096),
.B(n_509),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_6136),
.B(n_509),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6130),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_6235),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6258),
.Y(n_6387)
);

BUFx3_ASAP7_75t_L g6388 ( 
.A(n_6249),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_SL g6389 ( 
.A(n_6249),
.B(n_6219),
.Y(n_6389)
);

BUFx6f_ASAP7_75t_L g6390 ( 
.A(n_6243),
.Y(n_6390)
);

BUFx2_ASAP7_75t_L g6391 ( 
.A(n_6236),
.Y(n_6391)
);

OA21x2_ASAP7_75t_L g6392 ( 
.A1(n_6312),
.A2(n_6193),
.B(n_6173),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_6252),
.Y(n_6393)
);

AOI21xp33_ASAP7_75t_L g6394 ( 
.A1(n_6243),
.A2(n_6181),
.B(n_6158),
.Y(n_6394)
);

INVx4_ASAP7_75t_SL g6395 ( 
.A(n_6292),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_6247),
.Y(n_6396)
);

INVx2_ASAP7_75t_L g6397 ( 
.A(n_6247),
.Y(n_6397)
);

AOI21xp5_ASAP7_75t_L g6398 ( 
.A1(n_6277),
.A2(n_6181),
.B(n_6140),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6241),
.Y(n_6399)
);

AND2x4_ASAP7_75t_L g6400 ( 
.A(n_6288),
.B(n_6138),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_6248),
.Y(n_6401)
);

HB1xp67_ASAP7_75t_L g6402 ( 
.A(n_6251),
.Y(n_6402)
);

OAI21xp33_ASAP7_75t_L g6403 ( 
.A1(n_6351),
.A2(n_6143),
.B(n_6141),
.Y(n_6403)
);

NAND3xp33_ASAP7_75t_SL g6404 ( 
.A(n_6290),
.B(n_6135),
.C(n_6173),
.Y(n_6404)
);

INVx3_ASAP7_75t_L g6405 ( 
.A(n_6253),
.Y(n_6405)
);

AOI21xp5_ASAP7_75t_L g6406 ( 
.A1(n_6362),
.A2(n_6159),
.B(n_6148),
.Y(n_6406)
);

INVx2_ASAP7_75t_L g6407 ( 
.A(n_6272),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_6281),
.Y(n_6408)
);

HB1xp67_ASAP7_75t_L g6409 ( 
.A(n_6276),
.Y(n_6409)
);

OA21x2_ASAP7_75t_L g6410 ( 
.A1(n_6312),
.A2(n_6171),
.B(n_6163),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6348),
.B(n_6188),
.Y(n_6411)
);

INVx2_ASAP7_75t_L g6412 ( 
.A(n_6264),
.Y(n_6412)
);

OA21x2_ASAP7_75t_L g6413 ( 
.A1(n_6324),
.A2(n_6192),
.B(n_6191),
.Y(n_6413)
);

HB1xp67_ASAP7_75t_L g6414 ( 
.A(n_6279),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_6268),
.Y(n_6415)
);

INVx4_ASAP7_75t_SL g6416 ( 
.A(n_6254),
.Y(n_6416)
);

OR2x6_ASAP7_75t_L g6417 ( 
.A(n_6244),
.B(n_6099),
.Y(n_6417)
);

BUFx2_ASAP7_75t_L g6418 ( 
.A(n_6298),
.Y(n_6418)
);

OAI21xp5_ASAP7_75t_L g6419 ( 
.A1(n_6355),
.A2(n_6087),
.B(n_6201),
.Y(n_6419)
);

OR2x2_ASAP7_75t_SL g6420 ( 
.A(n_6257),
.B(n_6084),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_6269),
.Y(n_6421)
);

INVxp67_ASAP7_75t_L g6422 ( 
.A(n_6290),
.Y(n_6422)
);

A2O1A1Ixp33_ASAP7_75t_L g6423 ( 
.A1(n_6328),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6263),
.Y(n_6424)
);

BUFx2_ASAP7_75t_L g6425 ( 
.A(n_6284),
.Y(n_6425)
);

AND4x1_ASAP7_75t_L g6426 ( 
.A(n_6255),
.B(n_514),
.C(n_512),
.D(n_513),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_6286),
.Y(n_6427)
);

BUFx6f_ASAP7_75t_L g6428 ( 
.A(n_6273),
.Y(n_6428)
);

AND2x2_ASAP7_75t_L g6429 ( 
.A(n_6299),
.B(n_512),
.Y(n_6429)
);

INVx2_ASAP7_75t_L g6430 ( 
.A(n_6336),
.Y(n_6430)
);

INVx2_ASAP7_75t_L g6431 ( 
.A(n_6365),
.Y(n_6431)
);

A2O1A1Ixp33_ASAP7_75t_L g6432 ( 
.A1(n_6299),
.A2(n_516),
.B(n_512),
.C(n_515),
.Y(n_6432)
);

OR2x2_ASAP7_75t_L g6433 ( 
.A(n_6240),
.B(n_516),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6294),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6291),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6291),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_6239),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_6245),
.Y(n_6438)
);

OA21x2_ASAP7_75t_L g6439 ( 
.A1(n_6324),
.A2(n_517),
.B(n_518),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6274),
.Y(n_6440)
);

INVx8_ASAP7_75t_L g6441 ( 
.A(n_6310),
.Y(n_6441)
);

AOI21xp5_ASAP7_75t_L g6442 ( 
.A1(n_6256),
.A2(n_6346),
.B(n_6313),
.Y(n_6442)
);

OR2x2_ASAP7_75t_L g6443 ( 
.A(n_6267),
.B(n_6270),
.Y(n_6443)
);

INVx2_ASAP7_75t_L g6444 ( 
.A(n_6261),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6266),
.Y(n_6445)
);

OR2x2_ASAP7_75t_L g6446 ( 
.A(n_6271),
.B(n_517),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_6299),
.B(n_517),
.Y(n_6447)
);

AND2x2_ASAP7_75t_L g6448 ( 
.A(n_6319),
.B(n_518),
.Y(n_6448)
);

HB1xp67_ASAP7_75t_L g6449 ( 
.A(n_6275),
.Y(n_6449)
);

NAND3xp33_ASAP7_75t_SL g6450 ( 
.A(n_6356),
.B(n_6359),
.C(n_6383),
.Y(n_6450)
);

INVx1_ASAP7_75t_L g6451 ( 
.A(n_6238),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_6295),
.Y(n_6452)
);

BUFx2_ASAP7_75t_L g6453 ( 
.A(n_6306),
.Y(n_6453)
);

AOI21xp5_ASAP7_75t_L g6454 ( 
.A1(n_6368),
.A2(n_518),
.B(n_519),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_6309),
.B(n_519),
.Y(n_6455)
);

INVx2_ASAP7_75t_L g6456 ( 
.A(n_6310),
.Y(n_6456)
);

INVxp67_ASAP7_75t_SL g6457 ( 
.A(n_6345),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6356),
.Y(n_6458)
);

INVx2_ASAP7_75t_L g6459 ( 
.A(n_6265),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6359),
.Y(n_6460)
);

OR2x2_ASAP7_75t_L g6461 ( 
.A(n_6278),
.B(n_519),
.Y(n_6461)
);

OR2x2_ASAP7_75t_L g6462 ( 
.A(n_6289),
.B(n_520),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_6293),
.Y(n_6463)
);

OAI21xp5_ASAP7_75t_L g6464 ( 
.A1(n_6315),
.A2(n_520),
.B(n_521),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6320),
.Y(n_6465)
);

INVx1_ASAP7_75t_SL g6466 ( 
.A(n_6260),
.Y(n_6466)
);

INVx2_ASAP7_75t_L g6467 ( 
.A(n_6265),
.Y(n_6467)
);

INVx2_ASAP7_75t_L g6468 ( 
.A(n_6265),
.Y(n_6468)
);

INVx1_ASAP7_75t_SL g6469 ( 
.A(n_6262),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_6323),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_6352),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_6349),
.B(n_521),
.Y(n_6472)
);

INVx3_ASAP7_75t_L g6473 ( 
.A(n_6347),
.Y(n_6473)
);

BUFx2_ASAP7_75t_L g6474 ( 
.A(n_6265),
.Y(n_6474)
);

BUFx3_ASAP7_75t_L g6475 ( 
.A(n_6363),
.Y(n_6475)
);

OAI211xp5_ASAP7_75t_L g6476 ( 
.A1(n_6297),
.A2(n_524),
.B(n_522),
.C(n_523),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6360),
.Y(n_6477)
);

BUFx2_ASAP7_75t_L g6478 ( 
.A(n_6342),
.Y(n_6478)
);

HB1xp67_ASAP7_75t_L g6479 ( 
.A(n_6300),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_6380),
.Y(n_6480)
);

OAI21xp5_ASAP7_75t_SL g6481 ( 
.A1(n_6309),
.A2(n_522),
.B(n_523),
.Y(n_6481)
);

NAND2xp5_ASAP7_75t_L g6482 ( 
.A(n_6304),
.B(n_522),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_6316),
.Y(n_6483)
);

INVx3_ASAP7_75t_L g6484 ( 
.A(n_6347),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6301),
.Y(n_6485)
);

BUFx2_ASAP7_75t_L g6486 ( 
.A(n_6308),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6302),
.Y(n_6487)
);

AND2x2_ASAP7_75t_L g6488 ( 
.A(n_6333),
.B(n_523),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_6375),
.Y(n_6489)
);

INVx2_ASAP7_75t_SL g6490 ( 
.A(n_6305),
.Y(n_6490)
);

NAND4xp25_ASAP7_75t_L g6491 ( 
.A(n_6303),
.B(n_526),
.C(n_524),
.D(n_525),
.Y(n_6491)
);

INVx2_ASAP7_75t_L g6492 ( 
.A(n_6314),
.Y(n_6492)
);

INVx1_ASAP7_75t_SL g6493 ( 
.A(n_6343),
.Y(n_6493)
);

NAND2xp5_ASAP7_75t_L g6494 ( 
.A(n_6322),
.B(n_524),
.Y(n_6494)
);

OA21x2_ASAP7_75t_L g6495 ( 
.A1(n_6234),
.A2(n_525),
.B(n_526),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_6329),
.Y(n_6496)
);

INVx3_ASAP7_75t_L g6497 ( 
.A(n_6337),
.Y(n_6497)
);

NAND4xp25_ASAP7_75t_L g6498 ( 
.A(n_6307),
.B(n_529),
.C(n_527),
.D(n_528),
.Y(n_6498)
);

AND2x2_ASAP7_75t_L g6499 ( 
.A(n_6326),
.B(n_527),
.Y(n_6499)
);

OAI21xp5_ASAP7_75t_L g6500 ( 
.A1(n_6280),
.A2(n_527),
.B(n_528),
.Y(n_6500)
);

A2O1A1Ixp33_ASAP7_75t_L g6501 ( 
.A1(n_6283),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6340),
.Y(n_6502)
);

OR2x6_ASAP7_75t_L g6503 ( 
.A(n_6335),
.B(n_529),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6350),
.Y(n_6504)
);

NAND3xp33_ASAP7_75t_L g6505 ( 
.A(n_6237),
.B(n_530),
.C(n_531),
.Y(n_6505)
);

AND2x4_ASAP7_75t_L g6506 ( 
.A(n_6335),
.B(n_530),
.Y(n_6506)
);

NAND2xp5_ASAP7_75t_SL g6507 ( 
.A(n_6366),
.B(n_531),
.Y(n_6507)
);

INVxp67_ASAP7_75t_L g6508 ( 
.A(n_6287),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_6330),
.B(n_532),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6353),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6357),
.Y(n_6511)
);

OAI21xp33_ASAP7_75t_L g6512 ( 
.A1(n_6367),
.A2(n_6344),
.B(n_6370),
.Y(n_6512)
);

AO21x1_ASAP7_75t_L g6513 ( 
.A1(n_6246),
.A2(n_534),
.B(n_533),
.Y(n_6513)
);

AOI21xp33_ASAP7_75t_L g6514 ( 
.A1(n_6372),
.A2(n_532),
.B(n_533),
.Y(n_6514)
);

INVx2_ASAP7_75t_L g6515 ( 
.A(n_6361),
.Y(n_6515)
);

OR2x6_ASAP7_75t_L g6516 ( 
.A(n_6364),
.B(n_532),
.Y(n_6516)
);

INVx2_ASAP7_75t_L g6517 ( 
.A(n_6250),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_6259),
.Y(n_6518)
);

NAND2xp5_ASAP7_75t_L g6519 ( 
.A(n_6369),
.B(n_6373),
.Y(n_6519)
);

NOR2xp33_ASAP7_75t_L g6520 ( 
.A(n_6371),
.B(n_534),
.Y(n_6520)
);

NAND2xp5_ASAP7_75t_L g6521 ( 
.A(n_6381),
.B(n_535),
.Y(n_6521)
);

INVx2_ASAP7_75t_SL g6522 ( 
.A(n_6332),
.Y(n_6522)
);

INVx2_ASAP7_75t_L g6523 ( 
.A(n_6282),
.Y(n_6523)
);

HB1xp67_ASAP7_75t_L g6524 ( 
.A(n_6311),
.Y(n_6524)
);

INVx4_ASAP7_75t_L g6525 ( 
.A(n_6376),
.Y(n_6525)
);

INVx1_ASAP7_75t_L g6526 ( 
.A(n_6285),
.Y(n_6526)
);

A2O1A1Ixp33_ASAP7_75t_L g6527 ( 
.A1(n_6377),
.A2(n_537),
.B(n_535),
.C(n_536),
.Y(n_6527)
);

INVx2_ASAP7_75t_L g6528 ( 
.A(n_6341),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6318),
.B(n_535),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_6296),
.Y(n_6530)
);

OR2x2_ASAP7_75t_L g6531 ( 
.A(n_6374),
.B(n_536),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6321),
.B(n_6384),
.Y(n_6532)
);

INVx1_ASAP7_75t_SL g6533 ( 
.A(n_6339),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_6325),
.Y(n_6534)
);

AOI21xp5_ASAP7_75t_L g6535 ( 
.A1(n_6242),
.A2(n_6317),
.B(n_6334),
.Y(n_6535)
);

A2O1A1Ixp33_ASAP7_75t_L g6536 ( 
.A1(n_6338),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_6536)
);

INVx2_ASAP7_75t_L g6537 ( 
.A(n_6331),
.Y(n_6537)
);

NAND2x1_ASAP7_75t_L g6538 ( 
.A(n_6378),
.B(n_538),
.Y(n_6538)
);

AND2x2_ASAP7_75t_L g6539 ( 
.A(n_6358),
.B(n_539),
.Y(n_6539)
);

AOI21xp5_ASAP7_75t_L g6540 ( 
.A1(n_6382),
.A2(n_539),
.B(n_540),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6354),
.Y(n_6541)
);

INVx3_ASAP7_75t_L g6542 ( 
.A(n_6327),
.Y(n_6542)
);

INVx2_ASAP7_75t_L g6543 ( 
.A(n_6379),
.Y(n_6543)
);

NAND2xp5_ASAP7_75t_L g6544 ( 
.A(n_6385),
.B(n_540),
.Y(n_6544)
);

NAND3xp33_ASAP7_75t_L g6545 ( 
.A(n_6243),
.B(n_541),
.C(n_542),
.Y(n_6545)
);

OR2x2_ASAP7_75t_L g6546 ( 
.A(n_6362),
.B(n_542),
.Y(n_6546)
);

AOI22xp5_ASAP7_75t_L g6547 ( 
.A1(n_6236),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_6547)
);

AND4x1_ASAP7_75t_L g6548 ( 
.A(n_6255),
.B(n_545),
.C(n_543),
.D(n_544),
.Y(n_6548)
);

BUFx3_ASAP7_75t_L g6549 ( 
.A(n_6249),
.Y(n_6549)
);

BUFx6f_ASAP7_75t_L g6550 ( 
.A(n_6249),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_6236),
.B(n_545),
.Y(n_6551)
);

INVx1_ASAP7_75t_SL g6552 ( 
.A(n_6292),
.Y(n_6552)
);

A2O1A1Ixp33_ASAP7_75t_L g6553 ( 
.A1(n_6236),
.A2(n_547),
.B(n_545),
.C(n_546),
.Y(n_6553)
);

INVx2_ASAP7_75t_L g6554 ( 
.A(n_6236),
.Y(n_6554)
);

INVx2_ASAP7_75t_SL g6555 ( 
.A(n_6249),
.Y(n_6555)
);

AOI21xp5_ASAP7_75t_L g6556 ( 
.A1(n_6236),
.A2(n_546),
.B(n_548),
.Y(n_6556)
);

A2O1A1Ixp33_ASAP7_75t_L g6557 ( 
.A1(n_6236),
.A2(n_549),
.B(n_546),
.C(n_548),
.Y(n_6557)
);

OR2x2_ASAP7_75t_L g6558 ( 
.A(n_6362),
.B(n_548),
.Y(n_6558)
);

AO21x2_ASAP7_75t_L g6559 ( 
.A1(n_6362),
.A2(n_549),
.B(n_550),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6235),
.Y(n_6560)
);

INVx2_ASAP7_75t_SL g6561 ( 
.A(n_6249),
.Y(n_6561)
);

AOI21xp5_ASAP7_75t_SL g6562 ( 
.A1(n_6277),
.A2(n_551),
.B(n_552),
.Y(n_6562)
);

INVx2_ASAP7_75t_L g6563 ( 
.A(n_6236),
.Y(n_6563)
);

INVxp67_ASAP7_75t_SL g6564 ( 
.A(n_6236),
.Y(n_6564)
);

INVxp67_ASAP7_75t_L g6565 ( 
.A(n_6236),
.Y(n_6565)
);

INVx2_ASAP7_75t_L g6566 ( 
.A(n_6236),
.Y(n_6566)
);

OA21x2_ASAP7_75t_L g6567 ( 
.A1(n_6312),
.A2(n_551),
.B(n_552),
.Y(n_6567)
);

OAI21xp5_ASAP7_75t_SL g6568 ( 
.A1(n_6288),
.A2(n_551),
.B(n_552),
.Y(n_6568)
);

AND2x2_ASAP7_75t_L g6569 ( 
.A(n_6236),
.B(n_553),
.Y(n_6569)
);

INVxp67_ASAP7_75t_SL g6570 ( 
.A(n_6236),
.Y(n_6570)
);

AOI21x1_ASAP7_75t_L g6571 ( 
.A1(n_6324),
.A2(n_553),
.B(n_554),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_6551),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6569),
.Y(n_6573)
);

INVx2_ASAP7_75t_L g6574 ( 
.A(n_6391),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6409),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6395),
.B(n_554),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_6395),
.B(n_554),
.Y(n_6577)
);

AND2x2_ASAP7_75t_L g6578 ( 
.A(n_6564),
.B(n_555),
.Y(n_6578)
);

NAND3xp33_ASAP7_75t_L g6579 ( 
.A(n_6565),
.B(n_555),
.C(n_556),
.Y(n_6579)
);

INVxp67_ASAP7_75t_SL g6580 ( 
.A(n_6570),
.Y(n_6580)
);

NAND3xp33_ASAP7_75t_L g6581 ( 
.A(n_6550),
.B(n_555),
.C(n_556),
.Y(n_6581)
);

AND2x4_ASAP7_75t_L g6582 ( 
.A(n_6388),
.B(n_557),
.Y(n_6582)
);

OR2x2_ASAP7_75t_L g6583 ( 
.A(n_6422),
.B(n_557),
.Y(n_6583)
);

NOR3xp33_ASAP7_75t_L g6584 ( 
.A(n_6555),
.B(n_560),
.C(n_559),
.Y(n_6584)
);

AND2x2_ASAP7_75t_L g6585 ( 
.A(n_6552),
.B(n_558),
.Y(n_6585)
);

NAND2xp5_ASAP7_75t_SL g6586 ( 
.A(n_6550),
.B(n_558),
.Y(n_6586)
);

NAND3xp33_ASAP7_75t_L g6587 ( 
.A(n_6390),
.B(n_559),
.C(n_560),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6554),
.B(n_561),
.Y(n_6588)
);

AND2x2_ASAP7_75t_L g6589 ( 
.A(n_6563),
.B(n_561),
.Y(n_6589)
);

NOR2xp33_ASAP7_75t_L g6590 ( 
.A(n_6566),
.B(n_561),
.Y(n_6590)
);

NAND2xp5_ASAP7_75t_L g6591 ( 
.A(n_6455),
.B(n_562),
.Y(n_6591)
);

OR2x2_ASAP7_75t_L g6592 ( 
.A(n_6489),
.B(n_562),
.Y(n_6592)
);

AND2x2_ASAP7_75t_L g6593 ( 
.A(n_6549),
.B(n_562),
.Y(n_6593)
);

OR2x2_ASAP7_75t_L g6594 ( 
.A(n_6440),
.B(n_563),
.Y(n_6594)
);

BUFx2_ASAP7_75t_L g6595 ( 
.A(n_6561),
.Y(n_6595)
);

NOR2x1_ASAP7_75t_L g6596 ( 
.A(n_6439),
.B(n_563),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_SL g6597 ( 
.A(n_6390),
.B(n_563),
.Y(n_6597)
);

NOR3xp33_ASAP7_75t_L g6598 ( 
.A(n_6450),
.B(n_566),
.C(n_565),
.Y(n_6598)
);

NAND2xp5_ASAP7_75t_L g6599 ( 
.A(n_6429),
.B(n_564),
.Y(n_6599)
);

OR2x2_ASAP7_75t_L g6600 ( 
.A(n_6418),
.B(n_564),
.Y(n_6600)
);

NAND2xp5_ASAP7_75t_L g6601 ( 
.A(n_6447),
.B(n_564),
.Y(n_6601)
);

OR2x2_ASAP7_75t_L g6602 ( 
.A(n_6414),
.B(n_565),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6402),
.Y(n_6603)
);

AND2x2_ASAP7_75t_L g6604 ( 
.A(n_6425),
.B(n_565),
.Y(n_6604)
);

OR2x2_ASAP7_75t_L g6605 ( 
.A(n_6387),
.B(n_566),
.Y(n_6605)
);

AND2x2_ASAP7_75t_L g6606 ( 
.A(n_6453),
.B(n_566),
.Y(n_6606)
);

NAND3xp33_ASAP7_75t_L g6607 ( 
.A(n_6389),
.B(n_567),
.C(n_568),
.Y(n_6607)
);

AOI221xp5_ASAP7_75t_L g6608 ( 
.A1(n_6486),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.C(n_570),
.Y(n_6608)
);

OA211x2_ASAP7_75t_L g6609 ( 
.A1(n_6419),
.A2(n_571),
.B(n_567),
.C(n_569),
.Y(n_6609)
);

INVx2_ASAP7_75t_SL g6610 ( 
.A(n_6441),
.Y(n_6610)
);

OAI21xp33_ASAP7_75t_SL g6611 ( 
.A1(n_6490),
.A2(n_6438),
.B(n_6437),
.Y(n_6611)
);

AO21x2_ASAP7_75t_L g6612 ( 
.A1(n_6458),
.A2(n_571),
.B(n_572),
.Y(n_6612)
);

OAI211xp5_ASAP7_75t_SL g6613 ( 
.A1(n_6393),
.A2(n_573),
.B(n_571),
.C(n_572),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6449),
.Y(n_6614)
);

NOR2xp33_ASAP7_75t_L g6615 ( 
.A(n_6405),
.B(n_572),
.Y(n_6615)
);

NAND3xp33_ASAP7_75t_L g6616 ( 
.A(n_6432),
.B(n_6567),
.C(n_6442),
.Y(n_6616)
);

NAND2xp5_ASAP7_75t_L g6617 ( 
.A(n_6499),
.B(n_573),
.Y(n_6617)
);

NAND3xp33_ASAP7_75t_SL g6618 ( 
.A(n_6481),
.B(n_573),
.C(n_574),
.Y(n_6618)
);

NOR3xp33_ASAP7_75t_L g6619 ( 
.A(n_6404),
.B(n_577),
.C(n_576),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_L g6620 ( 
.A(n_6478),
.B(n_575),
.Y(n_6620)
);

OR2x2_ASAP7_75t_L g6621 ( 
.A(n_6462),
.B(n_575),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6416),
.B(n_576),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_6479),
.Y(n_6623)
);

OA21x2_ASAP7_75t_L g6624 ( 
.A1(n_6474),
.A2(n_576),
.B(n_577),
.Y(n_6624)
);

OR2x2_ASAP7_75t_L g6625 ( 
.A(n_6519),
.B(n_577),
.Y(n_6625)
);

AOI22xp33_ASAP7_75t_L g6626 ( 
.A1(n_6473),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6448),
.Y(n_6627)
);

NAND3xp33_ASAP7_75t_L g6628 ( 
.A(n_6459),
.B(n_578),
.C(n_579),
.Y(n_6628)
);

INVxp67_ASAP7_75t_SL g6629 ( 
.A(n_6520),
.Y(n_6629)
);

XNOR2xp5_ASAP7_75t_L g6630 ( 
.A(n_6426),
.B(n_578),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6416),
.B(n_579),
.Y(n_6631)
);

INVx1_ASAP7_75t_L g6632 ( 
.A(n_6435),
.Y(n_6632)
);

AOI22x1_ASAP7_75t_L g6633 ( 
.A1(n_6524),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_6633)
);

AO21x2_ASAP7_75t_L g6634 ( 
.A1(n_6460),
.A2(n_580),
.B(n_581),
.Y(n_6634)
);

NOR2xp33_ASAP7_75t_L g6635 ( 
.A(n_6484),
.B(n_582),
.Y(n_6635)
);

AOI211xp5_ASAP7_75t_L g6636 ( 
.A1(n_6562),
.A2(n_585),
.B(n_583),
.C(n_584),
.Y(n_6636)
);

OR2x2_ASAP7_75t_L g6637 ( 
.A(n_6521),
.B(n_583),
.Y(n_6637)
);

AOI22xp33_ASAP7_75t_SL g6638 ( 
.A1(n_6430),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.Y(n_6638)
);

NOR3xp33_ASAP7_75t_L g6639 ( 
.A(n_6476),
.B(n_587),
.C(n_586),
.Y(n_6639)
);

AND2x2_ASAP7_75t_L g6640 ( 
.A(n_6529),
.B(n_585),
.Y(n_6640)
);

AND2x2_ASAP7_75t_L g6641 ( 
.A(n_6431),
.B(n_587),
.Y(n_6641)
);

NAND2xp5_ASAP7_75t_L g6642 ( 
.A(n_6497),
.B(n_587),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6436),
.Y(n_6643)
);

NAND2xp5_ASAP7_75t_L g6644 ( 
.A(n_6556),
.B(n_588),
.Y(n_6644)
);

INVx2_ASAP7_75t_L g6645 ( 
.A(n_6467),
.Y(n_6645)
);

OR2x2_ASAP7_75t_L g6646 ( 
.A(n_6386),
.B(n_588),
.Y(n_6646)
);

NOR2xp33_ASAP7_75t_L g6647 ( 
.A(n_6428),
.B(n_588),
.Y(n_6647)
);

INVxp67_ASAP7_75t_SL g6648 ( 
.A(n_6472),
.Y(n_6648)
);

AOI22xp33_ASAP7_75t_L g6649 ( 
.A1(n_6417),
.A2(n_592),
.B1(n_589),
.B2(n_591),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_6493),
.B(n_589),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_6396),
.B(n_589),
.Y(n_6651)
);

NAND3xp33_ASAP7_75t_L g6652 ( 
.A(n_6468),
.B(n_591),
.C(n_592),
.Y(n_6652)
);

OR2x2_ASAP7_75t_L g6653 ( 
.A(n_6560),
.B(n_591),
.Y(n_6653)
);

AND2x2_ASAP7_75t_L g6654 ( 
.A(n_6397),
.B(n_592),
.Y(n_6654)
);

OAI211xp5_ASAP7_75t_SL g6655 ( 
.A1(n_6512),
.A2(n_595),
.B(n_593),
.C(n_594),
.Y(n_6655)
);

NAND4xp25_ASAP7_75t_L g6656 ( 
.A(n_6535),
.B(n_595),
.C(n_593),
.D(n_594),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_6466),
.B(n_593),
.Y(n_6657)
);

NOR2xp33_ASAP7_75t_L g6658 ( 
.A(n_6428),
.B(n_594),
.Y(n_6658)
);

OAI21xp33_ASAP7_75t_SL g6659 ( 
.A1(n_6445),
.A2(n_595),
.B(n_596),
.Y(n_6659)
);

AO21x2_ASAP7_75t_L g6660 ( 
.A1(n_6394),
.A2(n_596),
.B(n_597),
.Y(n_6660)
);

NAND2xp5_ASAP7_75t_L g6661 ( 
.A(n_6469),
.B(n_596),
.Y(n_6661)
);

AND2x2_ASAP7_75t_L g6662 ( 
.A(n_6411),
.B(n_597),
.Y(n_6662)
);

AO21x2_ASAP7_75t_L g6663 ( 
.A1(n_6398),
.A2(n_598),
.B(n_599),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6444),
.Y(n_6664)
);

AND2x2_ASAP7_75t_L g6665 ( 
.A(n_6475),
.B(n_598),
.Y(n_6665)
);

NOR3xp33_ASAP7_75t_L g6666 ( 
.A(n_6545),
.B(n_599),
.C(n_600),
.Y(n_6666)
);

NAND3xp33_ASAP7_75t_L g6667 ( 
.A(n_6427),
.B(n_599),
.C(n_600),
.Y(n_6667)
);

NAND2xp5_ASAP7_75t_L g6668 ( 
.A(n_6533),
.B(n_601),
.Y(n_6668)
);

NAND3xp33_ASAP7_75t_L g6669 ( 
.A(n_6434),
.B(n_602),
.C(n_603),
.Y(n_6669)
);

NAND3xp33_ASAP7_75t_L g6670 ( 
.A(n_6485),
.B(n_602),
.C(n_603),
.Y(n_6670)
);

OR2x2_ASAP7_75t_L g6671 ( 
.A(n_6492),
.B(n_602),
.Y(n_6671)
);

AND2x2_ASAP7_75t_L g6672 ( 
.A(n_6532),
.B(n_6542),
.Y(n_6672)
);

AND2x2_ASAP7_75t_L g6673 ( 
.A(n_6457),
.B(n_604),
.Y(n_6673)
);

AND2x2_ASAP7_75t_L g6674 ( 
.A(n_6407),
.B(n_604),
.Y(n_6674)
);

NAND2xp5_ASAP7_75t_L g6675 ( 
.A(n_6522),
.B(n_605),
.Y(n_6675)
);

NAND2xp5_ASAP7_75t_SL g6676 ( 
.A(n_6400),
.B(n_605),
.Y(n_6676)
);

NOR2x1_ASAP7_75t_L g6677 ( 
.A(n_6495),
.B(n_605),
.Y(n_6677)
);

AOI22xp33_ASAP7_75t_L g6678 ( 
.A1(n_6417),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.Y(n_6678)
);

AO21x2_ASAP7_75t_L g6679 ( 
.A1(n_6571),
.A2(n_606),
.B(n_607),
.Y(n_6679)
);

NOR2xp33_ASAP7_75t_L g6680 ( 
.A(n_6525),
.B(n_607),
.Y(n_6680)
);

NAND3xp33_ASAP7_75t_SL g6681 ( 
.A(n_6513),
.B(n_608),
.C(n_609),
.Y(n_6681)
);

AND2x2_ASAP7_75t_L g6682 ( 
.A(n_6412),
.B(n_608),
.Y(n_6682)
);

NAND3xp33_ASAP7_75t_L g6683 ( 
.A(n_6487),
.B(n_609),
.C(n_610),
.Y(n_6683)
);

NAND2xp33_ASAP7_75t_SL g6684 ( 
.A(n_6538),
.B(n_609),
.Y(n_6684)
);

BUFx3_ASAP7_75t_L g6685 ( 
.A(n_6496),
.Y(n_6685)
);

NAND4xp75_ASAP7_75t_L g6686 ( 
.A(n_6465),
.B(n_612),
.C(n_610),
.D(n_611),
.Y(n_6686)
);

NAND3xp33_ASAP7_75t_L g6687 ( 
.A(n_6504),
.B(n_610),
.C(n_611),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_L g6688 ( 
.A(n_6456),
.B(n_611),
.Y(n_6688)
);

AOI221xp5_ASAP7_75t_L g6689 ( 
.A1(n_6403),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.C(n_615),
.Y(n_6689)
);

OR2x2_ASAP7_75t_L g6690 ( 
.A(n_6502),
.B(n_613),
.Y(n_6690)
);

NOR2xp33_ASAP7_75t_L g6691 ( 
.A(n_6441),
.B(n_614),
.Y(n_6691)
);

NAND3xp33_ASAP7_75t_L g6692 ( 
.A(n_6510),
.B(n_616),
.C(n_617),
.Y(n_6692)
);

NAND3xp33_ASAP7_75t_L g6693 ( 
.A(n_6511),
.B(n_616),
.C(n_617),
.Y(n_6693)
);

NAND3xp33_ASAP7_75t_L g6694 ( 
.A(n_6423),
.B(n_616),
.C(n_618),
.Y(n_6694)
);

NAND2xp5_ASAP7_75t_SL g6695 ( 
.A(n_6515),
.B(n_618),
.Y(n_6695)
);

AOI22xp33_ASAP7_75t_L g6696 ( 
.A1(n_6451),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.Y(n_6696)
);

OR2x2_ASAP7_75t_L g6697 ( 
.A(n_6531),
.B(n_6446),
.Y(n_6697)
);

AND2x2_ASAP7_75t_L g6698 ( 
.A(n_6415),
.B(n_619),
.Y(n_6698)
);

NAND2xp5_ASAP7_75t_L g6699 ( 
.A(n_6568),
.B(n_619),
.Y(n_6699)
);

NAND4xp25_ASAP7_75t_L g6700 ( 
.A(n_6443),
.B(n_622),
.C(n_620),
.D(n_621),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6506),
.Y(n_6701)
);

OR2x2_ASAP7_75t_L g6702 ( 
.A(n_6461),
.B(n_620),
.Y(n_6702)
);

INVx1_ASAP7_75t_SL g6703 ( 
.A(n_6539),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_SL g6704 ( 
.A(n_6399),
.B(n_621),
.Y(n_6704)
);

NAND4xp75_ASAP7_75t_L g6705 ( 
.A(n_6470),
.B(n_623),
.C(n_621),
.D(n_622),
.Y(n_6705)
);

NAND2xp5_ASAP7_75t_L g6706 ( 
.A(n_6401),
.B(n_622),
.Y(n_6706)
);

AOI22xp5_ASAP7_75t_L g6707 ( 
.A1(n_6452),
.A2(n_6408),
.B1(n_6424),
.B2(n_6421),
.Y(n_6707)
);

NAND3xp33_ASAP7_75t_L g6708 ( 
.A(n_6480),
.B(n_623),
.C(n_624),
.Y(n_6708)
);

AND2x2_ASAP7_75t_L g6709 ( 
.A(n_6516),
.B(n_623),
.Y(n_6709)
);

NAND2xp5_ASAP7_75t_SL g6710 ( 
.A(n_6537),
.B(n_624),
.Y(n_6710)
);

INVx2_ASAP7_75t_L g6711 ( 
.A(n_6503),
.Y(n_6711)
);

NOR2xp33_ASAP7_75t_L g6712 ( 
.A(n_6471),
.B(n_625),
.Y(n_6712)
);

OR2x2_ASAP7_75t_L g6713 ( 
.A(n_6541),
.B(n_625),
.Y(n_6713)
);

AOI22xp33_ASAP7_75t_SL g6714 ( 
.A1(n_6534),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_6714)
);

NOR2x1_ASAP7_75t_L g6715 ( 
.A(n_6559),
.B(n_626),
.Y(n_6715)
);

AOI211xp5_ASAP7_75t_L g6716 ( 
.A1(n_6463),
.A2(n_629),
.B(n_627),
.C(n_628),
.Y(n_6716)
);

NAND2xp5_ASAP7_75t_L g6717 ( 
.A(n_6454),
.B(n_627),
.Y(n_6717)
);

CKINVDCx5p33_ASAP7_75t_R g6718 ( 
.A(n_6516),
.Y(n_6718)
);

AOI22xp33_ASAP7_75t_L g6719 ( 
.A1(n_6477),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6413),
.Y(n_6720)
);

AND2x2_ASAP7_75t_SL g6721 ( 
.A(n_6392),
.B(n_6410),
.Y(n_6721)
);

NAND3xp33_ASAP7_75t_L g6722 ( 
.A(n_6505),
.B(n_630),
.C(n_631),
.Y(n_6722)
);

AND2x2_ASAP7_75t_L g6723 ( 
.A(n_6483),
.B(n_631),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6488),
.Y(n_6724)
);

NAND3xp33_ASAP7_75t_L g6725 ( 
.A(n_6527),
.B(n_632),
.C(n_633),
.Y(n_6725)
);

AND2x2_ASAP7_75t_L g6726 ( 
.A(n_6518),
.B(n_632),
.Y(n_6726)
);

AND2x2_ASAP7_75t_SL g6727 ( 
.A(n_6523),
.B(n_6530),
.Y(n_6727)
);

NAND3xp33_ASAP7_75t_L g6728 ( 
.A(n_6553),
.B(n_633),
.C(n_634),
.Y(n_6728)
);

NAND3xp33_ASAP7_75t_L g6729 ( 
.A(n_6557),
.B(n_633),
.C(n_634),
.Y(n_6729)
);

AO21x2_ASAP7_75t_L g6730 ( 
.A1(n_6517),
.A2(n_634),
.B(n_635),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_6509),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6433),
.Y(n_6732)
);

AND2x2_ASAP7_75t_L g6733 ( 
.A(n_6585),
.B(n_6526),
.Y(n_6733)
);

INVx1_ASAP7_75t_SL g6734 ( 
.A(n_6576),
.Y(n_6734)
);

NAND3xp33_ASAP7_75t_L g6735 ( 
.A(n_6598),
.B(n_6508),
.C(n_6536),
.Y(n_6735)
);

INVx2_ASAP7_75t_L g6736 ( 
.A(n_6574),
.Y(n_6736)
);

OAI221xp5_ASAP7_75t_SL g6737 ( 
.A1(n_6580),
.A2(n_6528),
.B1(n_6543),
.B2(n_6406),
.C(n_6501),
.Y(n_6737)
);

NAND4xp75_ASAP7_75t_L g6738 ( 
.A(n_6610),
.B(n_6464),
.C(n_6500),
.D(n_6547),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_6578),
.Y(n_6739)
);

NAND2xp5_ASAP7_75t_L g6740 ( 
.A(n_6577),
.B(n_6540),
.Y(n_6740)
);

NAND2xp5_ASAP7_75t_L g6741 ( 
.A(n_6622),
.B(n_6503),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6595),
.B(n_6593),
.Y(n_6742)
);

OAI211xp5_ASAP7_75t_L g6743 ( 
.A1(n_6611),
.A2(n_6514),
.B(n_6498),
.C(n_6491),
.Y(n_6743)
);

INVx2_ASAP7_75t_L g6744 ( 
.A(n_6685),
.Y(n_6744)
);

INVxp67_ASAP7_75t_L g6745 ( 
.A(n_6631),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6604),
.Y(n_6746)
);

NAND2xp5_ASAP7_75t_SL g6747 ( 
.A(n_6721),
.B(n_6544),
.Y(n_6747)
);

INVxp67_ASAP7_75t_L g6748 ( 
.A(n_6606),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6720),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_6588),
.B(n_6546),
.Y(n_6750)
);

BUFx3_ASAP7_75t_L g6751 ( 
.A(n_6582),
.Y(n_6751)
);

AOI221xp5_ASAP7_75t_SL g6752 ( 
.A1(n_6575),
.A2(n_6420),
.B1(n_6507),
.B2(n_6494),
.C(n_6482),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6620),
.Y(n_6753)
);

NAND2xp5_ASAP7_75t_L g6754 ( 
.A(n_6582),
.B(n_6548),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_6645),
.Y(n_6755)
);

AND2x4_ASAP7_75t_L g6756 ( 
.A(n_6614),
.B(n_6558),
.Y(n_6756)
);

HB1xp67_ASAP7_75t_L g6757 ( 
.A(n_6623),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6709),
.Y(n_6758)
);

NOR3xp33_ASAP7_75t_L g6759 ( 
.A(n_6681),
.B(n_636),
.C(n_637),
.Y(n_6759)
);

NAND2xp5_ASAP7_75t_L g6760 ( 
.A(n_6673),
.B(n_636),
.Y(n_6760)
);

AOI211xp5_ASAP7_75t_L g6761 ( 
.A1(n_6616),
.A2(n_638),
.B(n_636),
.C(n_637),
.Y(n_6761)
);

INVx1_ASAP7_75t_L g6762 ( 
.A(n_6642),
.Y(n_6762)
);

AND2x2_ASAP7_75t_L g6763 ( 
.A(n_6589),
.B(n_6662),
.Y(n_6763)
);

XNOR2xp5_ASAP7_75t_L g6764 ( 
.A(n_6630),
.B(n_637),
.Y(n_6764)
);

HB1xp67_ASAP7_75t_L g6765 ( 
.A(n_6664),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6665),
.Y(n_6766)
);

NOR2xp33_ASAP7_75t_L g6767 ( 
.A(n_6659),
.B(n_638),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6701),
.Y(n_6768)
);

NAND2xp5_ASAP7_75t_L g6769 ( 
.A(n_6639),
.B(n_638),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6641),
.B(n_639),
.Y(n_6770)
);

AOI22xp33_ASAP7_75t_L g6771 ( 
.A1(n_6619),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.Y(n_6771)
);

INVx1_ASAP7_75t_L g6772 ( 
.A(n_6651),
.Y(n_6772)
);

CKINVDCx5p33_ASAP7_75t_R g6773 ( 
.A(n_6718),
.Y(n_6773)
);

AOI222xp33_ASAP7_75t_L g6774 ( 
.A1(n_6603),
.A2(n_642),
.B1(n_644),
.B2(n_640),
.C1(n_641),
.C2(n_643),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6654),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6602),
.Y(n_6776)
);

INVx1_ASAP7_75t_SL g6777 ( 
.A(n_6592),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6691),
.Y(n_6778)
);

AND2x2_ASAP7_75t_L g6779 ( 
.A(n_6672),
.B(n_640),
.Y(n_6779)
);

AOI33xp33_ASAP7_75t_L g6780 ( 
.A1(n_6632),
.A2(n_643),
.A3(n_645),
.B1(n_641),
.B2(n_642),
.B3(n_644),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6723),
.B(n_643),
.Y(n_6781)
);

AND2x2_ASAP7_75t_L g6782 ( 
.A(n_6726),
.B(n_644),
.Y(n_6782)
);

AO22x1_ASAP7_75t_L g6783 ( 
.A1(n_6596),
.A2(n_647),
.B1(n_645),
.B2(n_646),
.Y(n_6783)
);

OR2x2_ASAP7_75t_L g6784 ( 
.A(n_6600),
.B(n_6583),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6599),
.Y(n_6785)
);

OAI22xp5_ASAP7_75t_SL g6786 ( 
.A1(n_6711),
.A2(n_647),
.B1(n_645),
.B2(n_646),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_6601),
.Y(n_6787)
);

INVx1_ASAP7_75t_L g6788 ( 
.A(n_6624),
.Y(n_6788)
);

NAND2xp5_ASAP7_75t_L g6789 ( 
.A(n_6638),
.B(n_647),
.Y(n_6789)
);

AND2x2_ASAP7_75t_L g6790 ( 
.A(n_6682),
.B(n_648),
.Y(n_6790)
);

AND2x4_ASAP7_75t_L g6791 ( 
.A(n_6643),
.B(n_648),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6698),
.B(n_649),
.Y(n_6792)
);

AND2x2_ASAP7_75t_L g6793 ( 
.A(n_6674),
.B(n_6703),
.Y(n_6793)
);

AND2x2_ASAP7_75t_L g6794 ( 
.A(n_6629),
.B(n_649),
.Y(n_6794)
);

OAI33xp33_ASAP7_75t_L g6795 ( 
.A1(n_6627),
.A2(n_651),
.A3(n_653),
.B1(n_649),
.B2(n_650),
.B3(n_652),
.Y(n_6795)
);

INVxp67_ASAP7_75t_L g6796 ( 
.A(n_6684),
.Y(n_6796)
);

CKINVDCx16_ASAP7_75t_R g6797 ( 
.A(n_6625),
.Y(n_6797)
);

INVxp67_ASAP7_75t_L g6798 ( 
.A(n_6635),
.Y(n_6798)
);

AND2x6_ASAP7_75t_L g6799 ( 
.A(n_6647),
.B(n_650),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6624),
.Y(n_6800)
);

OR2x2_ASAP7_75t_L g6801 ( 
.A(n_6644),
.B(n_651),
.Y(n_6801)
);

AOI22xp33_ASAP7_75t_SL g6802 ( 
.A1(n_6727),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_6802)
);

OAI211xp5_ASAP7_75t_L g6803 ( 
.A1(n_6707),
.A2(n_656),
.B(n_654),
.C(n_655),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6594),
.Y(n_6804)
);

INVx2_ASAP7_75t_L g6805 ( 
.A(n_6671),
.Y(n_6805)
);

AOI22xp33_ASAP7_75t_L g6806 ( 
.A1(n_6572),
.A2(n_6573),
.B1(n_6731),
.B2(n_6724),
.Y(n_6806)
);

NAND2xp5_ASAP7_75t_L g6807 ( 
.A(n_6636),
.B(n_654),
.Y(n_6807)
);

INVx3_ASAP7_75t_L g6808 ( 
.A(n_6690),
.Y(n_6808)
);

NAND2xp5_ASAP7_75t_L g6809 ( 
.A(n_6584),
.B(n_655),
.Y(n_6809)
);

AND2x2_ASAP7_75t_L g6810 ( 
.A(n_6615),
.B(n_655),
.Y(n_6810)
);

NAND2xp5_ASAP7_75t_L g6811 ( 
.A(n_6663),
.B(n_657),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6633),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6633),
.Y(n_6813)
);

INVx2_ASAP7_75t_L g6814 ( 
.A(n_6730),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6686),
.Y(n_6815)
);

AOI221xp5_ASAP7_75t_L g6816 ( 
.A1(n_6648),
.A2(n_659),
.B1(n_657),
.B2(n_658),
.C(n_660),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6649),
.B(n_657),
.Y(n_6817)
);

OR2x2_ASAP7_75t_L g6818 ( 
.A(n_6702),
.B(n_658),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6640),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6675),
.Y(n_6820)
);

AOI22xp33_ASAP7_75t_L g6821 ( 
.A1(n_6732),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.Y(n_6821)
);

INVx2_ASAP7_75t_L g6822 ( 
.A(n_6705),
.Y(n_6822)
);

NAND2xp5_ASAP7_75t_L g6823 ( 
.A(n_6678),
.B(n_661),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_6688),
.Y(n_6824)
);

NAND2xp5_ASAP7_75t_L g6825 ( 
.A(n_6714),
.B(n_663),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_6650),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_6679),
.B(n_663),
.Y(n_6827)
);

INVx1_ASAP7_75t_L g6828 ( 
.A(n_6657),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6590),
.B(n_664),
.Y(n_6829)
);

CKINVDCx16_ASAP7_75t_R g6830 ( 
.A(n_6618),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6661),
.Y(n_6831)
);

OAI211xp5_ASAP7_75t_L g6832 ( 
.A1(n_6656),
.A2(n_666),
.B(n_664),
.C(n_665),
.Y(n_6832)
);

HB1xp67_ASAP7_75t_L g6833 ( 
.A(n_6658),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6712),
.B(n_664),
.Y(n_6834)
);

AND2x4_ASAP7_75t_L g6835 ( 
.A(n_6628),
.B(n_665),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6660),
.Y(n_6836)
);

OR2x2_ASAP7_75t_L g6837 ( 
.A(n_6621),
.B(n_666),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6677),
.Y(n_6838)
);

AOI221x1_ASAP7_75t_L g6839 ( 
.A1(n_6680),
.A2(n_669),
.B1(n_667),
.B2(n_668),
.C(n_670),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_6668),
.Y(n_6840)
);

INVx2_ASAP7_75t_L g6841 ( 
.A(n_6637),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6697),
.B(n_667),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6713),
.B(n_667),
.Y(n_6843)
);

INVx4_ASAP7_75t_L g6844 ( 
.A(n_6605),
.Y(n_6844)
);

AND2x2_ASAP7_75t_SL g6845 ( 
.A(n_6666),
.B(n_668),
.Y(n_6845)
);

AOI21xp5_ASAP7_75t_SL g6846 ( 
.A1(n_6612),
.A2(n_6634),
.B(n_6676),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6617),
.Y(n_6847)
);

AND2x2_ASAP7_75t_L g6848 ( 
.A(n_6646),
.B(n_6653),
.Y(n_6848)
);

OAI221xp5_ASAP7_75t_L g6849 ( 
.A1(n_6607),
.A2(n_671),
.B1(n_668),
.B2(n_669),
.C(n_672),
.Y(n_6849)
);

AOI33xp33_ASAP7_75t_L g6850 ( 
.A1(n_6719),
.A2(n_672),
.A3(n_674),
.B1(n_669),
.B2(n_671),
.B3(n_673),
.Y(n_6850)
);

AND2x4_ASAP7_75t_L g6851 ( 
.A(n_6652),
.B(n_671),
.Y(n_6851)
);

OR2x2_ASAP7_75t_L g6852 ( 
.A(n_6700),
.B(n_672),
.Y(n_6852)
);

HB1xp67_ASAP7_75t_L g6853 ( 
.A(n_6591),
.Y(n_6853)
);

AOI21xp5_ASAP7_75t_L g6854 ( 
.A1(n_6695),
.A2(n_673),
.B(n_674),
.Y(n_6854)
);

NAND2xp5_ASAP7_75t_L g6855 ( 
.A(n_6626),
.B(n_675),
.Y(n_6855)
);

AOI221xp5_ASAP7_75t_L g6856 ( 
.A1(n_6655),
.A2(n_677),
.B1(n_675),
.B2(n_676),
.C(n_678),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_6579),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6689),
.B(n_675),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_L g6859 ( 
.A(n_6608),
.B(n_676),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_6581),
.Y(n_6860)
);

AOI31xp33_ASAP7_75t_L g6861 ( 
.A1(n_6715),
.A2(n_678),
.A3(n_676),
.B(n_677),
.Y(n_6861)
);

AND2x2_ASAP7_75t_L g6862 ( 
.A(n_6717),
.B(n_678),
.Y(n_6862)
);

AOI22xp33_ASAP7_75t_L g6863 ( 
.A1(n_6609),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_6863)
);

AND2x4_ASAP7_75t_L g6864 ( 
.A(n_6587),
.B(n_679),
.Y(n_6864)
);

INVx2_ASAP7_75t_L g6865 ( 
.A(n_6586),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6670),
.Y(n_6866)
);

INVx2_ASAP7_75t_L g6867 ( 
.A(n_6597),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6683),
.Y(n_6868)
);

INVx3_ASAP7_75t_L g6869 ( 
.A(n_6706),
.Y(n_6869)
);

OR2x2_ASAP7_75t_L g6870 ( 
.A(n_6699),
.B(n_679),
.Y(n_6870)
);

INVx2_ASAP7_75t_SL g6871 ( 
.A(n_6710),
.Y(n_6871)
);

AOI22xp33_ASAP7_75t_SL g6872 ( 
.A1(n_6694),
.A2(n_682),
.B1(n_680),
.B2(n_681),
.Y(n_6872)
);

AND2x4_ASAP7_75t_L g6873 ( 
.A(n_6687),
.B(n_6692),
.Y(n_6873)
);

OR2x2_ASAP7_75t_L g6874 ( 
.A(n_6667),
.B(n_680),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6693),
.Y(n_6875)
);

HB1xp67_ASAP7_75t_L g6876 ( 
.A(n_6704),
.Y(n_6876)
);

OAI21xp5_ASAP7_75t_L g6877 ( 
.A1(n_6669),
.A2(n_682),
.B(n_683),
.Y(n_6877)
);

AOI221xp5_ASAP7_75t_L g6878 ( 
.A1(n_6725),
.A2(n_684),
.B1(n_682),
.B2(n_683),
.C(n_685),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6708),
.Y(n_6879)
);

OAI221xp5_ASAP7_75t_L g6880 ( 
.A1(n_6728),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.C(n_686),
.Y(n_6880)
);

AND2x2_ASAP7_75t_L g6881 ( 
.A(n_6696),
.B(n_684),
.Y(n_6881)
);

NAND3xp33_ASAP7_75t_L g6882 ( 
.A(n_6716),
.B(n_685),
.C(n_687),
.Y(n_6882)
);

NOR2xp33_ASAP7_75t_L g6883 ( 
.A(n_6722),
.B(n_687),
.Y(n_6883)
);

OAI33xp33_ASAP7_75t_L g6884 ( 
.A1(n_6729),
.A2(n_689),
.A3(n_691),
.B1(n_687),
.B2(n_688),
.B3(n_690),
.Y(n_6884)
);

AOI221xp5_ASAP7_75t_L g6885 ( 
.A1(n_6613),
.A2(n_690),
.B1(n_688),
.B2(n_689),
.C(n_691),
.Y(n_6885)
);

AOI31xp33_ASAP7_75t_L g6886 ( 
.A1(n_6580),
.A2(n_690),
.A3(n_688),
.B(n_689),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6580),
.Y(n_6887)
);

INVx2_ASAP7_75t_L g6888 ( 
.A(n_6574),
.Y(n_6888)
);

BUFx2_ASAP7_75t_L g6889 ( 
.A(n_6580),
.Y(n_6889)
);

AND2x2_ASAP7_75t_L g6890 ( 
.A(n_6585),
.B(n_691),
.Y(n_6890)
);

OAI31xp33_ASAP7_75t_L g6891 ( 
.A1(n_6616),
.A2(n_694),
.A3(n_692),
.B(n_693),
.Y(n_6891)
);

AND2x2_ASAP7_75t_L g6892 ( 
.A(n_6585),
.B(n_692),
.Y(n_6892)
);

INVx1_ASAP7_75t_L g6893 ( 
.A(n_6580),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6889),
.Y(n_6894)
);

OR2x2_ASAP7_75t_L g6895 ( 
.A(n_6744),
.B(n_692),
.Y(n_6895)
);

INVx2_ASAP7_75t_L g6896 ( 
.A(n_6751),
.Y(n_6896)
);

AND2x2_ASAP7_75t_L g6897 ( 
.A(n_6742),
.B(n_693),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6749),
.Y(n_6898)
);

AND2x2_ASAP7_75t_L g6899 ( 
.A(n_6779),
.B(n_694),
.Y(n_6899)
);

OR2x2_ASAP7_75t_L g6900 ( 
.A(n_6736),
.B(n_695),
.Y(n_6900)
);

INVx1_ASAP7_75t_L g6901 ( 
.A(n_6788),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_6890),
.B(n_695),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6800),
.Y(n_6903)
);

INVx1_ASAP7_75t_L g6904 ( 
.A(n_6765),
.Y(n_6904)
);

AND2x2_ASAP7_75t_L g6905 ( 
.A(n_6892),
.B(n_695),
.Y(n_6905)
);

NAND2x1p5_ASAP7_75t_L g6906 ( 
.A(n_6888),
.B(n_696),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6755),
.Y(n_6907)
);

AND2x2_ASAP7_75t_L g6908 ( 
.A(n_6790),
.B(n_697),
.Y(n_6908)
);

INVx1_ASAP7_75t_L g6909 ( 
.A(n_6770),
.Y(n_6909)
);

OR2x2_ASAP7_75t_L g6910 ( 
.A(n_6887),
.B(n_697),
.Y(n_6910)
);

OAI21xp33_ASAP7_75t_L g6911 ( 
.A1(n_6743),
.A2(n_6773),
.B(n_6767),
.Y(n_6911)
);

NAND3xp33_ASAP7_75t_L g6912 ( 
.A(n_6761),
.B(n_697),
.C(n_698),
.Y(n_6912)
);

INVx2_ASAP7_75t_SL g6913 ( 
.A(n_6768),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6893),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6786),
.Y(n_6915)
);

INVxp67_ASAP7_75t_L g6916 ( 
.A(n_6781),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_6792),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6757),
.Y(n_6918)
);

BUFx2_ASAP7_75t_L g6919 ( 
.A(n_6791),
.Y(n_6919)
);

AND2x2_ASAP7_75t_L g6920 ( 
.A(n_6763),
.B(n_698),
.Y(n_6920)
);

INVx1_ASAP7_75t_SL g6921 ( 
.A(n_6734),
.Y(n_6921)
);

NAND2x1_ASAP7_75t_L g6922 ( 
.A(n_6756),
.B(n_699),
.Y(n_6922)
);

OR2x2_ASAP7_75t_L g6923 ( 
.A(n_6852),
.B(n_699),
.Y(n_6923)
);

AOI22xp5_ASAP7_75t_L g6924 ( 
.A1(n_6830),
.A2(n_6759),
.B1(n_6832),
.B2(n_6796),
.Y(n_6924)
);

OR2x2_ASAP7_75t_L g6925 ( 
.A(n_6812),
.B(n_699),
.Y(n_6925)
);

NOR4xp25_ASAP7_75t_SL g6926 ( 
.A(n_6737),
.B(n_702),
.C(n_700),
.D(n_701),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6791),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6874),
.Y(n_6928)
);

NAND2x1p5_ASAP7_75t_L g6929 ( 
.A(n_6860),
.B(n_700),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6794),
.B(n_700),
.Y(n_6930)
);

NAND2xp5_ASAP7_75t_L g6931 ( 
.A(n_6783),
.B(n_701),
.Y(n_6931)
);

INVx2_ASAP7_75t_SL g6932 ( 
.A(n_6864),
.Y(n_6932)
);

INVxp67_ASAP7_75t_L g6933 ( 
.A(n_6782),
.Y(n_6933)
);

AND2x2_ASAP7_75t_L g6934 ( 
.A(n_6842),
.B(n_701),
.Y(n_6934)
);

OR2x2_ASAP7_75t_L g6935 ( 
.A(n_6813),
.B(n_702),
.Y(n_6935)
);

OR2x2_ASAP7_75t_L g6936 ( 
.A(n_6811),
.B(n_6809),
.Y(n_6936)
);

NAND2xp5_ASAP7_75t_L g6937 ( 
.A(n_6863),
.B(n_702),
.Y(n_6937)
);

AND2x2_ASAP7_75t_L g6938 ( 
.A(n_6793),
.B(n_703),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6862),
.Y(n_6939)
);

NAND2xp5_ASAP7_75t_L g6940 ( 
.A(n_6799),
.B(n_703),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_L g6941 ( 
.A(n_6799),
.B(n_703),
.Y(n_6941)
);

INVx1_ASAP7_75t_SL g6942 ( 
.A(n_6777),
.Y(n_6942)
);

O2A1O1Ixp5_ASAP7_75t_SL g6943 ( 
.A1(n_6747),
.A2(n_6838),
.B(n_6833),
.C(n_6778),
.Y(n_6943)
);

INVx1_ASAP7_75t_L g6944 ( 
.A(n_6810),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6733),
.B(n_704),
.Y(n_6945)
);

INVxp67_ASAP7_75t_SL g6946 ( 
.A(n_6760),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6801),
.Y(n_6947)
);

NOR2xp33_ASAP7_75t_L g6948 ( 
.A(n_6795),
.B(n_705),
.Y(n_6948)
);

NOR2xp67_ASAP7_75t_L g6949 ( 
.A(n_6745),
.B(n_705),
.Y(n_6949)
);

OR2x2_ASAP7_75t_L g6950 ( 
.A(n_6789),
.B(n_706),
.Y(n_6950)
);

AND2x2_ASAP7_75t_L g6951 ( 
.A(n_6829),
.B(n_706),
.Y(n_6951)
);

NAND2x1p5_ASAP7_75t_SL g6952 ( 
.A(n_6815),
.B(n_706),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_6843),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6780),
.Y(n_6954)
);

OR2x2_ASAP7_75t_L g6955 ( 
.A(n_6817),
.B(n_707),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6818),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6837),
.Y(n_6957)
);

NAND2xp5_ASAP7_75t_L g6958 ( 
.A(n_6799),
.B(n_707),
.Y(n_6958)
);

AND2x2_ASAP7_75t_L g6959 ( 
.A(n_6834),
.B(n_6750),
.Y(n_6959)
);

OR2x2_ASAP7_75t_L g6960 ( 
.A(n_6823),
.B(n_707),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_6756),
.Y(n_6961)
);

OR2x2_ASAP7_75t_L g6962 ( 
.A(n_6797),
.B(n_708),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_6835),
.Y(n_6963)
);

AO31x2_ASAP7_75t_L g6964 ( 
.A1(n_6836),
.A2(n_6844),
.A3(n_6758),
.B(n_6822),
.Y(n_6964)
);

INVx2_ASAP7_75t_L g6965 ( 
.A(n_6804),
.Y(n_6965)
);

AND2x2_ASAP7_75t_L g6966 ( 
.A(n_6881),
.B(n_6848),
.Y(n_6966)
);

AND2x2_ASAP7_75t_L g6967 ( 
.A(n_6845),
.B(n_6739),
.Y(n_6967)
);

INVx2_ASAP7_75t_SL g6968 ( 
.A(n_6805),
.Y(n_6968)
);

NOR2x1_ASAP7_75t_L g6969 ( 
.A(n_6846),
.B(n_708),
.Y(n_6969)
);

HB1xp67_ASAP7_75t_L g6970 ( 
.A(n_6766),
.Y(n_6970)
);

AND2x4_ASAP7_75t_L g6971 ( 
.A(n_6865),
.B(n_708),
.Y(n_6971)
);

NAND2xp5_ASAP7_75t_L g6972 ( 
.A(n_6802),
.B(n_709),
.Y(n_6972)
);

INVx2_ASAP7_75t_L g6973 ( 
.A(n_6808),
.Y(n_6973)
);

AND2x2_ASAP7_75t_L g6974 ( 
.A(n_6746),
.B(n_709),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6835),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6819),
.B(n_710),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6851),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6851),
.Y(n_6978)
);

NAND2xp5_ASAP7_75t_L g6979 ( 
.A(n_6891),
.B(n_710),
.Y(n_6979)
);

INVx2_ASAP7_75t_SL g6980 ( 
.A(n_6867),
.Y(n_6980)
);

INVx3_ASAP7_75t_L g6981 ( 
.A(n_6873),
.Y(n_6981)
);

INVx2_ASAP7_75t_L g6982 ( 
.A(n_6841),
.Y(n_6982)
);

INVx2_ASAP7_75t_SL g6983 ( 
.A(n_6741),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6886),
.Y(n_6984)
);

INVxp67_ASAP7_75t_L g6985 ( 
.A(n_6883),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6870),
.Y(n_6986)
);

INVxp67_ASAP7_75t_L g6987 ( 
.A(n_6827),
.Y(n_6987)
);

HB1xp67_ASAP7_75t_L g6988 ( 
.A(n_6876),
.Y(n_6988)
);

NOR2xp33_ASAP7_75t_L g6989 ( 
.A(n_6803),
.B(n_711),
.Y(n_6989)
);

AND2x2_ASAP7_75t_SL g6990 ( 
.A(n_6873),
.B(n_712),
.Y(n_6990)
);

AND2x2_ASAP7_75t_L g6991 ( 
.A(n_6748),
.B(n_712),
.Y(n_6991)
);

OR2x2_ASAP7_75t_L g6992 ( 
.A(n_6855),
.B(n_712),
.Y(n_6992)
);

NAND2x1p5_ASAP7_75t_L g6993 ( 
.A(n_6857),
.B(n_713),
.Y(n_6993)
);

NAND2xp67_ASAP7_75t_L g6994 ( 
.A(n_6814),
.B(n_713),
.Y(n_6994)
);

NOR2x1_ASAP7_75t_L g6995 ( 
.A(n_6735),
.B(n_713),
.Y(n_6995)
);

OR2x2_ASAP7_75t_L g6996 ( 
.A(n_6825),
.B(n_714),
.Y(n_6996)
);

INVx1_ASAP7_75t_L g6997 ( 
.A(n_6772),
.Y(n_6997)
);

INVx1_ASAP7_75t_SL g6998 ( 
.A(n_6754),
.Y(n_6998)
);

INVx1_ASAP7_75t_L g6999 ( 
.A(n_6775),
.Y(n_6999)
);

AND2x2_ASAP7_75t_L g7000 ( 
.A(n_6776),
.B(n_715),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6850),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6871),
.B(n_6879),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_L g7003 ( 
.A(n_6764),
.B(n_715),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6784),
.Y(n_7004)
);

AND2x4_ASAP7_75t_L g7005 ( 
.A(n_6877),
.B(n_715),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6866),
.B(n_716),
.Y(n_7006)
);

INVx2_ASAP7_75t_L g7007 ( 
.A(n_6738),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6807),
.Y(n_7008)
);

INVxp67_ASAP7_75t_L g7009 ( 
.A(n_6849),
.Y(n_7009)
);

OAI211xp5_ASAP7_75t_L g7010 ( 
.A1(n_6868),
.A2(n_718),
.B(n_716),
.C(n_717),
.Y(n_7010)
);

NAND2xp5_ASAP7_75t_L g7011 ( 
.A(n_6774),
.B(n_716),
.Y(n_7011)
);

NAND3xp33_ASAP7_75t_L g7012 ( 
.A(n_6816),
.B(n_6771),
.C(n_6839),
.Y(n_7012)
);

HB1xp67_ASAP7_75t_L g7013 ( 
.A(n_6875),
.Y(n_7013)
);

NAND2xp5_ASAP7_75t_L g7014 ( 
.A(n_6872),
.B(n_717),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6901),
.Y(n_7015)
);

INVx1_ASAP7_75t_L g7016 ( 
.A(n_6903),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6922),
.Y(n_7017)
);

HB1xp67_ASAP7_75t_L g7018 ( 
.A(n_6913),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6971),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6971),
.Y(n_7020)
);

OR2x2_ASAP7_75t_L g7021 ( 
.A(n_7007),
.B(n_6769),
.Y(n_7021)
);

OR4x1_ASAP7_75t_L g7022 ( 
.A(n_6980),
.B(n_6826),
.C(n_6831),
.D(n_6828),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6940),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6941),
.Y(n_7024)
);

INVxp67_ASAP7_75t_L g7025 ( 
.A(n_6897),
.Y(n_7025)
);

AND2x2_ASAP7_75t_L g7026 ( 
.A(n_6938),
.B(n_6798),
.Y(n_7026)
);

OAI32xp33_ASAP7_75t_L g7027 ( 
.A1(n_6998),
.A2(n_6740),
.A3(n_6840),
.B1(n_6753),
.B2(n_6824),
.Y(n_7027)
);

INVx2_ASAP7_75t_L g7028 ( 
.A(n_6896),
.Y(n_7028)
);

INVx2_ASAP7_75t_L g7029 ( 
.A(n_6907),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6958),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6906),
.Y(n_7031)
);

OAI22xp5_ASAP7_75t_L g7032 ( 
.A1(n_6924),
.A2(n_6806),
.B1(n_6858),
.B2(n_6882),
.Y(n_7032)
);

AND2x2_ASAP7_75t_L g7033 ( 
.A(n_6945),
.B(n_6853),
.Y(n_7033)
);

NAND2xp5_ASAP7_75t_L g7034 ( 
.A(n_6948),
.B(n_6861),
.Y(n_7034)
);

OR2x2_ASAP7_75t_L g7035 ( 
.A(n_6952),
.B(n_6859),
.Y(n_7035)
);

INVx1_ASAP7_75t_L g7036 ( 
.A(n_6925),
.Y(n_7036)
);

AOI21xp33_ASAP7_75t_L g7037 ( 
.A1(n_6911),
.A2(n_6954),
.B(n_6894),
.Y(n_7037)
);

INVx2_ASAP7_75t_SL g7038 ( 
.A(n_6961),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6899),
.B(n_6869),
.Y(n_7039)
);

INVx1_ASAP7_75t_L g7040 ( 
.A(n_6935),
.Y(n_7040)
);

NAND2xp5_ASAP7_75t_L g7041 ( 
.A(n_6930),
.B(n_6821),
.Y(n_7041)
);

HB1xp67_ASAP7_75t_L g7042 ( 
.A(n_6919),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6962),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6923),
.Y(n_7044)
);

NAND2xp5_ASAP7_75t_L g7045 ( 
.A(n_6920),
.B(n_6878),
.Y(n_7045)
);

INVx2_ASAP7_75t_SL g7046 ( 
.A(n_6965),
.Y(n_7046)
);

INVx1_ASAP7_75t_L g7047 ( 
.A(n_7006),
.Y(n_7047)
);

NAND2xp5_ASAP7_75t_L g7048 ( 
.A(n_6981),
.B(n_6752),
.Y(n_7048)
);

NOR2xp67_ASAP7_75t_L g7049 ( 
.A(n_6968),
.B(n_6932),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6895),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6910),
.Y(n_7051)
);

INVx1_ASAP7_75t_L g7052 ( 
.A(n_6931),
.Y(n_7052)
);

AND2x2_ASAP7_75t_L g7053 ( 
.A(n_6934),
.B(n_6847),
.Y(n_7053)
);

HB1xp67_ASAP7_75t_L g7054 ( 
.A(n_6993),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_6900),
.Y(n_7055)
);

NAND2x1p5_ASAP7_75t_L g7056 ( 
.A(n_6942),
.B(n_6785),
.Y(n_7056)
);

HB1xp67_ASAP7_75t_L g7057 ( 
.A(n_6963),
.Y(n_7057)
);

OAI322xp33_ASAP7_75t_L g7058 ( 
.A1(n_6921),
.A2(n_6820),
.A3(n_6787),
.B1(n_6762),
.B2(n_6880),
.C1(n_6854),
.C2(n_6884),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_7000),
.Y(n_7059)
);

OAI22xp33_ASAP7_75t_L g7060 ( 
.A1(n_6937),
.A2(n_6856),
.B1(n_6885),
.B2(n_720),
.Y(n_7060)
);

AOI33xp33_ASAP7_75t_L g7061 ( 
.A1(n_6926),
.A2(n_720),
.A3(n_722),
.B1(n_718),
.B2(n_719),
.B3(n_721),
.Y(n_7061)
);

INVx1_ASAP7_75t_SL g7062 ( 
.A(n_7002),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_L g7063 ( 
.A(n_6989),
.B(n_719),
.Y(n_7063)
);

INVx1_ASAP7_75t_L g7064 ( 
.A(n_6991),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6976),
.Y(n_7065)
);

AND2x2_ASAP7_75t_L g7066 ( 
.A(n_6902),
.B(n_719),
.Y(n_7066)
);

INVx2_ASAP7_75t_L g7067 ( 
.A(n_6982),
.Y(n_7067)
);

NAND2xp5_ASAP7_75t_L g7068 ( 
.A(n_6905),
.B(n_722),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6929),
.Y(n_7069)
);

INVx1_ASAP7_75t_SL g7070 ( 
.A(n_6927),
.Y(n_7070)
);

OAI22xp5_ASAP7_75t_L g7071 ( 
.A1(n_7009),
.A2(n_724),
.B1(n_722),
.B2(n_723),
.Y(n_7071)
);

AOI22xp33_ASAP7_75t_SL g7072 ( 
.A1(n_7001),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_7072)
);

A2O1A1Ixp33_ASAP7_75t_L g7073 ( 
.A1(n_6912),
.A2(n_726),
.B(n_723),
.C(n_725),
.Y(n_7073)
);

NAND2xp5_ASAP7_75t_L g7074 ( 
.A(n_6908),
.B(n_725),
.Y(n_7074)
);

NAND2xp5_ASAP7_75t_L g7075 ( 
.A(n_6984),
.B(n_726),
.Y(n_7075)
);

INVx1_ASAP7_75t_L g7076 ( 
.A(n_6988),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6974),
.Y(n_7077)
);

OAI22x1_ASAP7_75t_L g7078 ( 
.A1(n_7005),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_7078)
);

INVx2_ASAP7_75t_L g7079 ( 
.A(n_6973),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6994),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_6983),
.Y(n_7081)
);

INVx2_ASAP7_75t_SL g7082 ( 
.A(n_6975),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6951),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6979),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_7013),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6977),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6978),
.Y(n_7087)
);

INVx2_ASAP7_75t_L g7088 ( 
.A(n_6904),
.Y(n_7088)
);

NAND3xp33_ASAP7_75t_L g7089 ( 
.A(n_6943),
.B(n_727),
.C(n_728),
.Y(n_7089)
);

OR2x2_ASAP7_75t_L g7090 ( 
.A(n_7014),
.B(n_727),
.Y(n_7090)
);

AND2x4_ASAP7_75t_L g7091 ( 
.A(n_6914),
.B(n_729),
.Y(n_7091)
);

INVx2_ASAP7_75t_L g7092 ( 
.A(n_7004),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6959),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6970),
.Y(n_7094)
);

AND2x2_ASAP7_75t_L g7095 ( 
.A(n_6966),
.B(n_729),
.Y(n_7095)
);

NAND2xp5_ASAP7_75t_L g7096 ( 
.A(n_6990),
.B(n_729),
.Y(n_7096)
);

AND2x2_ASAP7_75t_L g7097 ( 
.A(n_6909),
.B(n_730),
.Y(n_7097)
);

AND2x2_ASAP7_75t_L g7098 ( 
.A(n_6917),
.B(n_730),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6972),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_L g7100 ( 
.A(n_6949),
.B(n_730),
.Y(n_7100)
);

NAND2xp5_ASAP7_75t_L g7101 ( 
.A(n_7005),
.B(n_731),
.Y(n_7101)
);

NAND2xp5_ASAP7_75t_SL g7102 ( 
.A(n_7011),
.B(n_731),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6918),
.Y(n_7103)
);

OAI22xp5_ASAP7_75t_L g7104 ( 
.A1(n_7012),
.A2(n_733),
.B1(n_731),
.B2(n_732),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6955),
.Y(n_7105)
);

OAI22xp33_ASAP7_75t_L g7106 ( 
.A1(n_6915),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.Y(n_7106)
);

AOI32xp33_ASAP7_75t_L g7107 ( 
.A1(n_6995),
.A2(n_735),
.A3(n_733),
.B1(n_734),
.B2(n_736),
.Y(n_7107)
);

AND2x2_ASAP7_75t_L g7108 ( 
.A(n_6944),
.B(n_734),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6960),
.Y(n_7109)
);

OR2x6_ASAP7_75t_L g7110 ( 
.A(n_7003),
.B(n_735),
.Y(n_7110)
);

NAND2xp5_ASAP7_75t_L g7111 ( 
.A(n_6939),
.B(n_735),
.Y(n_7111)
);

INVx1_ASAP7_75t_L g7112 ( 
.A(n_6992),
.Y(n_7112)
);

NOR2xp67_ASAP7_75t_SL g7113 ( 
.A(n_7010),
.B(n_736),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6964),
.Y(n_7114)
);

OR2x2_ASAP7_75t_L g7115 ( 
.A(n_6950),
.B(n_737),
.Y(n_7115)
);

OR2x2_ASAP7_75t_L g7116 ( 
.A(n_6996),
.B(n_6953),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6964),
.Y(n_7117)
);

AND2x2_ASAP7_75t_L g7118 ( 
.A(n_6916),
.B(n_737),
.Y(n_7118)
);

OAI22xp5_ASAP7_75t_L g7119 ( 
.A1(n_6933),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.Y(n_7119)
);

INVx1_ASAP7_75t_L g7120 ( 
.A(n_6969),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_6956),
.Y(n_7121)
);

INVx1_ASAP7_75t_L g7122 ( 
.A(n_6957),
.Y(n_7122)
);

AOI21xp5_ASAP7_75t_L g7123 ( 
.A1(n_6946),
.A2(n_738),
.B(n_739),
.Y(n_7123)
);

AOI32xp33_ASAP7_75t_L g7124 ( 
.A1(n_6967),
.A2(n_741),
.A3(n_739),
.B1(n_740),
.B2(n_743),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6928),
.Y(n_7125)
);

AND2x2_ASAP7_75t_L g7126 ( 
.A(n_6947),
.B(n_740),
.Y(n_7126)
);

INVx3_ASAP7_75t_SL g7127 ( 
.A(n_6936),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_6898),
.Y(n_7128)
);

OAI222xp33_ASAP7_75t_L g7129 ( 
.A1(n_6997),
.A2(n_743),
.B1(n_745),
.B2(n_740),
.C1(n_741),
.C2(n_744),
.Y(n_7129)
);

NAND2xp5_ASAP7_75t_SL g7130 ( 
.A(n_6999),
.B(n_743),
.Y(n_7130)
);

INVx2_ASAP7_75t_SL g7131 ( 
.A(n_6986),
.Y(n_7131)
);

HB1xp67_ASAP7_75t_L g7132 ( 
.A(n_6985),
.Y(n_7132)
);

AND2x2_ASAP7_75t_L g7133 ( 
.A(n_7008),
.B(n_744),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6987),
.Y(n_7134)
);

XNOR2xp5_ASAP7_75t_L g7135 ( 
.A(n_6924),
.B(n_744),
.Y(n_7135)
);

NAND2xp5_ASAP7_75t_L g7136 ( 
.A(n_6901),
.B(n_745),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6901),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_7028),
.Y(n_7138)
);

NOR2xp33_ASAP7_75t_L g7139 ( 
.A(n_7062),
.B(n_746),
.Y(n_7139)
);

INVxp67_ASAP7_75t_L g7140 ( 
.A(n_7018),
.Y(n_7140)
);

OR2x2_ASAP7_75t_L g7141 ( 
.A(n_7038),
.B(n_746),
.Y(n_7141)
);

INVxp67_ASAP7_75t_SL g7142 ( 
.A(n_7049),
.Y(n_7142)
);

BUFx2_ASAP7_75t_L g7143 ( 
.A(n_7067),
.Y(n_7143)
);

INVx1_ASAP7_75t_SL g7144 ( 
.A(n_7070),
.Y(n_7144)
);

INVx1_ASAP7_75t_SL g7145 ( 
.A(n_7029),
.Y(n_7145)
);

AND2x2_ASAP7_75t_L g7146 ( 
.A(n_7095),
.B(n_748),
.Y(n_7146)
);

OR2x2_ASAP7_75t_L g7147 ( 
.A(n_7046),
.B(n_7081),
.Y(n_7147)
);

INVx4_ASAP7_75t_L g7148 ( 
.A(n_7127),
.Y(n_7148)
);

INVx1_ASAP7_75t_L g7149 ( 
.A(n_7042),
.Y(n_7149)
);

INVx1_ASAP7_75t_L g7150 ( 
.A(n_7101),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_7079),
.Y(n_7151)
);

AND2x2_ASAP7_75t_L g7152 ( 
.A(n_7066),
.B(n_749),
.Y(n_7152)
);

NAND2xp33_ASAP7_75t_L g7153 ( 
.A(n_7054),
.B(n_749),
.Y(n_7153)
);

NAND2xp5_ASAP7_75t_L g7154 ( 
.A(n_7061),
.B(n_749),
.Y(n_7154)
);

AND2x2_ASAP7_75t_L g7155 ( 
.A(n_7093),
.B(n_750),
.Y(n_7155)
);

OR2x2_ASAP7_75t_L g7156 ( 
.A(n_7092),
.B(n_750),
.Y(n_7156)
);

OR2x2_ASAP7_75t_L g7157 ( 
.A(n_7076),
.B(n_751),
.Y(n_7157)
);

AND2x2_ASAP7_75t_L g7158 ( 
.A(n_7118),
.B(n_751),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_7113),
.B(n_7072),
.Y(n_7159)
);

OR2x2_ASAP7_75t_L g7160 ( 
.A(n_7019),
.B(n_751),
.Y(n_7160)
);

INVx2_ASAP7_75t_L g7161 ( 
.A(n_7082),
.Y(n_7161)
);

AND2x2_ASAP7_75t_L g7162 ( 
.A(n_7108),
.B(n_752),
.Y(n_7162)
);

OR2x2_ASAP7_75t_L g7163 ( 
.A(n_7020),
.B(n_752),
.Y(n_7163)
);

INVx3_ASAP7_75t_L g7164 ( 
.A(n_7091),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_L g7165 ( 
.A(n_7091),
.B(n_752),
.Y(n_7165)
);

INVx2_ASAP7_75t_L g7166 ( 
.A(n_7088),
.Y(n_7166)
);

HB1xp67_ASAP7_75t_L g7167 ( 
.A(n_7057),
.Y(n_7167)
);

NAND2xp5_ASAP7_75t_L g7168 ( 
.A(n_7097),
.B(n_753),
.Y(n_7168)
);

BUFx2_ASAP7_75t_L g7169 ( 
.A(n_7056),
.Y(n_7169)
);

INVx2_ASAP7_75t_L g7170 ( 
.A(n_7131),
.Y(n_7170)
);

NAND2xp5_ASAP7_75t_L g7171 ( 
.A(n_7098),
.B(n_753),
.Y(n_7171)
);

INVxp67_ASAP7_75t_L g7172 ( 
.A(n_7078),
.Y(n_7172)
);

INVx4_ASAP7_75t_L g7173 ( 
.A(n_7110),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_SL g7174 ( 
.A(n_7106),
.B(n_7060),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_7135),
.Y(n_7175)
);

HB1xp67_ASAP7_75t_L g7176 ( 
.A(n_7094),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_7126),
.Y(n_7177)
);

AND2x4_ASAP7_75t_SL g7178 ( 
.A(n_7031),
.B(n_753),
.Y(n_7178)
);

AOI22xp33_ASAP7_75t_L g7179 ( 
.A1(n_7085),
.A2(n_756),
.B1(n_754),
.B2(n_755),
.Y(n_7179)
);

NAND2xp5_ASAP7_75t_L g7180 ( 
.A(n_7133),
.B(n_754),
.Y(n_7180)
);

NAND2xp5_ASAP7_75t_L g7181 ( 
.A(n_7123),
.B(n_754),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_7069),
.Y(n_7182)
);

OR2x2_ASAP7_75t_L g7183 ( 
.A(n_7068),
.B(n_755),
.Y(n_7183)
);

OAI22xp5_ASAP7_75t_L g7184 ( 
.A1(n_7048),
.A2(n_757),
.B1(n_755),
.B2(n_756),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_7074),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_7114),
.Y(n_7186)
);

INVx2_ASAP7_75t_L g7187 ( 
.A(n_7086),
.Y(n_7187)
);

HB1xp67_ASAP7_75t_L g7188 ( 
.A(n_7017),
.Y(n_7188)
);

INVx1_ASAP7_75t_SL g7189 ( 
.A(n_7087),
.Y(n_7189)
);

AND2x2_ASAP7_75t_L g7190 ( 
.A(n_7033),
.B(n_756),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_7117),
.Y(n_7191)
);

AND2x2_ASAP7_75t_L g7192 ( 
.A(n_7026),
.B(n_758),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_7089),
.Y(n_7193)
);

INVx1_ASAP7_75t_SL g7194 ( 
.A(n_7115),
.Y(n_7194)
);

INVxp67_ASAP7_75t_L g7195 ( 
.A(n_7075),
.Y(n_7195)
);

NAND2xp5_ASAP7_75t_L g7196 ( 
.A(n_7124),
.B(n_758),
.Y(n_7196)
);

BUFx2_ASAP7_75t_L g7197 ( 
.A(n_7110),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_7136),
.Y(n_7198)
);

INVx1_ASAP7_75t_SL g7199 ( 
.A(n_7116),
.Y(n_7199)
);

INVxp67_ASAP7_75t_L g7200 ( 
.A(n_7096),
.Y(n_7200)
);

AO21x2_ASAP7_75t_L g7201 ( 
.A1(n_7037),
.A2(n_7103),
.B(n_7016),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_7071),
.Y(n_7202)
);

INVxp67_ASAP7_75t_L g7203 ( 
.A(n_7111),
.Y(n_7203)
);

AOI22xp33_ASAP7_75t_L g7204 ( 
.A1(n_7104),
.A2(n_761),
.B1(n_759),
.B2(n_760),
.Y(n_7204)
);

OR2x6_ASAP7_75t_L g7205 ( 
.A(n_7121),
.B(n_759),
.Y(n_7205)
);

OR2x2_ASAP7_75t_L g7206 ( 
.A(n_7119),
.B(n_759),
.Y(n_7206)
);

NAND2xp5_ASAP7_75t_L g7207 ( 
.A(n_7107),
.B(n_760),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_7039),
.Y(n_7208)
);

NOR2xp33_ASAP7_75t_L g7209 ( 
.A(n_7148),
.B(n_7058),
.Y(n_7209)
);

AOI22xp5_ASAP7_75t_L g7210 ( 
.A1(n_7145),
.A2(n_7032),
.B1(n_7043),
.B2(n_7034),
.Y(n_7210)
);

INVxp67_ASAP7_75t_L g7211 ( 
.A(n_7167),
.Y(n_7211)
);

OAI22xp5_ASAP7_75t_L g7212 ( 
.A1(n_7140),
.A2(n_7025),
.B1(n_7035),
.B2(n_7063),
.Y(n_7212)
);

NAND2xp5_ASAP7_75t_L g7213 ( 
.A(n_7148),
.B(n_7073),
.Y(n_7213)
);

NAND2xp5_ASAP7_75t_L g7214 ( 
.A(n_7138),
.B(n_7053),
.Y(n_7214)
);

INVxp67_ASAP7_75t_SL g7215 ( 
.A(n_7147),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_7151),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_7142),
.Y(n_7217)
);

AOI22xp33_ASAP7_75t_SL g7218 ( 
.A1(n_7169),
.A2(n_7132),
.B1(n_7125),
.B2(n_7122),
.Y(n_7218)
);

OAI21xp5_ASAP7_75t_L g7219 ( 
.A1(n_7154),
.A2(n_7045),
.B(n_7130),
.Y(n_7219)
);

INVxp67_ASAP7_75t_L g7220 ( 
.A(n_7143),
.Y(n_7220)
);

INVx1_ASAP7_75t_L g7221 ( 
.A(n_7178),
.Y(n_7221)
);

AOI221xp5_ASAP7_75t_L g7222 ( 
.A1(n_7184),
.A2(n_7027),
.B1(n_7129),
.B2(n_7022),
.C(n_7015),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_7165),
.Y(n_7223)
);

INVx3_ASAP7_75t_SL g7224 ( 
.A(n_7144),
.Y(n_7224)
);

NAND2xp5_ASAP7_75t_L g7225 ( 
.A(n_7190),
.B(n_7064),
.Y(n_7225)
);

OAI21xp33_ASAP7_75t_L g7226 ( 
.A1(n_7161),
.A2(n_7041),
.B(n_7084),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_7141),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_7160),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_7163),
.Y(n_7229)
);

OAI21xp5_ASAP7_75t_L g7230 ( 
.A1(n_7139),
.A2(n_7102),
.B(n_7120),
.Y(n_7230)
);

NAND2xp5_ASAP7_75t_L g7231 ( 
.A(n_7192),
.B(n_7047),
.Y(n_7231)
);

OR4x1_ASAP7_75t_L g7232 ( 
.A(n_7149),
.B(n_7099),
.C(n_7052),
.D(n_7040),
.Y(n_7232)
);

NAND3xp33_ASAP7_75t_L g7233 ( 
.A(n_7179),
.B(n_7137),
.C(n_7128),
.Y(n_7233)
);

NOR2xp33_ASAP7_75t_L g7234 ( 
.A(n_7173),
.B(n_7100),
.Y(n_7234)
);

AND2x2_ASAP7_75t_L g7235 ( 
.A(n_7146),
.B(n_7083),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_7166),
.Y(n_7236)
);

INVx1_ASAP7_75t_SL g7237 ( 
.A(n_7199),
.Y(n_7237)
);

NAND2xp5_ASAP7_75t_L g7238 ( 
.A(n_7155),
.B(n_7065),
.Y(n_7238)
);

OR2x2_ASAP7_75t_L g7239 ( 
.A(n_7208),
.B(n_7182),
.Y(n_7239)
);

AND2x2_ASAP7_75t_L g7240 ( 
.A(n_7162),
.B(n_7158),
.Y(n_7240)
);

AND2x2_ASAP7_75t_SL g7241 ( 
.A(n_7153),
.B(n_7173),
.Y(n_7241)
);

INVx2_ASAP7_75t_L g7242 ( 
.A(n_7170),
.Y(n_7242)
);

NOR2xp33_ASAP7_75t_L g7243 ( 
.A(n_7193),
.B(n_7077),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_7188),
.Y(n_7244)
);

INVx1_ASAP7_75t_SL g7245 ( 
.A(n_7189),
.Y(n_7245)
);

AOI211xp5_ASAP7_75t_SL g7246 ( 
.A1(n_7172),
.A2(n_7134),
.B(n_7023),
.C(n_7030),
.Y(n_7246)
);

OAI22xp5_ASAP7_75t_L g7247 ( 
.A1(n_7196),
.A2(n_7090),
.B1(n_7021),
.B2(n_7036),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_7157),
.Y(n_7248)
);

OAI22xp5_ASAP7_75t_L g7249 ( 
.A1(n_7159),
.A2(n_7050),
.B1(n_7044),
.B2(n_7055),
.Y(n_7249)
);

OAI221xp5_ASAP7_75t_L g7250 ( 
.A1(n_7204),
.A2(n_7059),
.B1(n_7051),
.B2(n_7024),
.C(n_7105),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_7176),
.Y(n_7251)
);

AND2x2_ASAP7_75t_L g7252 ( 
.A(n_7152),
.B(n_7164),
.Y(n_7252)
);

INVxp67_ASAP7_75t_SL g7253 ( 
.A(n_7156),
.Y(n_7253)
);

NOR3xp33_ASAP7_75t_L g7254 ( 
.A(n_7187),
.B(n_7080),
.C(n_7109),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_7205),
.Y(n_7255)
);

INVx1_ASAP7_75t_L g7256 ( 
.A(n_7205),
.Y(n_7256)
);

INVx1_ASAP7_75t_SL g7257 ( 
.A(n_7194),
.Y(n_7257)
);

NOR2xp33_ASAP7_75t_L g7258 ( 
.A(n_7168),
.B(n_7112),
.Y(n_7258)
);

NOR3xp33_ASAP7_75t_L g7259 ( 
.A(n_7181),
.B(n_761),
.C(n_762),
.Y(n_7259)
);

OAI22xp5_ASAP7_75t_L g7260 ( 
.A1(n_7207),
.A2(n_763),
.B1(n_761),
.B2(n_762),
.Y(n_7260)
);

OAI22xp33_ASAP7_75t_L g7261 ( 
.A1(n_7171),
.A2(n_765),
.B1(n_763),
.B2(n_764),
.Y(n_7261)
);

AOI22xp5_ASAP7_75t_L g7262 ( 
.A1(n_7202),
.A2(n_7175),
.B1(n_7174),
.B2(n_7180),
.Y(n_7262)
);

INVx3_ASAP7_75t_SL g7263 ( 
.A(n_7183),
.Y(n_7263)
);

O2A1O1Ixp5_ASAP7_75t_L g7264 ( 
.A1(n_7177),
.A2(n_765),
.B(n_763),
.C(n_764),
.Y(n_7264)
);

INVx2_ASAP7_75t_L g7265 ( 
.A(n_7186),
.Y(n_7265)
);

AOI21xp33_ASAP7_75t_L g7266 ( 
.A1(n_7206),
.A2(n_7201),
.B(n_7150),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_7197),
.Y(n_7267)
);

OAI21xp33_ASAP7_75t_L g7268 ( 
.A1(n_7185),
.A2(n_765),
.B(n_766),
.Y(n_7268)
);

AOI221xp5_ASAP7_75t_L g7269 ( 
.A1(n_7195),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.C(n_769),
.Y(n_7269)
);

AOI22xp33_ASAP7_75t_L g7270 ( 
.A1(n_7198),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.Y(n_7270)
);

NAND2xp5_ASAP7_75t_SL g7271 ( 
.A(n_7191),
.B(n_767),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_7203),
.Y(n_7272)
);

OR2x2_ASAP7_75t_L g7273 ( 
.A(n_7200),
.B(n_768),
.Y(n_7273)
);

AND2x2_ASAP7_75t_L g7274 ( 
.A(n_7148),
.B(n_769),
.Y(n_7274)
);

INVx1_ASAP7_75t_L g7275 ( 
.A(n_7147),
.Y(n_7275)
);

INVx2_ASAP7_75t_L g7276 ( 
.A(n_7148),
.Y(n_7276)
);

AOI22xp5_ASAP7_75t_L g7277 ( 
.A1(n_7145),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_7277)
);

OAI211xp5_ASAP7_75t_SL g7278 ( 
.A1(n_7140),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_7278)
);

OR2x2_ASAP7_75t_L g7279 ( 
.A(n_7148),
.B(n_770),
.Y(n_7279)
);

INVx2_ASAP7_75t_L g7280 ( 
.A(n_7148),
.Y(n_7280)
);

NAND2xp5_ASAP7_75t_L g7281 ( 
.A(n_7148),
.B(n_771),
.Y(n_7281)
);

AOI322xp5_ASAP7_75t_L g7282 ( 
.A1(n_7145),
.A2(n_772),
.A3(n_773),
.B1(n_774),
.B2(n_775),
.C1(n_776),
.C2(n_777),
.Y(n_7282)
);

AND2x2_ASAP7_75t_L g7283 ( 
.A(n_7148),
.B(n_773),
.Y(n_7283)
);

INVx1_ASAP7_75t_SL g7284 ( 
.A(n_7147),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_7147),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_7147),
.Y(n_7286)
);

OAI21xp5_ASAP7_75t_L g7287 ( 
.A1(n_7140),
.A2(n_773),
.B(n_774),
.Y(n_7287)
);

INVx2_ASAP7_75t_L g7288 ( 
.A(n_7148),
.Y(n_7288)
);

OAI22xp33_ASAP7_75t_L g7289 ( 
.A1(n_7145),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_7289)
);

OAI21xp33_ASAP7_75t_L g7290 ( 
.A1(n_7144),
.A2(n_776),
.B(n_777),
.Y(n_7290)
);

OAI22xp5_ASAP7_75t_L g7291 ( 
.A1(n_7140),
.A2(n_779),
.B1(n_777),
.B2(n_778),
.Y(n_7291)
);

INVx1_ASAP7_75t_SL g7292 ( 
.A(n_7147),
.Y(n_7292)
);

AND2x2_ASAP7_75t_L g7293 ( 
.A(n_7148),
.B(n_778),
.Y(n_7293)
);

INVxp67_ASAP7_75t_L g7294 ( 
.A(n_7215),
.Y(n_7294)
);

AND2x2_ASAP7_75t_L g7295 ( 
.A(n_7284),
.B(n_7292),
.Y(n_7295)
);

NAND2xp5_ASAP7_75t_L g7296 ( 
.A(n_7224),
.B(n_778),
.Y(n_7296)
);

OAI21xp33_ASAP7_75t_SL g7297 ( 
.A1(n_7209),
.A2(n_779),
.B(n_780),
.Y(n_7297)
);

OAI22xp5_ASAP7_75t_L g7298 ( 
.A1(n_7239),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_7214),
.Y(n_7299)
);

AND2x2_ASAP7_75t_L g7300 ( 
.A(n_7276),
.B(n_7280),
.Y(n_7300)
);

OA21x2_ASAP7_75t_L g7301 ( 
.A1(n_7281),
.A2(n_780),
.B(n_781),
.Y(n_7301)
);

NAND3xp33_ASAP7_75t_L g7302 ( 
.A(n_7282),
.B(n_781),
.C(n_782),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_7275),
.Y(n_7303)
);

AOI22xp5_ASAP7_75t_L g7304 ( 
.A1(n_7285),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_7286),
.Y(n_7305)
);

AND2x4_ASAP7_75t_L g7306 ( 
.A(n_7288),
.B(n_783),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7274),
.Y(n_7307)
);

OR2x2_ASAP7_75t_L g7308 ( 
.A(n_7237),
.B(n_784),
.Y(n_7308)
);

AOI222xp33_ASAP7_75t_L g7309 ( 
.A1(n_7236),
.A2(n_786),
.B1(n_788),
.B2(n_784),
.C1(n_785),
.C2(n_787),
.Y(n_7309)
);

AND2x2_ASAP7_75t_L g7310 ( 
.A(n_7242),
.B(n_785),
.Y(n_7310)
);

OR2x2_ASAP7_75t_L g7311 ( 
.A(n_7216),
.B(n_786),
.Y(n_7311)
);

AND2x2_ASAP7_75t_L g7312 ( 
.A(n_7252),
.B(n_787),
.Y(n_7312)
);

NAND2xp5_ASAP7_75t_L g7313 ( 
.A(n_7283),
.B(n_7293),
.Y(n_7313)
);

OAI221xp5_ASAP7_75t_L g7314 ( 
.A1(n_7218),
.A2(n_7290),
.B1(n_7270),
.B2(n_7210),
.C(n_7269),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_7279),
.Y(n_7315)
);

INVx2_ASAP7_75t_SL g7316 ( 
.A(n_7221),
.Y(n_7316)
);

O2A1O1Ixp33_ASAP7_75t_L g7317 ( 
.A1(n_7291),
.A2(n_790),
.B(n_788),
.C(n_789),
.Y(n_7317)
);

INVx1_ASAP7_75t_SL g7318 ( 
.A(n_7245),
.Y(n_7318)
);

A2O1A1Ixp33_ASAP7_75t_L g7319 ( 
.A1(n_7264),
.A2(n_7268),
.B(n_7226),
.C(n_7220),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_7277),
.Y(n_7320)
);

NOR3xp33_ASAP7_75t_L g7321 ( 
.A(n_7213),
.B(n_788),
.C(n_789),
.Y(n_7321)
);

NAND2xp5_ASAP7_75t_L g7322 ( 
.A(n_7277),
.B(n_790),
.Y(n_7322)
);

INVx2_ASAP7_75t_L g7323 ( 
.A(n_7217),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_7273),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_7244),
.Y(n_7325)
);

INVx1_ASAP7_75t_L g7326 ( 
.A(n_7251),
.Y(n_7326)
);

AOI221xp5_ASAP7_75t_L g7327 ( 
.A1(n_7289),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.C(n_794),
.Y(n_7327)
);

OAI21xp33_ASAP7_75t_L g7328 ( 
.A1(n_7262),
.A2(n_7257),
.B(n_7243),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_7253),
.Y(n_7329)
);

OR2x2_ASAP7_75t_L g7330 ( 
.A(n_7211),
.B(n_791),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_7235),
.Y(n_7331)
);

INVx1_ASAP7_75t_L g7332 ( 
.A(n_7231),
.Y(n_7332)
);

AND2x2_ASAP7_75t_L g7333 ( 
.A(n_7240),
.B(n_792),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_7225),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_7238),
.Y(n_7335)
);

CKINVDCx14_ASAP7_75t_R g7336 ( 
.A(n_7234),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_7241),
.Y(n_7337)
);

NOR2x1_ASAP7_75t_L g7338 ( 
.A(n_7302),
.B(n_7233),
.Y(n_7338)
);

AND2x2_ASAP7_75t_L g7339 ( 
.A(n_7295),
.B(n_7267),
.Y(n_7339)
);

NAND2xp5_ASAP7_75t_L g7340 ( 
.A(n_7300),
.B(n_7222),
.Y(n_7340)
);

NAND2xp5_ASAP7_75t_L g7341 ( 
.A(n_7294),
.B(n_7261),
.Y(n_7341)
);

INVx3_ASAP7_75t_SL g7342 ( 
.A(n_7316),
.Y(n_7342)
);

AND2x2_ASAP7_75t_L g7343 ( 
.A(n_7312),
.B(n_7263),
.Y(n_7343)
);

AND2x2_ASAP7_75t_L g7344 ( 
.A(n_7318),
.B(n_7227),
.Y(n_7344)
);

NOR2xp33_ASAP7_75t_L g7345 ( 
.A(n_7299),
.B(n_7265),
.Y(n_7345)
);

NOR2xp33_ASAP7_75t_L g7346 ( 
.A(n_7328),
.B(n_7260),
.Y(n_7346)
);

NOR2xp33_ASAP7_75t_L g7347 ( 
.A(n_7303),
.B(n_7250),
.Y(n_7347)
);

INVx1_ASAP7_75t_SL g7348 ( 
.A(n_7306),
.Y(n_7348)
);

AND2x2_ASAP7_75t_L g7349 ( 
.A(n_7333),
.B(n_7228),
.Y(n_7349)
);

OR2x2_ASAP7_75t_L g7350 ( 
.A(n_7331),
.B(n_7229),
.Y(n_7350)
);

NAND2x1_ASAP7_75t_L g7351 ( 
.A(n_7323),
.B(n_7255),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_7310),
.Y(n_7352)
);

NAND2xp5_ASAP7_75t_L g7353 ( 
.A(n_7309),
.B(n_7254),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_7296),
.Y(n_7354)
);

CKINVDCx5p33_ASAP7_75t_R g7355 ( 
.A(n_7336),
.Y(n_7355)
);

NAND2x1_ASAP7_75t_L g7356 ( 
.A(n_7305),
.B(n_7256),
.Y(n_7356)
);

HB1xp67_ASAP7_75t_L g7357 ( 
.A(n_7329),
.Y(n_7357)
);

INVx2_ASAP7_75t_L g7358 ( 
.A(n_7325),
.Y(n_7358)
);

NAND2xp5_ASAP7_75t_L g7359 ( 
.A(n_7304),
.B(n_7259),
.Y(n_7359)
);

INVx2_ASAP7_75t_SL g7360 ( 
.A(n_7337),
.Y(n_7360)
);

NAND2xp5_ASAP7_75t_L g7361 ( 
.A(n_7332),
.B(n_7246),
.Y(n_7361)
);

NAND2xp5_ASAP7_75t_L g7362 ( 
.A(n_7334),
.B(n_7248),
.Y(n_7362)
);

INVx2_ASAP7_75t_SL g7363 ( 
.A(n_7311),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_7330),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_7322),
.Y(n_7365)
);

OR2x2_ASAP7_75t_L g7366 ( 
.A(n_7313),
.B(n_7249),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_L g7367 ( 
.A(n_7321),
.B(n_7258),
.Y(n_7367)
);

NAND2xp5_ASAP7_75t_L g7368 ( 
.A(n_7301),
.B(n_7287),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_7308),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_7301),
.Y(n_7370)
);

INVxp67_ASAP7_75t_L g7371 ( 
.A(n_7326),
.Y(n_7371)
);

NAND2xp5_ASAP7_75t_SL g7372 ( 
.A(n_7297),
.B(n_7320),
.Y(n_7372)
);

AND2x2_ASAP7_75t_L g7373 ( 
.A(n_7335),
.B(n_7219),
.Y(n_7373)
);

NOR2xp33_ASAP7_75t_L g7374 ( 
.A(n_7314),
.B(n_7271),
.Y(n_7374)
);

AND2x4_ASAP7_75t_L g7375 ( 
.A(n_7315),
.B(n_7272),
.Y(n_7375)
);

NAND2xp5_ASAP7_75t_L g7376 ( 
.A(n_7327),
.B(n_7212),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_7298),
.Y(n_7377)
);

INVx1_ASAP7_75t_SL g7378 ( 
.A(n_7324),
.Y(n_7378)
);

INVxp67_ASAP7_75t_L g7379 ( 
.A(n_7307),
.Y(n_7379)
);

NOR2xp33_ASAP7_75t_L g7380 ( 
.A(n_7319),
.B(n_7266),
.Y(n_7380)
);

OR2x2_ASAP7_75t_L g7381 ( 
.A(n_7317),
.B(n_7247),
.Y(n_7381)
);

NAND2xp5_ASAP7_75t_L g7382 ( 
.A(n_7295),
.B(n_7223),
.Y(n_7382)
);

NOR2xp33_ASAP7_75t_L g7383 ( 
.A(n_7294),
.B(n_7278),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_7300),
.Y(n_7384)
);

AOI211xp5_ASAP7_75t_L g7385 ( 
.A1(n_7342),
.A2(n_7230),
.B(n_7232),
.C(n_794),
.Y(n_7385)
);

NOR4xp25_ASAP7_75t_L g7386 ( 
.A(n_7340),
.B(n_795),
.C(n_792),
.D(n_793),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_7384),
.Y(n_7387)
);

NOR3x1_ASAP7_75t_L g7388 ( 
.A(n_7361),
.B(n_793),
.C(n_795),
.Y(n_7388)
);

NOR3xp33_ASAP7_75t_L g7389 ( 
.A(n_7372),
.B(n_796),
.C(n_797),
.Y(n_7389)
);

NAND3xp33_ASAP7_75t_L g7390 ( 
.A(n_7380),
.B(n_796),
.C(n_797),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_7339),
.Y(n_7391)
);

AOI221xp5_ASAP7_75t_L g7392 ( 
.A1(n_7347),
.A2(n_7345),
.B1(n_7371),
.B2(n_7374),
.C(n_7346),
.Y(n_7392)
);

NOR2x1_ASAP7_75t_L g7393 ( 
.A(n_7370),
.B(n_796),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7357),
.Y(n_7394)
);

AOI221xp5_ASAP7_75t_L g7395 ( 
.A1(n_7379),
.A2(n_7383),
.B1(n_7355),
.B2(n_7378),
.C(n_7353),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_7366),
.Y(n_7396)
);

AOI211xp5_ASAP7_75t_L g7397 ( 
.A1(n_7344),
.A2(n_799),
.B(n_797),
.C(n_798),
.Y(n_7397)
);

NAND2x1_ASAP7_75t_L g7398 ( 
.A(n_7375),
.B(n_798),
.Y(n_7398)
);

NAND3xp33_ASAP7_75t_L g7399 ( 
.A(n_7338),
.B(n_798),
.C(n_799),
.Y(n_7399)
);

INVxp67_ASAP7_75t_SL g7400 ( 
.A(n_7382),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_L g7401 ( 
.A(n_7343),
.B(n_799),
.Y(n_7401)
);

NAND2xp5_ASAP7_75t_L g7402 ( 
.A(n_7375),
.B(n_800),
.Y(n_7402)
);

NOR3xp33_ASAP7_75t_L g7403 ( 
.A(n_7362),
.B(n_800),
.C(n_801),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_7349),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_7350),
.Y(n_7405)
);

NOR2xp33_ASAP7_75t_SL g7406 ( 
.A(n_7348),
.B(n_800),
.Y(n_7406)
);

NAND3xp33_ASAP7_75t_SL g7407 ( 
.A(n_7351),
.B(n_801),
.C(n_802),
.Y(n_7407)
);

NAND2xp5_ASAP7_75t_L g7408 ( 
.A(n_7358),
.B(n_802),
.Y(n_7408)
);

NAND3xp33_ASAP7_75t_SL g7409 ( 
.A(n_7356),
.B(n_803),
.C(n_804),
.Y(n_7409)
);

OAI21xp33_ASAP7_75t_SL g7410 ( 
.A1(n_7376),
.A2(n_7341),
.B(n_7360),
.Y(n_7410)
);

INVx1_ASAP7_75t_SL g7411 ( 
.A(n_7373),
.Y(n_7411)
);

NAND3xp33_ASAP7_75t_L g7412 ( 
.A(n_7377),
.B(n_803),
.C(n_804),
.Y(n_7412)
);

AOI21xp5_ASAP7_75t_L g7413 ( 
.A1(n_7368),
.A2(n_803),
.B(n_806),
.Y(n_7413)
);

AOI221x1_ASAP7_75t_L g7414 ( 
.A1(n_7364),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.C(n_809),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_7381),
.Y(n_7415)
);

NOR2xp33_ASAP7_75t_L g7416 ( 
.A(n_7352),
.B(n_807),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7396),
.Y(n_7417)
);

AND4x1_ASAP7_75t_L g7418 ( 
.A(n_7395),
.B(n_7392),
.C(n_7385),
.D(n_7406),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_7400),
.Y(n_7419)
);

OR2x2_ASAP7_75t_L g7420 ( 
.A(n_7411),
.B(n_7363),
.Y(n_7420)
);

NAND3xp33_ASAP7_75t_L g7421 ( 
.A(n_7397),
.B(n_7369),
.C(n_7367),
.Y(n_7421)
);

NAND3xp33_ASAP7_75t_SL g7422 ( 
.A(n_7389),
.B(n_7359),
.C(n_7365),
.Y(n_7422)
);

NOR4xp25_ASAP7_75t_L g7423 ( 
.A(n_7410),
.B(n_7354),
.C(n_810),
.D(n_808),
.Y(n_7423)
);

INVx1_ASAP7_75t_L g7424 ( 
.A(n_7393),
.Y(n_7424)
);

NOR2x1_ASAP7_75t_L g7425 ( 
.A(n_7415),
.B(n_808),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_7402),
.Y(n_7426)
);

NAND2xp5_ASAP7_75t_SL g7427 ( 
.A(n_7391),
.B(n_809),
.Y(n_7427)
);

AO221x1_ASAP7_75t_L g7428 ( 
.A1(n_7405),
.A2(n_7387),
.B1(n_7404),
.B2(n_7394),
.C(n_7388),
.Y(n_7428)
);

AND2x2_ASAP7_75t_L g7429 ( 
.A(n_7416),
.B(n_809),
.Y(n_7429)
);

AOI21xp5_ASAP7_75t_L g7430 ( 
.A1(n_7413),
.A2(n_810),
.B(n_811),
.Y(n_7430)
);

NOR3xp33_ASAP7_75t_L g7431 ( 
.A(n_7412),
.B(n_810),
.C(n_811),
.Y(n_7431)
);

NAND2x1_ASAP7_75t_SL g7432 ( 
.A(n_7386),
.B(n_812),
.Y(n_7432)
);

NOR3x1_ASAP7_75t_L g7433 ( 
.A(n_7401),
.B(n_7390),
.C(n_7399),
.Y(n_7433)
);

NOR2xp33_ASAP7_75t_L g7434 ( 
.A(n_7408),
.B(n_812),
.Y(n_7434)
);

NOR3xp33_ASAP7_75t_L g7435 ( 
.A(n_7409),
.B(n_812),
.C(n_813),
.Y(n_7435)
);

INVx1_ASAP7_75t_SL g7436 ( 
.A(n_7398),
.Y(n_7436)
);

NAND2xp5_ASAP7_75t_L g7437 ( 
.A(n_7403),
.B(n_813),
.Y(n_7437)
);

NAND4xp25_ASAP7_75t_L g7438 ( 
.A(n_7414),
.B(n_815),
.C(n_813),
.D(n_814),
.Y(n_7438)
);

NAND2xp5_ASAP7_75t_L g7439 ( 
.A(n_7407),
.B(n_814),
.Y(n_7439)
);

CKINVDCx5p33_ASAP7_75t_R g7440 ( 
.A(n_7411),
.Y(n_7440)
);

HB1xp67_ASAP7_75t_L g7441 ( 
.A(n_7396),
.Y(n_7441)
);

AND2x2_ASAP7_75t_L g7442 ( 
.A(n_7400),
.B(n_814),
.Y(n_7442)
);

INVx2_ASAP7_75t_L g7443 ( 
.A(n_7396),
.Y(n_7443)
);

NOR4xp25_ASAP7_75t_L g7444 ( 
.A(n_7410),
.B(n_817),
.C(n_815),
.D(n_816),
.Y(n_7444)
);

NAND2xp5_ASAP7_75t_L g7445 ( 
.A(n_7396),
.B(n_816),
.Y(n_7445)
);

INVx2_ASAP7_75t_L g7446 ( 
.A(n_7396),
.Y(n_7446)
);

NOR3xp33_ASAP7_75t_L g7447 ( 
.A(n_7410),
.B(n_817),
.C(n_819),
.Y(n_7447)
);

INVxp67_ASAP7_75t_L g7448 ( 
.A(n_7406),
.Y(n_7448)
);

NOR3xp33_ASAP7_75t_L g7449 ( 
.A(n_7410),
.B(n_819),
.C(n_820),
.Y(n_7449)
);

NAND2xp5_ASAP7_75t_L g7450 ( 
.A(n_7396),
.B(n_819),
.Y(n_7450)
);

AOI211xp5_ASAP7_75t_L g7451 ( 
.A1(n_7410),
.A2(n_822),
.B(n_820),
.C(n_821),
.Y(n_7451)
);

AND2x2_ASAP7_75t_L g7452 ( 
.A(n_7400),
.B(n_821),
.Y(n_7452)
);

NAND3xp33_ASAP7_75t_SL g7453 ( 
.A(n_7385),
.B(n_822),
.C(n_823),
.Y(n_7453)
);

OAI211xp5_ASAP7_75t_SL g7454 ( 
.A1(n_7395),
.A2(n_824),
.B(n_822),
.C(n_823),
.Y(n_7454)
);

NAND4xp25_ASAP7_75t_L g7455 ( 
.A(n_7395),
.B(n_826),
.C(n_824),
.D(n_825),
.Y(n_7455)
);

OR2x6_ASAP7_75t_L g7456 ( 
.A(n_7396),
.B(n_825),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7442),
.Y(n_7457)
);

NOR2xp33_ASAP7_75t_L g7458 ( 
.A(n_7419),
.B(n_825),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_7452),
.Y(n_7459)
);

OA22x2_ASAP7_75t_L g7460 ( 
.A1(n_7428),
.A2(n_828),
.B1(n_826),
.B2(n_827),
.Y(n_7460)
);

NAND2xp33_ASAP7_75t_L g7461 ( 
.A(n_7440),
.B(n_826),
.Y(n_7461)
);

AOI32xp33_ASAP7_75t_L g7462 ( 
.A1(n_7417),
.A2(n_829),
.A3(n_827),
.B1(n_828),
.B2(n_830),
.Y(n_7462)
);

INVxp67_ASAP7_75t_L g7463 ( 
.A(n_7441),
.Y(n_7463)
);

NOR3xp33_ASAP7_75t_L g7464 ( 
.A(n_7453),
.B(n_827),
.C(n_828),
.Y(n_7464)
);

AOI211xp5_ASAP7_75t_SL g7465 ( 
.A1(n_7434),
.A2(n_832),
.B(n_829),
.C(n_831),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_7445),
.Y(n_7466)
);

AOI221xp5_ASAP7_75t_L g7467 ( 
.A1(n_7444),
.A2(n_832),
.B1(n_829),
.B2(n_831),
.C(n_833),
.Y(n_7467)
);

O2A1O1Ixp33_ASAP7_75t_L g7468 ( 
.A1(n_7427),
.A2(n_833),
.B(n_831),
.C(n_832),
.Y(n_7468)
);

NOR2xp33_ASAP7_75t_L g7469 ( 
.A(n_7443),
.B(n_834),
.Y(n_7469)
);

AOI222xp33_ASAP7_75t_L g7470 ( 
.A1(n_7446),
.A2(n_834),
.B1(n_835),
.B2(n_836),
.C1(n_837),
.C2(n_838),
.Y(n_7470)
);

NAND2xp33_ASAP7_75t_SL g7471 ( 
.A(n_7420),
.B(n_835),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_7450),
.Y(n_7472)
);

NOR2x1_ASAP7_75t_L g7473 ( 
.A(n_7421),
.B(n_835),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_7451),
.B(n_836),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7456),
.Y(n_7475)
);

NAND4xp25_ASAP7_75t_L g7476 ( 
.A(n_7433),
.B(n_839),
.C(n_836),
.D(n_837),
.Y(n_7476)
);

NAND2xp5_ASAP7_75t_L g7477 ( 
.A(n_7447),
.B(n_837),
.Y(n_7477)
);

OAI22xp33_ASAP7_75t_L g7478 ( 
.A1(n_7439),
.A2(n_841),
.B1(n_839),
.B2(n_840),
.Y(n_7478)
);

BUFx2_ASAP7_75t_L g7479 ( 
.A(n_7456),
.Y(n_7479)
);

OAI21xp5_ASAP7_75t_L g7480 ( 
.A1(n_7430),
.A2(n_839),
.B(n_840),
.Y(n_7480)
);

OA22x2_ASAP7_75t_L g7481 ( 
.A1(n_7437),
.A2(n_842),
.B1(n_840),
.B2(n_841),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_7425),
.Y(n_7482)
);

NAND2xp5_ASAP7_75t_L g7483 ( 
.A(n_7449),
.B(n_842),
.Y(n_7483)
);

INVx2_ASAP7_75t_L g7484 ( 
.A(n_7426),
.Y(n_7484)
);

NAND2xp5_ASAP7_75t_L g7485 ( 
.A(n_7423),
.B(n_843),
.Y(n_7485)
);

OR2x2_ASAP7_75t_L g7486 ( 
.A(n_7455),
.B(n_843),
.Y(n_7486)
);

OAI21xp5_ASAP7_75t_L g7487 ( 
.A1(n_7431),
.A2(n_844),
.B(n_845),
.Y(n_7487)
);

HB1xp67_ASAP7_75t_L g7488 ( 
.A(n_7418),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_7429),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_7432),
.Y(n_7490)
);

OAI211xp5_ASAP7_75t_L g7491 ( 
.A1(n_7454),
.A2(n_846),
.B(n_844),
.C(n_845),
.Y(n_7491)
);

INVx1_ASAP7_75t_SL g7492 ( 
.A(n_7436),
.Y(n_7492)
);

INVxp67_ASAP7_75t_SL g7493 ( 
.A(n_7463),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_7460),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7485),
.Y(n_7495)
);

INVxp67_ASAP7_75t_SL g7496 ( 
.A(n_7468),
.Y(n_7496)
);

AOI221xp5_ASAP7_75t_L g7497 ( 
.A1(n_7478),
.A2(n_7435),
.B1(n_7438),
.B2(n_7422),
.C(n_7448),
.Y(n_7497)
);

INVx2_ASAP7_75t_L g7498 ( 
.A(n_7492),
.Y(n_7498)
);

AOI221xp5_ASAP7_75t_L g7499 ( 
.A1(n_7476),
.A2(n_7424),
.B1(n_846),
.B2(n_844),
.C(n_845),
.Y(n_7499)
);

AO22x2_ASAP7_75t_L g7500 ( 
.A1(n_7457),
.A2(n_848),
.B1(n_846),
.B2(n_847),
.Y(n_7500)
);

NOR2xp67_ASAP7_75t_L g7501 ( 
.A(n_7488),
.B(n_847),
.Y(n_7501)
);

NOR2x1_ASAP7_75t_L g7502 ( 
.A(n_7473),
.B(n_847),
.Y(n_7502)
);

AOI22xp5_ASAP7_75t_L g7503 ( 
.A1(n_7458),
.A2(n_850),
.B1(n_848),
.B2(n_849),
.Y(n_7503)
);

AO22x2_ASAP7_75t_L g7504 ( 
.A1(n_7459),
.A2(n_850),
.B1(n_848),
.B2(n_849),
.Y(n_7504)
);

NOR4xp25_ASAP7_75t_L g7505 ( 
.A(n_7491),
.B(n_852),
.C(n_850),
.D(n_851),
.Y(n_7505)
);

NAND2xp5_ASAP7_75t_L g7506 ( 
.A(n_7470),
.B(n_851),
.Y(n_7506)
);

AOI22xp5_ASAP7_75t_L g7507 ( 
.A1(n_7469),
.A2(n_853),
.B1(n_851),
.B2(n_852),
.Y(n_7507)
);

INVx1_ASAP7_75t_L g7508 ( 
.A(n_7481),
.Y(n_7508)
);

OAI22xp5_ASAP7_75t_SL g7509 ( 
.A1(n_7477),
.A2(n_855),
.B1(n_853),
.B2(n_854),
.Y(n_7509)
);

AOI22xp5_ASAP7_75t_L g7510 ( 
.A1(n_7484),
.A2(n_856),
.B1(n_854),
.B2(n_855),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_7483),
.Y(n_7511)
);

AOI22xp5_ASAP7_75t_L g7512 ( 
.A1(n_7464),
.A2(n_858),
.B1(n_856),
.B2(n_857),
.Y(n_7512)
);

NAND2xp5_ASAP7_75t_L g7513 ( 
.A(n_7462),
.B(n_857),
.Y(n_7513)
);

AOI22xp5_ASAP7_75t_L g7514 ( 
.A1(n_7489),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_7514)
);

AO22x1_ASAP7_75t_L g7515 ( 
.A1(n_7487),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_7515)
);

INVxp67_ASAP7_75t_SL g7516 ( 
.A(n_7474),
.Y(n_7516)
);

NOR2x1_ASAP7_75t_L g7517 ( 
.A(n_7486),
.B(n_859),
.Y(n_7517)
);

NAND2xp5_ASAP7_75t_SL g7518 ( 
.A(n_7498),
.B(n_7475),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_7504),
.Y(n_7519)
);

NAND2xp5_ASAP7_75t_L g7520 ( 
.A(n_7493),
.B(n_7467),
.Y(n_7520)
);

NOR3xp33_ASAP7_75t_L g7521 ( 
.A(n_7497),
.B(n_7472),
.C(n_7466),
.Y(n_7521)
);

AOI221xp5_ASAP7_75t_L g7522 ( 
.A1(n_7499),
.A2(n_7471),
.B1(n_7480),
.B2(n_7461),
.C(n_7490),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7504),
.Y(n_7523)
);

INVx1_ASAP7_75t_SL g7524 ( 
.A(n_7506),
.Y(n_7524)
);

NAND2xp5_ASAP7_75t_L g7525 ( 
.A(n_7501),
.B(n_7465),
.Y(n_7525)
);

INVxp33_ASAP7_75t_L g7526 ( 
.A(n_7517),
.Y(n_7526)
);

OR2x2_ASAP7_75t_L g7527 ( 
.A(n_7513),
.B(n_7479),
.Y(n_7527)
);

AND2x4_ASAP7_75t_L g7528 ( 
.A(n_7496),
.B(n_7482),
.Y(n_7528)
);

NOR2x1_ASAP7_75t_L g7529 ( 
.A(n_7494),
.B(n_860),
.Y(n_7529)
);

INVx1_ASAP7_75t_L g7530 ( 
.A(n_7500),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7514),
.Y(n_7531)
);

INVx3_ASAP7_75t_L g7532 ( 
.A(n_7508),
.Y(n_7532)
);

NAND2xp5_ASAP7_75t_L g7533 ( 
.A(n_7510),
.B(n_860),
.Y(n_7533)
);

OAI22xp5_ASAP7_75t_L g7534 ( 
.A1(n_7495),
.A2(n_863),
.B1(n_861),
.B2(n_862),
.Y(n_7534)
);

INVx1_ASAP7_75t_L g7535 ( 
.A(n_7509),
.Y(n_7535)
);

NOR2x1_ASAP7_75t_L g7536 ( 
.A(n_7502),
.B(n_861),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7529),
.Y(n_7537)
);

NOR3xp33_ASAP7_75t_L g7538 ( 
.A(n_7521),
.B(n_7516),
.C(n_7511),
.Y(n_7538)
);

NAND2x1p5_ASAP7_75t_L g7539 ( 
.A(n_7532),
.B(n_7512),
.Y(n_7539)
);

AND2x2_ASAP7_75t_L g7540 ( 
.A(n_7528),
.B(n_7505),
.Y(n_7540)
);

AND2x2_ASAP7_75t_L g7541 ( 
.A(n_7518),
.B(n_7526),
.Y(n_7541)
);

INVx2_ASAP7_75t_L g7542 ( 
.A(n_7530),
.Y(n_7542)
);

NOR2x1_ASAP7_75t_L g7543 ( 
.A(n_7520),
.B(n_7515),
.Y(n_7543)
);

NOR4xp25_ASAP7_75t_L g7544 ( 
.A(n_7524),
.B(n_7507),
.C(n_7503),
.D(n_863),
.Y(n_7544)
);

NAND4xp25_ASAP7_75t_L g7545 ( 
.A(n_7527),
.B(n_863),
.C(n_861),
.D(n_862),
.Y(n_7545)
);

BUFx2_ASAP7_75t_L g7546 ( 
.A(n_7519),
.Y(n_7546)
);

NOR2x1_ASAP7_75t_L g7547 ( 
.A(n_7523),
.B(n_1008),
.Y(n_7547)
);

AND2x2_ASAP7_75t_L g7548 ( 
.A(n_7538),
.B(n_7535),
.Y(n_7548)
);

NAND3x1_ASAP7_75t_L g7549 ( 
.A(n_7543),
.B(n_7536),
.C(n_7525),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7542),
.Y(n_7550)
);

INVx2_ASAP7_75t_L g7551 ( 
.A(n_7541),
.Y(n_7551)
);

NAND3x1_ASAP7_75t_L g7552 ( 
.A(n_7548),
.B(n_7540),
.C(n_7522),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_7551),
.Y(n_7553)
);

OAI22xp5_ASAP7_75t_L g7554 ( 
.A1(n_7552),
.A2(n_7539),
.B1(n_7549),
.B2(n_7531),
.Y(n_7554)
);

INVx2_ASAP7_75t_L g7555 ( 
.A(n_7553),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7554),
.Y(n_7556)
);

NAND2xp33_ASAP7_75t_R g7557 ( 
.A(n_7555),
.B(n_7546),
.Y(n_7557)
);

NAND2xp5_ASAP7_75t_SL g7558 ( 
.A(n_7557),
.B(n_7550),
.Y(n_7558)
);

OR2x2_ASAP7_75t_L g7559 ( 
.A(n_7556),
.B(n_7537),
.Y(n_7559)
);

INVx1_ASAP7_75t_L g7560 ( 
.A(n_7558),
.Y(n_7560)
);

INVx2_ASAP7_75t_SL g7561 ( 
.A(n_7559),
.Y(n_7561)
);

AOI21xp5_ASAP7_75t_L g7562 ( 
.A1(n_7561),
.A2(n_7544),
.B(n_7533),
.Y(n_7562)
);

OA21x2_ASAP7_75t_L g7563 ( 
.A1(n_7562),
.A2(n_7560),
.B(n_7545),
.Y(n_7563)
);

HB1xp67_ASAP7_75t_L g7564 ( 
.A(n_7563),
.Y(n_7564)
);

AOI21xp5_ASAP7_75t_L g7565 ( 
.A1(n_7564),
.A2(n_7547),
.B(n_7534),
.Y(n_7565)
);

AOI21xp5_ASAP7_75t_L g7566 ( 
.A1(n_7565),
.A2(n_864),
.B(n_865),
.Y(n_7566)
);

NAND3xp33_ASAP7_75t_L g7567 ( 
.A(n_7566),
.B(n_864),
.C(n_865),
.Y(n_7567)
);

AOI322xp5_ASAP7_75t_L g7568 ( 
.A1(n_7567),
.A2(n_864),
.A3(n_866),
.B1(n_867),
.B2(n_868),
.C1(n_869),
.C2(n_870),
.Y(n_7568)
);

OAI221xp5_ASAP7_75t_R g7569 ( 
.A1(n_7568),
.A2(n_866),
.B1(n_867),
.B2(n_868),
.C(n_869),
.Y(n_7569)
);

AOI22xp5_ASAP7_75t_L g7570 ( 
.A1(n_7569),
.A2(n_870),
.B1(n_867),
.B2(n_868),
.Y(n_7570)
);

AOI211xp5_ASAP7_75t_L g7571 ( 
.A1(n_7570),
.A2(n_873),
.B(n_870),
.C(n_871),
.Y(n_7571)
);


endmodule