module fake_jpeg_31565_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_70),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_2),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_76),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_52),
.B(n_58),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_45),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_58),
.B(n_53),
.C(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_89),
.B1(n_10),
.B2(n_13),
.Y(n_122)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_75),
.B1(n_56),
.B2(n_45),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_60),
.C(n_57),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_95),
.C(n_2),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_50),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_47),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_97),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_110),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_7),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_8),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_121),
.B(n_16),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_42),
.B1(n_28),
.B2(n_12),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_18),
.B(n_19),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_9),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_14),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_9),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_10),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_130),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_15),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_133),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_122),
.C(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_134),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_118),
.B1(n_113),
.B2(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_113),
.B(n_24),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_139),
.A2(n_125),
.B(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_126),
.C(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_131),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_136),
.B1(n_140),
.B2(n_139),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_126),
.C(n_142),
.Y(n_149)
);

AOI322xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_146),
.A3(n_141),
.B1(n_125),
.B2(n_135),
.C1(n_32),
.C2(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_25),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_30),
.A3(n_31),
.B1(n_34),
.B2(n_35),
.C1(n_36),
.C2(n_37),
.Y(n_153)
);


endmodule