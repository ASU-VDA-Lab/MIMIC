module fake_jpeg_8940_n_92 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_92);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_22),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_15),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_15),
.C(n_25),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_22),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_20),
.B1(n_15),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_20),
.B2(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_20),
.B1(n_19),
.B2(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_45),
.B1(n_14),
.B2(n_11),
.Y(n_55)
);

OAI22x1_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_25),
.B1(n_33),
.B2(n_10),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_33),
.C(n_23),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_49),
.C(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_26),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_30),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_58),
.B1(n_10),
.B2(n_16),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_57),
.B(n_13),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_18),
.B1(n_13),
.B2(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_46),
.C(n_18),
.Y(n_65)
);

XNOR2x1_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.C(n_68),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_16),
.B(n_4),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_54),
.A3(n_56),
.B1(n_61),
.B2(n_16),
.C(n_8),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_1),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_16),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_67),
.C(n_4),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_3),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_76),
.C(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_5),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_73),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_82),
.B1(n_81),
.B2(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_90),
.Y(n_92)
);


endmodule