module fake_aes_9806_n_613 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_613);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_613;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_384;
wire n_434;
wire n_227;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_54), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_22), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_25), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_2), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_56), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_27), .Y(n_82) );
INVx3_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
INVx3_ASAP7_75t_L g84 ( .A(n_66), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_38), .Y(n_85) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_23), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_76), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_72), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_21), .Y(n_90) );
BUFx2_ASAP7_75t_L g91 ( .A(n_63), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_61), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_50), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_73), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_59), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_0), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_47), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_35), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_52), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_4), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_33), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_14), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_36), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_18), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_19), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_65), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_45), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_5), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_12), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_43), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_24), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_92), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_91), .B(n_0), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_84), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_91), .B(n_1), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_83), .B(n_1), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_116), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_93), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_86), .B(n_3), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
NOR2x1_ASAP7_75t_L g137 ( .A(n_78), .B(n_3), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_90), .B(n_4), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_90), .B(n_5), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_117), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_96), .B(n_6), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_78), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_88), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_96), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_79), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_103), .B(n_6), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_101), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_113), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_82), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_113), .B(n_7), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_146), .B(n_103), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_122), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_146), .B(n_106), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_120), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_122), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_123), .A2(n_106), .B1(n_108), .B2(n_109), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_123), .B(n_114), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_130), .B(n_114), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_122), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_138), .B(n_108), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_127), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_138), .B(n_85), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_127), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_130), .A2(n_109), .B1(n_111), .B2(n_112), .Y(n_184) );
INVx8_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_127), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_142), .B(n_104), .Y(n_187) );
BUFx2_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_128), .B(n_111), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_142), .B(n_100), .Y(n_192) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_127), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_145), .B(n_87), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_143), .B(n_144), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_121), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_185), .A2(n_149), .B1(n_139), .B2(n_153), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_173), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_188), .B(n_139), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_164), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_178), .B(n_139), .Y(n_206) );
AND3x1_ASAP7_75t_L g207 ( .A(n_184), .B(n_135), .C(n_125), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_166), .Y(n_208) );
BUFx12f_ASAP7_75t_SL g209 ( .A(n_156), .Y(n_209) );
BUFx4f_ASAP7_75t_L g210 ( .A(n_185), .Y(n_210) );
INVxp67_ASAP7_75t_SL g211 ( .A(n_182), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_197), .B(n_143), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_195), .B(n_144), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_178), .A2(n_149), .B1(n_154), .B2(n_153), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_195), .B(n_147), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_188), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_185), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_195), .B(n_147), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_197), .B(n_154), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_194), .B(n_149), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_178), .B(n_149), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_194), .B(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_156), .B(n_141), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_185), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_178), .B(n_137), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_162), .Y(n_228) );
AND2x6_ASAP7_75t_SL g229 ( .A(n_156), .B(n_155), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_170), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_161), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_163), .B(n_136), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_162), .B(n_119), .Y(n_233) );
BUFx4f_ASAP7_75t_L g234 ( .A(n_185), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_163), .B(n_136), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_161), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_175), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_163), .B(n_136), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_178), .B(n_134), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_175), .Y(n_241) );
NAND2x1p5_ASAP7_75t_L g242 ( .A(n_162), .B(n_126), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_177), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_177), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_191), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_191), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_174), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_185), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_196), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
INVx5_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_226), .A2(n_162), .B1(n_165), .B2(n_182), .Y(n_252) );
AOI21xp33_ASAP7_75t_L g253 ( .A1(n_248), .A2(n_174), .B(n_190), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_225), .B(n_165), .Y(n_254) );
NAND3xp33_ASAP7_75t_L g255 ( .A(n_207), .B(n_184), .C(n_190), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_221), .A2(n_165), .B(n_182), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_218), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_211), .A2(n_182), .B1(n_165), .B2(n_187), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_224), .B(n_190), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_201), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_207), .B(n_168), .C(n_165), .Y(n_262) );
CKINVDCx11_ASAP7_75t_R g263 ( .A(n_204), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_225), .B(n_187), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_225), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_218), .B(n_137), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_210), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_248), .B(n_192), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_241), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_201), .Y(n_271) );
NAND2xp33_ASAP7_75t_L g272 ( .A(n_198), .B(n_131), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_210), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_210), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_206), .A2(n_192), .B1(n_168), .B2(n_171), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_214), .A2(n_171), .B(n_172), .C(n_134), .Y(n_277) );
BUFx2_ASAP7_75t_SL g278 ( .A(n_206), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_241), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_247), .B(n_172), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_231), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_226), .B(n_102), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_234), .A2(n_151), .B1(n_94), .B2(n_95), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_234), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_244), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_234), .B(n_193), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_203), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_244), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_199), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_199), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_205), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_199), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_214), .A2(n_151), .B1(n_94), .B2(n_95), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_205), .Y(n_294) );
AOI21xp33_ASAP7_75t_L g295 ( .A1(n_212), .A2(n_193), .B(n_89), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_209), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_199), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_228), .Y(n_298) );
CKINVDCx6p67_ASAP7_75t_R g299 ( .A(n_251), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_255), .A2(n_209), .B1(n_237), .B2(n_226), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_276), .A2(n_213), .B1(n_219), .B2(n_216), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_280), .B(n_220), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_260), .A2(n_232), .B1(n_239), .B2(n_235), .C(n_223), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_262), .A2(n_226), .B1(n_206), .B2(n_222), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_280), .B(n_206), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_281), .A2(n_222), .B1(n_202), .B2(n_228), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_276), .A2(n_238), .B1(n_208), .B2(n_246), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_281), .A2(n_222), .B1(n_228), .B2(n_246), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_253), .A2(n_222), .B1(n_228), .B2(n_245), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_269), .B(n_208), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_258), .B(n_215), .Y(n_313) );
AOI222xp33_ASAP7_75t_L g314 ( .A1(n_272), .A2(n_238), .B1(n_215), .B2(n_245), .C1(n_243), .C2(n_230), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_272), .A2(n_243), .B1(n_230), .B2(n_250), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_279), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_265), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_282), .A2(n_250), .B1(n_249), .B2(n_240), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g319 ( .A1(n_278), .A2(n_249), .B1(n_229), .B2(n_133), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_261), .B(n_229), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_251), .B(n_242), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_261), .A2(n_151), .B1(n_133), .B2(n_242), .Y(n_322) );
OAI222xp33_ASAP7_75t_L g323 ( .A1(n_293), .A2(n_105), .B1(n_97), .B2(n_118), .C1(n_115), .C2(n_110), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_251), .B(n_268), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_271), .Y(n_325) );
BUFx12f_ASAP7_75t_L g326 ( .A(n_263), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_271), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_273), .B(n_242), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_279), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_251), .A2(n_233), .B1(n_133), .B2(n_97), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_273), .Y(n_331) );
BUFx4f_ASAP7_75t_SL g332 ( .A(n_296), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g333 ( .A1(n_304), .A2(n_277), .B1(n_283), .B2(n_259), .C(n_252), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_302), .A2(n_266), .B1(n_282), .B2(n_278), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_325), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_320), .B(n_296), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_320), .A2(n_259), .B1(n_265), .B2(n_251), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_303), .B(n_312), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_302), .A2(n_266), .B1(n_282), .B2(n_269), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_304), .A2(n_266), .B1(n_269), .B2(n_287), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_303), .B(n_291), .Y(n_341) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_309), .A2(n_322), .B(n_328), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_314), .A2(n_287), .B1(n_295), .B2(n_291), .Y(n_343) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_309), .B(n_294), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_301), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_315), .A2(n_319), .B1(n_317), .B2(n_318), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
OR2x2_ASAP7_75t_SL g348 ( .A(n_313), .B(n_294), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_313), .B(n_285), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_300), .A2(n_256), .B1(n_264), .B2(n_284), .C(n_274), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_314), .A2(n_288), .B1(n_285), .B2(n_257), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_319), .A2(n_267), .B1(n_297), .B2(n_290), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
AND2x6_ASAP7_75t_SL g355 ( .A(n_326), .B(n_254), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_315), .A2(n_305), .B1(n_312), .B2(n_306), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_306), .A2(n_267), .B1(n_297), .B2(n_290), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_325), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_311), .A2(n_297), .B1(n_289), .B2(n_257), .Y(n_360) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_358), .B(n_299), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_341), .B(n_301), .Y(n_362) );
OAI21x1_ASAP7_75t_L g363 ( .A1(n_344), .A2(n_322), .B(n_329), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_335), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_333), .A2(n_323), .B(n_328), .Y(n_365) );
OAI321xp33_ASAP7_75t_L g366 ( .A1(n_346), .A2(n_310), .A3(n_89), .B1(n_100), .B2(n_118), .C(n_107), .Y(n_366) );
OA222x2_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_348), .B1(n_349), .B2(n_335), .C1(n_359), .C2(n_355), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_339), .A2(n_334), .B1(n_340), .B2(n_336), .C(n_308), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_359), .Y(n_369) );
OAI31xp33_ASAP7_75t_L g370 ( .A1(n_333), .A2(n_323), .A3(n_331), .B(n_327), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_338), .A2(n_327), .B1(n_331), .B2(n_330), .C(n_110), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_344), .A2(n_329), .B(n_316), .Y(n_373) );
NAND3xp33_ASAP7_75t_SL g374 ( .A(n_354), .B(n_104), .C(n_99), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_345), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_338), .A2(n_99), .B1(n_105), .B2(n_107), .C(n_115), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_341), .B(n_332), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_345), .B(n_307), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_352), .A2(n_329), .B1(n_307), .B2(n_316), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_347), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_355), .B(n_326), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_342), .A2(n_321), .B(n_316), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_324), .B1(n_307), .B2(n_288), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_343), .A2(n_264), .B1(n_275), .B2(n_289), .C(n_98), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_351), .B(n_324), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_352), .A2(n_264), .B1(n_275), .B2(n_98), .C(n_274), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_370), .B(n_376), .C(n_381), .D(n_385), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_383), .B(n_354), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_389), .A2(n_348), .B1(n_353), .B2(n_337), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_362), .B(n_342), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_391), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_362), .B(n_342), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_364), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_387), .Y(n_403) );
OAI211xp5_ASAP7_75t_SL g404 ( .A1(n_377), .A2(n_357), .B(n_360), .C(n_350), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_371), .B(n_342), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_387), .B(n_358), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_371), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_375), .B(n_358), .Y(n_409) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_366), .B(n_268), .C(n_326), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_380), .B(n_358), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_366), .B(n_324), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_380), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_368), .A2(n_324), .B1(n_268), .B2(n_254), .Y(n_415) );
AOI33xp33_ASAP7_75t_L g416 ( .A1(n_367), .A2(n_7), .A3(n_8), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_370), .A2(n_148), .B1(n_150), .B2(n_152), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_365), .A2(n_148), .B1(n_150), .B2(n_152), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_374), .B(n_286), .C(n_181), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_390), .B(n_148), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_148), .B1(n_150), .B2(n_152), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_390), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
AO221x2_ASAP7_75t_L g425 ( .A1(n_367), .A2(n_8), .B1(n_9), .B2(n_10), .C(n_11), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_384), .B(n_148), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_388), .B(n_148), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_386), .A2(n_254), .A3(n_14), .B(n_15), .Y(n_429) );
OAI33xp33_ASAP7_75t_L g430 ( .A1(n_379), .A2(n_13), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_361), .A2(n_387), .A3(n_372), .B(n_17), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_382), .B(n_152), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_402), .B(n_373), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_392), .A2(n_150), .B1(n_152), .B2(n_169), .C(n_181), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_396), .B(n_405), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_396), .B(n_373), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_419), .B(n_363), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_405), .B(n_363), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_398), .B(n_152), .Y(n_443) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_400), .A2(n_13), .A3(n_16), .B1(n_19), .B2(n_20), .B3(n_21), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_397), .B(n_150), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
NAND3xp33_ASAP7_75t_SL g447 ( .A(n_416), .B(n_20), .C(n_189), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_401), .Y(n_449) );
AO21x1_ASAP7_75t_L g450 ( .A1(n_432), .A2(n_189), .B(n_183), .Y(n_450) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_430), .B(n_181), .C(n_169), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_393), .B(n_150), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_413), .A2(n_193), .B(n_292), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_409), .B(n_28), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_409), .B(n_30), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_423), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_412), .B(n_31), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_412), .B(n_32), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_431), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_425), .B(n_180), .C(n_158), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_432), .B(n_298), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_424), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_403), .B(n_34), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_403), .B(n_37), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_401), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_401), .B(n_298), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_426), .B(n_39), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_429), .B(n_183), .C(n_167), .D(n_179), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_421), .B(n_41), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_421), .B(n_42), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_427), .B(n_44), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_395), .B(n_298), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_395), .B(n_51), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_428), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_407), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_395), .B(n_176), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_395), .B(n_298), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_463), .A2(n_410), .B1(n_429), .B2(n_415), .C(n_394), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_437), .B(n_443), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_478), .A2(n_415), .B(n_407), .C(n_425), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_437), .B(n_425), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_480), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_438), .B(n_425), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_443), .B(n_417), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_444), .A2(n_404), .B1(n_418), .B2(n_422), .C(n_420), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_476), .B(n_53), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_449), .Y(n_495) );
OAI31xp33_ASAP7_75t_L g496 ( .A1(n_478), .A2(n_468), .A3(n_466), .B(n_467), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_466), .A2(n_183), .A3(n_179), .B(n_176), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_452), .B(n_158), .C(n_186), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_438), .B(n_55), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_447), .A2(n_193), .B(n_167), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_442), .B(n_57), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_457), .B(n_58), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_448), .B(n_167), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_454), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_476), .B(n_62), .Y(n_507) );
AOI211xp5_ASAP7_75t_L g508 ( .A1(n_450), .A2(n_186), .B(n_180), .C(n_159), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_446), .A2(n_169), .B1(n_181), .B2(n_186), .C(n_180), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_464), .A2(n_64), .B(n_67), .C(n_68), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_457), .B(n_70), .Y(n_511) );
OAI211xp5_ASAP7_75t_L g512 ( .A1(n_445), .A2(n_179), .B(n_186), .C(n_180), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_458), .B(n_71), .Y(n_513) );
OAI21xp5_ASAP7_75t_SL g514 ( .A1(n_467), .A2(n_459), .B(n_460), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_461), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_455), .B(n_456), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_74), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_434), .B(n_75), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_435), .A2(n_193), .B1(n_158), .B2(n_159), .C(n_157), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_459), .B(n_181), .Y(n_520) );
BUFx12f_ASAP7_75t_L g521 ( .A(n_459), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_456), .B(n_169), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_462), .B(n_157), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_460), .B(n_157), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_489), .A2(n_450), .B1(n_440), .B2(n_473), .C(n_465), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_490), .B(n_434), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_521), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_491), .B(n_473), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_485), .B(n_479), .Y(n_530) );
NOR2xp33_ASAP7_75t_R g531 ( .A(n_495), .B(n_482), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_505), .B(n_479), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_515), .B(n_525), .Y(n_533) );
NAND4xp25_ASAP7_75t_SL g534 ( .A(n_486), .B(n_453), .C(n_472), .D(n_474), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_516), .B(n_470), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_483), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_487), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_496), .B(n_477), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_488), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_497), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_508), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_514), .A2(n_481), .B(n_469), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_484), .A2(n_481), .B(n_471), .C(n_451), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_500), .B(n_472), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_506), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_484), .B(n_475), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_500), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_502), .B(n_475), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_520), .A2(n_292), .B1(n_158), .B2(n_159), .Y(n_549) );
AND3x1_ASAP7_75t_L g550 ( .A(n_501), .B(n_236), .C(n_227), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_499), .B(n_157), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_518), .B(n_157), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_492), .B(n_157), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_492), .B(n_158), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_SL g555 ( .A1(n_501), .A2(n_200), .B(n_236), .C(n_227), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_512), .A2(n_292), .B(n_159), .Y(n_556) );
OAI211xp5_ASAP7_75t_L g557 ( .A1(n_493), .A2(n_158), .B(n_159), .C(n_180), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_522), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_524), .A2(n_159), .B1(n_180), .B2(n_186), .C(n_292), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_510), .A2(n_292), .B(n_180), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_523), .B(n_159), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_503), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_494), .A2(n_186), .B(n_200), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_498), .A2(n_186), .B(n_507), .C(n_519), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_519), .A2(n_509), .B(n_517), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_513), .A2(n_514), .B1(n_486), .B2(n_463), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_511), .A2(n_514), .B1(n_486), .B2(n_463), .Y(n_568) );
AOI222xp33_ASAP7_75t_L g569 ( .A1(n_504), .A2(n_489), .B1(n_491), .B2(n_484), .C1(n_444), .C2(n_447), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_491), .A2(n_425), .B1(n_489), .B2(n_514), .Y(n_570) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_515), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_495), .B(n_381), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_485), .B(n_437), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_490), .B(n_495), .Y(n_574) );
AO221x1_ASAP7_75t_L g575 ( .A1(n_567), .A2(n_568), .B1(n_528), .B2(n_531), .C(n_570), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_541), .A2(n_534), .B(n_538), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_526), .B(n_527), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_546), .A2(n_543), .B1(n_538), .B2(n_527), .C(n_542), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_541), .A2(n_557), .B(n_569), .C(n_528), .Y(n_579) );
AND3x1_ASAP7_75t_L g580 ( .A(n_528), .B(n_546), .C(n_572), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_573), .B(n_571), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_571), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
NAND4xp75_ASAP7_75t_L g584 ( .A(n_574), .B(n_550), .C(n_566), .D(n_529), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_574), .A2(n_558), .B1(n_547), .B2(n_535), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_531), .A2(n_544), .B1(n_548), .B2(n_562), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_537), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_533), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_532), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_579), .B(n_554), .C(n_553), .Y(n_590) );
OAI211xp5_ASAP7_75t_L g591 ( .A1(n_579), .A2(n_565), .B(n_564), .C(n_551), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_576), .A2(n_563), .B1(n_545), .B2(n_536), .C(n_540), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_584), .B(n_551), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_588), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_582), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_578), .B(n_539), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_578), .B(n_555), .C(n_559), .D(n_549), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_587), .Y(n_598) );
AO22x2_ASAP7_75t_L g599 ( .A1(n_596), .A2(n_575), .B1(n_577), .B2(n_589), .Y(n_599) );
NAND5xp2_ASAP7_75t_L g600 ( .A(n_591), .B(n_586), .C(n_580), .D(n_585), .E(n_556), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_594), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_593), .B(n_552), .C(n_561), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_590), .B(n_583), .Y(n_603) );
NAND5xp2_ASAP7_75t_L g604 ( .A(n_599), .B(n_592), .C(n_597), .D(n_598), .E(n_560), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_601), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_603), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_606), .A2(n_599), .B1(n_595), .B2(n_600), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_604), .B(n_602), .C(n_581), .Y(n_608) );
XOR2xp5_ASAP7_75t_L g609 ( .A(n_607), .B(n_605), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_608), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_610), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_611), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_612), .A2(n_609), .B(n_605), .Y(n_613) );
endmodule