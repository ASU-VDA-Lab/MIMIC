module fake_jpeg_5405_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_7),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_18),
.B(n_26),
.C(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_54),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_21),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_44),
.B(n_18),
.C(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_20),
.B1(n_36),
.B2(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_57),
.B1(n_68),
.B2(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_31),
.B1(n_32),
.B2(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_31),
.B1(n_32),
.B2(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_20),
.B1(n_23),
.B2(n_32),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_83),
.B1(n_96),
.B2(n_54),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_23),
.B1(n_20),
.B2(n_36),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_91),
.B1(n_65),
.B2(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_86),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_58),
.B1(n_55),
.B2(n_66),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_60),
.B(n_59),
.C(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_65),
.B1(n_50),
.B2(n_70),
.Y(n_103)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_23),
.B1(n_20),
.B2(n_44),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_26),
.C(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_100),
.B1(n_102),
.B2(n_104),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_114),
.B1(n_77),
.B2(n_84),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_49),
.B1(n_50),
.B2(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_73),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_50),
.B1(n_52),
.B2(n_46),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_53),
.B1(n_65),
.B2(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_113),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_41),
.B1(n_19),
.B2(n_28),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_112),
.B1(n_117),
.B2(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_119),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_78),
.B1(n_72),
.B2(n_86),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_41),
.B1(n_25),
.B2(n_27),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_28),
.B(n_34),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_77),
.C(n_81),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_56),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_95),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_80),
.B1(n_90),
.B2(n_94),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_41),
.B1(n_24),
.B2(n_64),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_76),
.B1(n_84),
.B2(n_64),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_76),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_101),
.C(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_133),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_139),
.B(n_142),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_138),
.B1(n_146),
.B2(n_141),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_81),
.C(n_73),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_33),
.Y(n_178)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_34),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_0),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_147),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_56),
.C(n_24),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_0),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_0),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_106),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_124),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_148),
.B(n_129),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_175),
.C(n_140),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_103),
.B(n_99),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_143),
.B(n_132),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_98),
.B1(n_104),
.B2(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_112),
.C(n_117),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_173),
.B1(n_177),
.B2(n_182),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_134),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_178),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_113),
.B1(n_110),
.B2(n_56),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_174),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_24),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_24),
.B1(n_33),
.B2(n_111),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_1),
.Y(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_188),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_190),
.B(n_136),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_194),
.Y(n_214)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_144),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_129),
.C(n_128),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_200),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_128),
.C(n_147),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_158),
.C(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_164),
.B1(n_168),
.B2(n_158),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_217),
.B1(n_222),
.B2(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_216),
.C(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_167),
.C(n_170),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_170),
.B1(n_174),
.B2(n_160),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_181),
.B1(n_131),
.B2(n_153),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_154),
.C(n_172),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_229),
.C(n_200),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_172),
.C(n_163),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_149),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_192),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_153),
.B1(n_161),
.B2(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_145),
.C(n_111),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_231),
.C(n_225),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_145),
.C(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_189),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_191),
.B1(n_194),
.B2(n_203),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_247),
.C(n_242),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_250),
.B(n_252),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_184),
.B1(n_186),
.B2(n_189),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_254),
.B1(n_218),
.B2(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_245),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_216),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_229),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_255),
.Y(n_257)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_217),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_230),
.C(n_215),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_262),
.C(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_266),
.B1(n_243),
.B2(n_237),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_185),
.B1(n_202),
.B2(n_190),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_231),
.C(n_207),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_235),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_278),
.B1(n_10),
.B2(n_11),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_243),
.B1(n_236),
.B2(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_284),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_211),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_202),
.B(n_246),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_249),
.B(n_191),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_193),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_4),
.Y(n_290)
);

AOI321xp33_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_193),
.A3(n_10),
.B1(n_11),
.B2(n_5),
.C(n_6),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_290),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_262),
.B1(n_261),
.B2(n_260),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_294),
.C(n_279),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_5),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_7),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_297),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_279),
.C(n_272),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_302),
.B(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_11),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_286),
.A3(n_289),
.B1(n_15),
.B2(n_16),
.C1(n_13),
.C2(n_14),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_16),
.B(n_13),
.C(n_15),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_300),
.C(n_15),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_311),
.Y(n_313)
);

NOR3xp33_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_310),
.C(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_16),
.Y(n_315)
);


endmodule