module fake_jpeg_20367_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_48),
.B1(n_46),
.B2(n_58),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_70),
.B1(n_47),
.B2(n_73),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_49),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_50),
.B(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_65),
.B1(n_45),
.B2(n_56),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_74),
.B1(n_54),
.B2(n_53),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_0),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_47),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_120),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_25),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_62),
.B1(n_67),
.B2(n_71),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_138),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_72),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_131),
.B(n_20),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_132),
.B1(n_136),
.B2(n_9),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_63),
.B(n_1),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_61),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_137),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_115),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_144),
.B(n_147),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_26),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_131),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_146),
.B(n_151),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_139),
.C(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_130),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_36),
.Y(n_164)
);


endmodule