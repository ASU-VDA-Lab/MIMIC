module fake_jpeg_16608_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_17),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_27),
.B1(n_26),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_95)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_29),
.B1(n_23),
.B2(n_30),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_19),
.B(n_21),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_24),
.B(n_20),
.C(n_28),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_23),
.B1(n_21),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_21),
.B1(n_30),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_24),
.B1(n_31),
.B2(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_70),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_49),
.C(n_51),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_40),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_18),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_83),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_94),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_88),
.B(n_50),
.Y(n_112)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_40),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_43),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_22),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_22),
.B(n_20),
.C(n_17),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_43),
.A2(n_20),
.B1(n_25),
.B2(n_18),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_124)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_109),
.Y(n_135)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_43),
.B(n_50),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_112),
.B(n_96),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_53),
.B1(n_44),
.B2(n_52),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_77),
.B1(n_65),
.B2(n_75),
.Y(n_133)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_82),
.Y(n_127)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_136),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_95),
.C(n_80),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_104),
.C(n_107),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_82),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_87),
.B1(n_70),
.B2(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_140),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_88),
.B1(n_78),
.B2(n_64),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_93),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_118),
.B(n_110),
.C(n_122),
.D(n_103),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_78),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_147),
.B(n_149),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_32),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_145),
.C(n_26),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_32),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_150),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_65),
.B(n_77),
.C(n_66),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_14),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_121),
.B1(n_107),
.B2(n_102),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_154),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_134),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_161),
.C(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_106),
.C(n_99),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_143),
.B1(n_138),
.B2(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_171),
.B1(n_2),
.B2(n_4),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_145),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_106),
.C(n_99),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_67),
.B1(n_100),
.B2(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_26),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_176),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

OR2x6_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_143),
.Y(n_178)
);

NAND2x1_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_164),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_181),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_147),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_159),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_67),
.B1(n_129),
.B2(n_3),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_185),
.B1(n_188),
.B2(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_173),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_156),
.C(n_157),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_194),
.C(n_199),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_161),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_193),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_192),
.B1(n_198),
.B2(n_201),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_165),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_158),
.B(n_168),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_155),
.B1(n_6),
.B2(n_7),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_208),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_174),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_177),
.B1(n_175),
.B2(n_186),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_194),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.C(n_199),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_198),
.C(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_214),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_193),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_205),
.B(n_191),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

AOI31xp67_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_206),
.A3(n_210),
.B(n_211),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_219),
.A2(n_220),
.B(n_221),
.C(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_213),
.B(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_10),
.B(n_226),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_10),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_228),
.Y(n_229)
);


endmodule