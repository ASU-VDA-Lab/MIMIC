module fake_jpeg_21526_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_22),
.B1(n_17),
.B2(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_38),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_24),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_17),
.B1(n_22),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_30),
.B1(n_19),
.B2(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_55),
.A2(n_78),
.B1(n_48),
.B2(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_68),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_69),
.B(n_25),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_23),
.B1(n_30),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_44),
.B1(n_43),
.B2(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_80),
.B1(n_46),
.B2(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_19),
.B1(n_26),
.B2(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_39),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_52),
.B(n_44),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_38),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_103),
.B1(n_107),
.B2(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_108),
.B1(n_82),
.B2(n_73),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_34),
.C(n_39),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_70),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_77),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_58),
.C(n_61),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_80),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_105),
.B1(n_82),
.B2(n_75),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_41),
.B1(n_48),
.B2(n_19),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_44),
.B1(n_52),
.B2(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_26),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_62),
.B1(n_57),
.B2(n_63),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_115),
.B1(n_119),
.B2(n_127),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_111),
.B(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_134),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_94),
.B1(n_86),
.B2(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_92),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_122),
.B(n_87),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_70),
.B1(n_66),
.B2(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_70),
.B1(n_66),
.B2(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_101),
.A3(n_92),
.B1(n_88),
.B2(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_70),
.B1(n_83),
.B2(n_67),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_136),
.B1(n_135),
.B2(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_34),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_15),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_15),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_101),
.C(n_94),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_28),
.C(n_21),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_145),
.A2(n_147),
.B(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_122),
.B(n_126),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_110),
.B1(n_91),
.B2(n_59),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_125),
.B1(n_23),
.B2(n_24),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_103),
.B1(n_108),
.B2(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_152),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_108),
.B1(n_93),
.B2(n_110),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_104),
.B(n_16),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_104),
.A3(n_31),
.B1(n_20),
.B2(n_27),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_21),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_100),
.B(n_26),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_130),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_31),
.B(n_27),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_169),
.B(n_5),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_85),
.B1(n_31),
.B2(n_27),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_170),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_85),
.B1(n_29),
.B2(n_25),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_168),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_85),
.B1(n_24),
.B2(n_21),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_116),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_175),
.B(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_176),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_139),
.B1(n_123),
.B2(n_133),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_124),
.A3(n_125),
.B1(n_120),
.B2(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_192),
.C(n_160),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_194),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_28),
.B1(n_15),
.B2(n_23),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_15),
.A3(n_28),
.B1(n_23),
.B2(n_14),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_187),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_14),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_193),
.B1(n_196),
.B2(n_198),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_143),
.C(n_150),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_159),
.B(n_3),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_6),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_144),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_159),
.B1(n_167),
.B2(n_157),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_162),
.B1(n_144),
.B2(n_157),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_161),
.B(n_145),
.Y(n_210)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_200),
.A2(n_166),
.B1(n_7),
.B2(n_8),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_208),
.C(n_219),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_146),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_206),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_221),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_146),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_155),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_167),
.B1(n_158),
.B2(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_216),
.B1(n_186),
.B2(n_178),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_152),
.B1(n_150),
.B2(n_156),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_181),
.B1(n_197),
.B2(n_177),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_8),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_8),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_227),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_207),
.B(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_184),
.B1(n_175),
.B2(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_175),
.B1(n_185),
.B2(n_199),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_175),
.B1(n_190),
.B2(n_188),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_187),
.B(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_239),
.B(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_204),
.C(n_201),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_246),
.C(n_248),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_220),
.C(n_208),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_219),
.C(n_221),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_210),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_227),
.C(n_231),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_214),
.B(n_202),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_226),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_262),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_211),
.B1(n_217),
.B2(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_248),
.C(n_245),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_229),
.B1(n_230),
.B2(n_202),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_233),
.C(n_211),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_263),
.C(n_265),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.C(n_193),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_249),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_274),
.B1(n_250),
.B2(n_171),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_252),
.B1(n_254),
.B2(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_243),
.C(n_251),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_253),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_257),
.B(n_243),
.Y(n_278)
);

AOI21x1_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_280),
.B(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_191),
.C(n_183),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_196),
.C(n_10),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_9),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_9),
.C(n_10),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_269),
.B(n_11),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_284),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_280),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_287),
.B(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_10),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_293),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_12),
.B(n_13),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_12),
.C(n_13),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_12),
.B(n_282),
.Y(n_300)
);


endmodule