module fake_jpeg_14846_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_54),
.Y(n_74)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_64),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_26),
.C(n_30),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_26),
.C(n_17),
.Y(n_72)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_33),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_43),
.B1(n_38),
.B2(n_23),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_42),
.B1(n_43),
.B2(n_23),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_42),
.B1(n_16),
.B2(n_25),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_42),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_58),
.C(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_49),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_102),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_75),
.B1(n_87),
.B2(n_69),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_115),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_103),
.C(n_107),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_48),
.B1(n_51),
.B2(n_44),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_114),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_71),
.Y(n_102)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_57),
.B1(n_50),
.B2(n_47),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_58),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_57),
.B1(n_66),
.B2(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_50),
.B1(n_47),
.B2(n_45),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_86),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_33),
.B1(n_25),
.B2(n_20),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_26),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_59),
.B(n_0),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_18),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_135),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_85),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_74),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_74),
.B1(n_67),
.B2(n_73),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_113),
.B1(n_111),
.B2(n_38),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_R g133 ( 
.A(n_116),
.B(n_73),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_21),
.B(n_30),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_70),
.B1(n_81),
.B2(n_80),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_10),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_140),
.A2(n_141),
.B(n_18),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_8),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_127),
.C(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_98),
.C(n_86),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_167),
.C(n_120),
.Y(n_175)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_80),
.B1(n_105),
.B2(n_70),
.Y(n_148)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_79),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_157),
.B(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_172),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_121),
.B(n_125),
.C(n_122),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_161),
.B(n_2),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_113),
.B1(n_93),
.B2(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_93),
.B1(n_38),
.B2(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_0),
.Y(n_159)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_82),
.B(n_21),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_82),
.C(n_24),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_21),
.B(n_24),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_121),
.B(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_31),
.B1(n_27),
.B2(n_17),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_166),
.C(n_164),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_186),
.B(n_191),
.Y(n_219)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_195),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_123),
.B(n_129),
.C(n_140),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_193),
.B(n_197),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_161),
.B(n_21),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_189),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_1),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_31),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_199),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_165),
.B1(n_162),
.B2(n_152),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_157),
.B1(n_155),
.B2(n_147),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_158),
.B1(n_154),
.B2(n_148),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_224),
.B(n_191),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_151),
.C(n_149),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_168),
.C(n_153),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_154),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_167),
.C(n_156),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_172),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_184),
.C(n_176),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_170),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_199),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_200),
.B1(n_180),
.B2(n_193),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_235),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_230),
.C(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_193),
.B1(n_178),
.B2(n_186),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_178),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_185),
.B(n_187),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_219),
.B(n_205),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_188),
.C(n_182),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_188),
.C(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_230),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_228),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_214),
.C(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_257),
.C(n_258),
.Y(n_264)
);

XNOR2x2_ASAP7_75t_SL g252 ( 
.A(n_234),
.B(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_207),
.C(n_212),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_219),
.C(n_220),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_209),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_239),
.CI(n_244),
.CON(n_266),
.SN(n_266)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_268),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_221),
.B(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_236),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_227),
.C(n_235),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_247),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_274),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_254),
.B(n_203),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_281),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_262),
.B1(n_255),
.B2(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.C(n_286),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_249),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_177),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_4),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_9),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_264),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_283),
.C(n_284),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_288),
.A2(n_265),
.B(n_266),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_11),
.B(n_12),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_295),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_275),
.C(n_10),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_9),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_15),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_301),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_9),
.B(n_10),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_12),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_297),
.B(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_309),
.A2(n_307),
.B(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_306),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_13),
.B(n_15),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_312),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_13),
.Y(n_314)
);


endmodule