module real_jpeg_17555_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AO22x1_ASAP7_75t_SL g14 ( 
.A1(n_0),
.A2(n_5),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_3),
.B1(n_16),
.B2(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_29),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_12),
.B(n_21),
.Y(n_7)
);

INVx1_ASAP7_75t_SL g8 ( 
.A(n_9),
.Y(n_8)
);

AND2x4_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

OR2x4_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_17),
.B(n_18),
.Y(n_13)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_19),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);


endmodule