module fake_aes_4939_n_473 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_473);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_473;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g72 ( .A(n_36), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_52), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_39), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_56), .Y(n_75) );
INVxp33_ASAP7_75t_SL g76 ( .A(n_23), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_4), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_43), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_8), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_31), .Y(n_80) );
INVx1_ASAP7_75t_SL g81 ( .A(n_54), .Y(n_81) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_12), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_20), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_68), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_11), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_42), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_28), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_8), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_47), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_4), .Y(n_92) );
INVxp33_ASAP7_75t_L g93 ( .A(n_33), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_21), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_45), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_18), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_37), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_35), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_71), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_67), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_51), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g104 ( .A(n_94), .B(n_0), .Y(n_104) );
INVx3_ASAP7_75t_L g105 ( .A(n_82), .Y(n_105) );
NAND2x1_ASAP7_75t_L g106 ( .A(n_82), .B(n_0), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_94), .B(n_1), .Y(n_107) );
BUFx8_ASAP7_75t_L g108 ( .A(n_94), .Y(n_108) );
NOR2x1_ASAP7_75t_L g109 ( .A(n_72), .B(n_1), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_89), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_103), .B(n_2), .Y(n_113) );
NOR2x1_ASAP7_75t_L g114 ( .A(n_74), .B(n_75), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_86), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_94), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
INVx4_ASAP7_75t_L g118 ( .A(n_94), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_95), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_80), .B(n_2), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_93), .B(n_3), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
BUFx8_ASAP7_75t_SL g123 ( .A(n_110), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_115), .B(n_93), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_120), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_108), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_108), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_112), .B(n_86), .Y(n_131) );
INVx2_ASAP7_75t_SL g132 ( .A(n_108), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_116), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_116), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_114), .B(n_77), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_113), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_118), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_120), .B(n_83), .Y(n_143) );
INVx2_ASAP7_75t_SL g144 ( .A(n_114), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_106), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_131), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_127), .B(n_121), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_134), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_123), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_134), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_140), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_134), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_125), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
AND3x1_ASAP7_75t_L g157 ( .A(n_124), .B(n_109), .C(n_79), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_144), .B(n_76), .Y(n_158) );
INVx3_ASAP7_75t_SL g159 ( .A(n_129), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_143), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_127), .Y(n_161) );
BUFx12f_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
HB1xp67_ASAP7_75t_SL g163 ( .A(n_130), .Y(n_163) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_125), .B(n_84), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_131), .B(n_111), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_141), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_150), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_128), .B(n_145), .C(n_136), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_152), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_162), .B(n_132), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_146), .B(n_136), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_155), .A2(n_145), .B(n_136), .C(n_106), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_162), .Y(n_182) );
BUFx12f_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_159), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_146), .B(n_143), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_165), .Y(n_187) );
OR2x6_ASAP7_75t_L g188 ( .A(n_167), .B(n_160), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_167), .B(n_160), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_165), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_164), .A2(n_104), .B1(n_107), .B2(n_92), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_165), .B(n_87), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_163), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_160), .B(n_85), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_192), .B(n_171), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_187), .B(n_171), .Y(n_201) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_175), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_180), .A2(n_148), .B(n_158), .C(n_159), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_177), .A2(n_149), .B1(n_160), .B2(n_170), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_181), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_182), .B(n_170), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_179), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_186), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_195), .A2(n_169), .B1(n_161), .B2(n_154), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_181), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_178), .Y(n_211) );
AOI211xp5_ASAP7_75t_L g212 ( .A1(n_194), .A2(n_82), .B(n_111), .C(n_157), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_174), .A2(n_166), .B(n_156), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_185), .A2(n_156), .B1(n_166), .B2(n_169), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_185), .B(n_174), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_188), .A2(n_161), .B1(n_169), .B2(n_154), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_193), .A2(n_161), .B1(n_88), .B2(n_97), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_207), .Y(n_219) );
OAI211xp5_ASAP7_75t_L g220 ( .A1(n_212), .A2(n_180), .B(n_184), .C(n_173), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g221 ( .A(n_212), .B(n_199), .C(n_181), .Y(n_221) );
OAI211xp5_ASAP7_75t_L g222 ( .A1(n_218), .A2(n_173), .B(n_101), .C(n_99), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_202), .A2(n_198), .B1(n_178), .B2(n_197), .Y(n_223) );
BUFx4f_ASAP7_75t_SL g224 ( .A(n_206), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_210), .Y(n_225) );
OAI21xp33_ASAP7_75t_L g226 ( .A1(n_218), .A2(n_200), .B(n_213), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_210), .Y(n_227) );
INVx1_ASAP7_75t_SL g228 ( .A(n_201), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_210), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_215), .A2(n_188), .B1(n_191), .B2(n_176), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_207), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_200), .A2(n_198), .B1(n_197), .B2(n_196), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_214), .A2(n_191), .B1(n_188), .B2(n_176), .Y(n_233) );
AOI221xp5_ASAP7_75t_L g234 ( .A1(n_203), .A2(n_189), .B1(n_196), .B2(n_182), .C(n_102), .Y(n_234) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_210), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_201), .B(n_208), .Y(n_236) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_205), .B(n_216), .Y(n_237) );
NOR2x1_ASAP7_75t_SL g238 ( .A(n_230), .B(n_210), .Y(n_238) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_221), .A2(n_209), .B(n_216), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_228), .A2(n_236), .B1(n_233), .B2(n_224), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_228), .B(n_205), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_225), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_219), .B(n_211), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_219), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g245 ( .A(n_220), .B(n_119), .C(n_95), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_231), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_226), .B(n_217), .Y(n_247) );
OAI31xp33_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_91), .A3(n_96), .B(n_98), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_225), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_231), .B(n_211), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_227), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_227), .B(n_211), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_229), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_226), .A2(n_206), .B1(n_188), .B2(n_191), .Y(n_256) );
AOI21xp5_ASAP7_75t_SL g257 ( .A1(n_234), .A2(n_176), .B(n_191), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_244), .B(n_229), .Y(n_258) );
NOR3xp33_ASAP7_75t_SL g259 ( .A(n_248), .B(n_240), .C(n_88), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_246), .B(n_229), .Y(n_261) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_256), .B(n_232), .Y(n_262) );
BUFx6f_ASAP7_75t_SL g263 ( .A(n_253), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_246), .B(n_223), .Y(n_264) );
OAI31xp33_ASAP7_75t_L g265 ( .A1(n_248), .A2(n_100), .A3(n_81), .B(n_206), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_241), .B(n_235), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_249), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_249), .B(n_3), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_242), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_252), .B(n_5), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_241), .B(n_95), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_252), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_241), .B(n_95), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_243), .B(n_189), .Y(n_276) );
AOI33xp33_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_204), .A3(n_7), .B1(n_9), .B2(n_10), .B3(n_13), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_242), .B(n_6), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_243), .B(n_95), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_242), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_250), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_243), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_251), .B(n_7), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_245), .B(n_251), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_266), .B(n_250), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_266), .B(n_255), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_267), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_260), .B(n_255), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_283), .B(n_9), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_271), .B(n_255), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_263), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_283), .B(n_251), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_269), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_271), .B(n_238), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_273), .Y(n_299) );
AO221x1_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_238), .B1(n_257), .B2(n_245), .C(n_247), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_282), .B(n_253), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_284), .A2(n_237), .B(n_239), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_279), .B(n_253), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_275), .B(n_237), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_273), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_275), .B(n_237), .Y(n_306) );
OR2x4_ASAP7_75t_L g307 ( .A(n_268), .B(n_119), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_274), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_280), .B(n_237), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_258), .B(n_253), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_269), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_268), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_258), .B(n_239), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_270), .Y(n_315) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_265), .B(n_183), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_280), .B(n_237), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_278), .B(n_239), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_281), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_285), .B(n_119), .Y(n_323) );
OAI31xp33_ASAP7_75t_L g324 ( .A1(n_264), .A2(n_105), .A3(n_117), .B(n_122), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_262), .B(n_10), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_312), .B(n_262), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_314), .B(n_285), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_314), .B(n_276), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_298), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_315), .B(n_277), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_323), .B(n_263), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_310), .B(n_259), .Y(n_336) );
NAND2xp67_ASAP7_75t_L g337 ( .A(n_325), .B(n_263), .Y(n_337) );
AOI21xp33_ASAP7_75t_L g338 ( .A1(n_291), .A2(n_90), .B(n_97), .Y(n_338) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_317), .A2(n_105), .A3(n_117), .B1(n_122), .B2(n_13), .C1(n_14), .C2(n_90), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_316), .B(n_118), .C(n_105), .D(n_122), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_290), .B(n_14), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_310), .B(n_118), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_310), .B(n_118), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_296), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_311), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_293), .B(n_199), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g347 ( .A(n_323), .B(n_139), .C(n_135), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_286), .B(n_287), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_286), .B(n_16), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_294), .B(n_17), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_287), .B(n_19), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_308), .B(n_22), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_307), .B(n_24), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_321), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_297), .B(n_25), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_319), .B(n_26), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_300), .A2(n_183), .B1(n_182), .B2(n_176), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_297), .B(n_199), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_301), .B(n_27), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_292), .B(n_289), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_313), .B(n_29), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_289), .B(n_292), .Y(n_365) );
NAND2xp33_ASAP7_75t_R g366 ( .A(n_293), .B(n_30), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_303), .B(n_32), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_307), .B(n_34), .Y(n_368) );
NAND3xp33_ASAP7_75t_L g369 ( .A(n_324), .B(n_302), .C(n_320), .Y(n_369) );
NOR2xp33_ASAP7_75t_R g370 ( .A(n_300), .B(n_38), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_366), .A2(n_313), .B1(n_306), .B2(n_304), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_346), .A2(n_306), .B(n_304), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_330), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_362), .B(n_313), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_335), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_326), .B(n_318), .Y(n_377) );
OAI21xp5_ASAP7_75t_SL g378 ( .A1(n_359), .A2(n_309), .B(n_318), .Y(n_378) );
NOR3xp33_ASAP7_75t_L g379 ( .A(n_369), .B(n_309), .C(n_139), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_348), .B(n_40), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_334), .B(n_41), .Y(n_381) );
XNOR2xp5_ASAP7_75t_L g382 ( .A(n_365), .B(n_46), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_356), .B(n_48), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_329), .B(n_49), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_330), .B(n_50), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_364), .B(n_53), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_370), .B(n_199), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_337), .B(n_55), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_328), .B(n_57), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_366), .B(n_126), .C(n_139), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_327), .B(n_58), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_339), .A2(n_346), .B(n_368), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_328), .B(n_59), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_333), .B(n_61), .Y(n_397) );
XOR2x2_ASAP7_75t_L g398 ( .A(n_335), .B(n_63), .Y(n_398) );
XNOR2xp5_ASAP7_75t_L g399 ( .A(n_336), .B(n_64), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_345), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_340), .B(n_65), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_363), .B(n_66), .Y(n_402) );
XNOR2x1_ASAP7_75t_L g403 ( .A(n_357), .B(n_69), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_370), .B(n_190), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_332), .Y(n_406) );
OAI332xp33_ASAP7_75t_L g407 ( .A1(n_341), .A2(n_138), .A3(n_142), .B1(n_133), .B2(n_135), .B3(n_137), .C1(n_70), .C2(n_168), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_342), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_343), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_355), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_368), .B(n_190), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_361), .Y(n_413) );
XNOR2xp5_ASAP7_75t_L g414 ( .A(n_349), .B(n_135), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_354), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_347), .B(n_126), .C(n_137), .Y(n_416) );
XNOR2x1_ASAP7_75t_L g417 ( .A(n_351), .B(n_190), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_352), .B(n_138), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_358), .Y(n_419) );
NAND2xp33_ASAP7_75t_SL g420 ( .A(n_367), .B(n_154), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_338), .B(n_126), .Y(n_421) );
AO22x1_ASAP7_75t_L g422 ( .A1(n_347), .A2(n_154), .B1(n_126), .B2(n_168), .Y(n_422) );
XNOR2xp5_ASAP7_75t_L g423 ( .A(n_359), .B(n_172), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_330), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_344), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_333), .B(n_356), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_348), .Y(n_427) );
XOR2x2_ASAP7_75t_L g428 ( .A(n_335), .B(n_150), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_326), .A2(n_369), .B(n_328), .Y(n_429) );
XOR2xp5_ASAP7_75t_L g430 ( .A(n_329), .B(n_150), .Y(n_430) );
AO21x1_ASAP7_75t_L g431 ( .A1(n_366), .A2(n_346), .B(n_326), .Y(n_431) );
NAND4xp75_ASAP7_75t_L g432 ( .A(n_431), .B(n_395), .C(n_389), .D(n_405), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_395), .A2(n_408), .B1(n_409), .B2(n_429), .Y(n_433) );
INVxp33_ASAP7_75t_L g434 ( .A(n_428), .Y(n_434) );
XOR2x2_ASAP7_75t_SL g435 ( .A(n_398), .B(n_372), .Y(n_435) );
XOR2xp5_ASAP7_75t_L g436 ( .A(n_430), .B(n_399), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_426), .Y(n_437) );
NOR2x1p5_ASAP7_75t_L g438 ( .A(n_376), .B(n_393), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_373), .B(n_378), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_393), .B(n_378), .Y(n_440) );
AOI211xp5_ASAP7_75t_L g441 ( .A1(n_382), .A2(n_379), .B(n_410), .C(n_381), .Y(n_441) );
AOI322xp5_ASAP7_75t_L g442 ( .A1(n_427), .A2(n_424), .A3(n_374), .B1(n_377), .B2(n_375), .C1(n_413), .C2(n_371), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_419), .A2(n_415), .B1(n_374), .B2(n_403), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_400), .Y(n_444) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_426), .A2(n_388), .B(n_425), .Y(n_445) );
INVxp33_ASAP7_75t_SL g446 ( .A(n_423), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_385), .Y(n_447) );
CKINVDCx6p67_ASAP7_75t_R g448 ( .A(n_402), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_386), .Y(n_449) );
INVxp33_ASAP7_75t_L g450 ( .A(n_434), .Y(n_450) );
AOI211xp5_ASAP7_75t_SL g451 ( .A1(n_439), .A2(n_391), .B(n_407), .C(n_380), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_440), .A2(n_402), .B(n_404), .Y(n_452) );
OAI211xp5_ASAP7_75t_SL g453 ( .A1(n_433), .A2(n_384), .B(n_394), .C(n_411), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_433), .A2(n_390), .B1(n_404), .B2(n_396), .Y(n_454) );
O2A1O1Ixp5_ASAP7_75t_L g455 ( .A1(n_435), .A2(n_420), .B(n_422), .C(n_412), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_448), .B(n_404), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_432), .B(n_407), .C(n_401), .Y(n_457) );
AOI21xp33_ASAP7_75t_SL g458 ( .A1(n_443), .A2(n_417), .B(n_392), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_442), .A2(n_416), .B(n_414), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_459), .A2(n_446), .B1(n_444), .B2(n_449), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_450), .A2(n_441), .B(n_444), .C(n_445), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_456), .A2(n_436), .B1(n_438), .B2(n_416), .Y(n_462) );
AO22x2_ASAP7_75t_L g463 ( .A1(n_452), .A2(n_447), .B1(n_437), .B2(n_406), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_457), .B(n_421), .C(n_383), .Y(n_464) );
OR3x2_ASAP7_75t_L g465 ( .A(n_460), .B(n_458), .C(n_455), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_464), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_466), .Y(n_468) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_467), .B(n_462), .Y(n_469) );
OR2x6_ASAP7_75t_L g470 ( .A(n_468), .B(n_463), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_470), .A2(n_465), .B1(n_469), .B2(n_454), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_471), .A2(n_451), .B1(n_453), .B2(n_387), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_472), .A2(n_418), .B(n_397), .Y(n_473) );
endmodule