module real_jpeg_1723_n_16 (n_5, n_4, n_8, n_0, n_12, n_325, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_325;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_1),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_1),
.B(n_29),
.C(n_43),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_1),
.B(n_32),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_1),
.B(n_64),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_1),
.A2(n_64),
.B(n_182),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_1),
.B(n_126),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_1),
.A2(n_58),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_29),
.B1(n_36),
.B2(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_2),
.A2(n_48),
.B1(n_58),
.B2(n_60),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_4),
.A2(n_58),
.B1(n_60),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_29),
.B1(n_36),
.B2(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_109),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_5),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_5),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_5),
.A2(n_35),
.B1(n_58),
.B2(n_60),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_58),
.B1(n_60),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_67),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_205)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_11),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_11),
.A2(n_39),
.B1(n_58),
.B2(n_60),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_12),
.A2(n_58),
.B1(n_60),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_69),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_13),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_13),
.A2(n_29),
.B1(n_36),
.B2(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_13),
.A2(n_58),
.B1(n_60),
.B2(n_72),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_315),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_305),
.B(n_314),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_271),
.B(n_302),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_248),
.B(n_270),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_135),
.B(n_247),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_110),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_22),
.B(n_110),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_93),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_23),
.B(n_82),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_55),
.C(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_26),
.B(n_40),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_37),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_27),
.A2(n_31),
.B(n_86),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_31),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_27),
.A2(n_37),
.B(n_86),
.Y(n_184)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_28),
.B(n_38),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_28),
.A2(n_85),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_32),
.B1(n_98),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_28),
.A2(n_32),
.B1(n_162),
.B2(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_29),
.B(n_160),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_31),
.A2(n_88),
.B(n_102),
.Y(n_210)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_44),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_41),
.A2(n_91),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_41),
.B(n_199),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_52)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_46),
.B1(n_75),
.B2(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_45),
.B(n_77),
.Y(n_183)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_46),
.B(n_152),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_46),
.A2(n_64),
.A3(n_75),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_49),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_50),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_51),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_51),
.A2(n_119),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_51),
.A2(n_119),
.B1(n_147),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_51),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_51),
.A2(n_119),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_70),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_56),
.A2(n_68),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_56),
.A2(n_62),
.B1(n_108),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_56),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_56),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_56),
.A2(n_62),
.B1(n_276),
.B2(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_56),
.A2(n_259),
.B(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_63),
.B(n_97),
.C(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_98),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_61),
.C(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_62),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_64),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B(n_79),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_71),
.A2(n_73),
.B(n_78),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_73),
.A2(n_78),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_73),
.A2(n_78),
.B1(n_104),
.B2(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_79),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_81),
.A2(n_131),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_81),
.A2(n_131),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_92),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_91),
.A2(n_118),
.B(n_199),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_93),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_107),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_94),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_227),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_100),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_103),
.B(n_107),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_105),
.B(n_130),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_134),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_114),
.B(n_121),
.C(n_134),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_115),
.A2(n_116),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_116),
.B(n_117),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_116),
.A2(n_256),
.B(n_261),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_124),
.B(n_128),
.C(n_133),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_125),
.B(n_277),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_126),
.B(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_127),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_129),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_131),
.A2(n_267),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

AOI321xp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_229),
.A3(n_239),
.B1(n_245),
.B2(n_246),
.C(n_325),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_213),
.B(n_228),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_193),
.B(n_212),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_175),
.B(n_192),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_156),
.B(n_174),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_146),
.C(n_177),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_168),
.B(n_173),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_166),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_178),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_186),
.C(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_211),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_211),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_200),
.C(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_208),
.C(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_215),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_223),
.B2(n_224),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_225),
.C(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_217),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_221),
.CI(n_222),
.CON(n_217),
.SN(n_217)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_238),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_234),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_269),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_269),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_254),
.C(n_262),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_262),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_265),
.B(n_268),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_294),
.C(n_298),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_268),
.B(n_294),
.CI(n_298),
.CON(n_301),
.SN(n_301)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_299),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_293),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_275),
.C(n_292),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.C(n_281),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_284),
.B1(n_291),
.B2(n_292),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_291),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_281),
.B1(n_290),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_285),
.C(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_307),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_311),
.C(n_313),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);


endmodule