module fake_jpeg_13022_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_54),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_13),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_84),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_13),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_0),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_102),
.Y(n_175)
);

BUFx12f_ASAP7_75t_SL g102 ( 
.A(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_54),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_108),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_28),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_28),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_117),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_128),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_18),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_46),
.A2(n_20),
.B1(n_43),
.B2(n_39),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_41),
.B1(n_31),
.B2(n_20),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_61),
.B(n_23),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_52),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_91),
.B(n_41),
.Y(n_148)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_164),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_107),
.A2(n_93),
.B1(n_89),
.B2(n_83),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_125),
.B1(n_101),
.B2(n_140),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_62),
.B1(n_76),
.B2(n_74),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_166),
.B1(n_185),
.B2(n_191),
.Y(n_210)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_67),
.B1(n_73),
.B2(n_71),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_165),
.A2(n_187),
.B(n_104),
.C(n_151),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_69),
.B1(n_66),
.B2(n_65),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

BUFx4f_ASAP7_75t_SL g170 ( 
.A(n_113),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_174),
.Y(n_212)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_190),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_105),
.B(n_108),
.C(n_98),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_184),
.B(n_142),
.CI(n_133),
.CON(n_209),
.SN(n_209)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_105),
.A2(n_64),
.B1(n_55),
.B2(n_81),
.Y(n_185)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_126),
.A2(n_53),
.B1(n_20),
.B2(n_23),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_95),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_114),
.B(n_45),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_131),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_95),
.A2(n_26),
.B1(n_37),
.B2(n_28),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_201),
.B1(n_134),
.B2(n_115),
.Y(n_231)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_195),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_117),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_120),
.A2(n_37),
.B1(n_45),
.B2(n_47),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_203),
.B(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_205),
.A2(n_182),
.B1(n_178),
.B2(n_180),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_162),
.C(n_155),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_223),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_176),
.A2(n_97),
.B1(n_123),
.B2(n_153),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_140),
.B1(n_125),
.B2(n_118),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_231),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_153),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_158),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_188),
.B(n_184),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_238),
.B(n_243),
.Y(n_298)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_192),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_192),
.A3(n_187),
.B1(n_161),
.B2(n_190),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_269),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_187),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_160),
.B(n_157),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_251),
.B(n_253),
.Y(n_273)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_157),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_244),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_165),
.B(n_187),
.C(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_259),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_165),
.B(n_170),
.C(n_198),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_258),
.B1(n_220),
.B2(n_228),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_227),
.A2(n_165),
.B1(n_196),
.B2(n_163),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_264),
.B1(n_235),
.B2(n_206),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_167),
.B1(n_173),
.B2(n_159),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_207),
.A2(n_172),
.B1(n_171),
.B2(n_174),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_123),
.B1(n_97),
.B2(n_151),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_207),
.A2(n_216),
.B1(n_232),
.B2(n_202),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_226),
.B(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_220),
.B1(n_228),
.B2(n_203),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_210),
.A2(n_177),
.B1(n_195),
.B2(n_168),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_268),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_212),
.B(n_204),
.Y(n_284)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_154),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_237),
.B1(n_231),
.B2(n_215),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_279),
.B1(n_281),
.B2(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_271),
.B(n_278),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_287),
.B(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_249),
.B(n_224),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_204),
.B1(n_202),
.B2(n_220),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_283),
.B(n_253),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_293),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_228),
.B1(n_208),
.B2(n_233),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_217),
.B(n_233),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_230),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_295),
.C(n_251),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_247),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_278),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_217),
.B(n_235),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_221),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_211),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_301),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_246),
.A2(n_208),
.B1(n_234),
.B2(n_211),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_254),
.B1(n_259),
.B2(n_269),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_221),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_270),
.A2(n_266),
.B1(n_262),
.B2(n_261),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_305),
.A2(n_310),
.B(n_326),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_307),
.A2(n_289),
.B1(n_281),
.B2(n_288),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_270),
.A2(n_240),
.B1(n_242),
.B2(n_241),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_309),
.A2(n_316),
.B1(n_320),
.B2(n_273),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_313),
.B(n_333),
.Y(n_344)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_265),
.Y(n_315)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_263),
.B1(n_253),
.B2(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_248),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_323),
.C(n_330),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_319),
.B(n_318),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_253),
.B1(n_251),
.B2(n_245),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_332),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_239),
.Y(n_322)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_206),
.C(n_251),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_277),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_327),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_253),
.B1(n_208),
.B2(n_112),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_211),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_234),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_329),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_234),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_170),
.C(n_136),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_333),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_301),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_271),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_285),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_218),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_335),
.B(n_274),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_336),
.A2(n_352),
.B1(n_306),
.B2(n_307),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_312),
.A2(n_273),
.B(n_320),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_337),
.A2(n_312),
.B(n_326),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_347),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_353),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_290),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_349),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_351),
.A2(n_355),
.B1(n_358),
.B2(n_361),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_289),
.B1(n_273),
.B2(n_288),
.Y(n_352)
);

INVx6_ASAP7_75t_SL g353 ( 
.A(n_325),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_303),
.A2(n_282),
.B1(n_283),
.B2(n_297),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_290),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_362),
.C(n_366),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_298),
.B(n_287),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_357),
.A2(n_314),
.B(n_308),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_303),
.A2(n_282),
.B1(n_283),
.B2(n_276),
.Y(n_358)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_305),
.A2(n_282),
.B1(n_292),
.B2(n_299),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_295),
.C(n_298),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_324),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_280),
.Y(n_364)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_364),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_280),
.C(n_136),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_286),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_367),
.B(n_328),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_340),
.B(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_374),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_302),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_375),
.B(n_387),
.Y(n_409)
);

AO21x1_ASAP7_75t_L g417 ( 
.A1(n_377),
.A2(n_218),
.B(n_1),
.Y(n_417)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_361),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_316),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_309),
.B1(n_306),
.B2(n_302),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_352),
.A2(n_363),
.B1(n_337),
.B2(n_365),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_385),
.A2(n_392),
.B1(n_393),
.B2(n_355),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_365),
.B(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_329),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_341),
.B(n_327),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_390),
.B(n_395),
.Y(n_420)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_394),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_339),
.A2(n_331),
.B1(n_317),
.B2(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_353),
.B(n_367),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_286),
.B1(n_141),
.B2(n_124),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_396),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_354),
.C(n_343),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_399),
.B(n_402),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g401 ( 
.A1(n_377),
.A2(n_342),
.B(n_357),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_354),
.C(n_386),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_366),
.C(n_356),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_382),
.C(n_373),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_380),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_339),
.B1(n_360),
.B2(n_351),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_411),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_408),
.A2(n_415),
.B1(n_422),
.B2(n_378),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_394),
.B(n_387),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_397),
.A2(n_340),
.B1(n_358),
.B2(n_362),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_371),
.A2(n_346),
.B1(n_347),
.B2(n_218),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_421),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_392),
.A2(n_346),
.B1(n_218),
.B2(n_2),
.Y(n_415)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_0),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_418),
.B(n_388),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_369),
.A2(n_28),
.B1(n_32),
.B2(n_2),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_372),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_426),
.B(n_437),
.Y(n_451)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_420),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_442),
.Y(n_455)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_430),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_441),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_369),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_433),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_374),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_423),
.Y(n_435)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_438),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_382),
.C(n_393),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_445),
.C(n_446),
.Y(n_454)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_424),
.Y(n_440)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_424),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_406),
.A2(n_408),
.B1(n_400),
.B2(n_414),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_444),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_391),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_410),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_412),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_448),
.A2(n_417),
.B1(n_389),
.B2(n_384),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_427),
.A2(n_414),
.B1(n_403),
.B2(n_416),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_450),
.A2(n_453),
.B1(n_460),
.B2(n_429),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_427),
.A2(n_403),
.B1(n_398),
.B2(n_419),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_407),
.C(n_398),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_458),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_418),
.C(n_419),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_425),
.A2(n_412),
.B(n_381),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_459),
.A2(n_464),
.B(n_368),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_439),
.A2(n_370),
.B1(n_368),
.B2(n_421),
.Y(n_463)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_370),
.C(n_415),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_456),
.A2(n_426),
.B1(n_436),
.B2(n_446),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_470),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_452),
.A2(n_436),
.B1(n_445),
.B2(n_444),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_472),
.A2(n_483),
.B(n_466),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_432),
.C(n_431),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_475),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_467),
.A2(n_441),
.B1(n_422),
.B2(n_4),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_481),
.B1(n_482),
.B2(n_483),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_11),
.C(n_3),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_478),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_11),
.C(n_3),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_480),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_455),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_4),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_467),
.A2(n_6),
.B(n_7),
.Y(n_483)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_485),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_473),
.B(n_464),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_488),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_461),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_468),
.B(n_461),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_489),
.A2(n_490),
.B(n_491),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_453),
.C(n_458),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_470),
.A2(n_463),
.B(n_465),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_494),
.Y(n_503)
);

BUFx4f_ASAP7_75t_SL g494 ( 
.A(n_475),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_477),
.A2(n_449),
.B(n_450),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_496),
.A2(n_8),
.B(n_9),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_478),
.C(n_481),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_502),
.Y(n_511)
);

AO21x1_ASAP7_75t_L g500 ( 
.A1(n_495),
.A2(n_476),
.B(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_500),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g501 ( 
.A1(n_492),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_501),
.A2(n_486),
.B(n_494),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_6),
.C(n_8),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_6),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_504),
.B(n_8),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_497),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_499),
.Y(n_508)
);

O2A1O1Ixp33_ASAP7_75t_SL g518 ( 
.A1(n_508),
.A2(n_500),
.B(n_501),
.C(n_11),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_503),
.C(n_507),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_513),
.B(n_514),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_484),
.C(n_494),
.Y(n_513)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_515),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_503),
.C(n_511),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_516),
.A2(n_518),
.B(n_9),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_520),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_517),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_519),
.C(n_10),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_523),
.B(n_9),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_9),
.B(n_11),
.Y(n_525)
);


endmodule