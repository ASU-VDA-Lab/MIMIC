module fake_jpeg_30316_n_515 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_64),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_55),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_49),
.Y(n_124)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_72),
.Y(n_134)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_97),
.Y(n_152)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_37),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_19),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_125),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_41),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_19),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_147),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_73),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_26),
.C(n_47),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_21),
.C(n_25),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_20),
.Y(n_147)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_55),
.B(n_29),
.Y(n_149)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_130),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_86),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_20),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_21),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_161),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_109),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_163),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_181),
.Y(n_227)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_166),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_29),
.B1(n_36),
.B2(n_43),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_178),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_104),
.A2(n_92),
.B1(n_131),
.B2(n_36),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_117),
.A2(n_71),
.B1(n_98),
.B2(n_96),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_182),
.B1(n_187),
.B2(n_192),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_176),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_104),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_77),
.B1(n_95),
.B2(n_91),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_185),
.B(n_208),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_131),
.A2(n_32),
.B1(n_31),
.B2(n_47),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_211),
.B1(n_215),
.B2(n_153),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_75),
.B1(n_82),
.B2(n_81),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_116),
.A2(n_80),
.B1(n_79),
.B2(n_101),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_191),
.A2(n_138),
.B1(n_116),
.B2(n_56),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_134),
.A2(n_68),
.B1(n_63),
.B2(n_57),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_198),
.Y(n_251)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_106),
.B(n_39),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_195),
.B(n_212),
.Y(n_244)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_210),
.B1(n_189),
.B2(n_207),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_106),
.B(n_39),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_134),
.B(n_39),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_213),
.B(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_126),
.B(n_39),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_39),
.Y(n_215)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_185),
.A2(n_149),
.B1(n_118),
.B2(n_122),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_175),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_226),
.A2(n_245),
.B1(n_250),
.B2(n_252),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_231),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_167),
.A2(n_149),
.B(n_86),
.C(n_141),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_232),
.A2(n_199),
.B(n_161),
.C(n_206),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_138),
.B1(n_112),
.B2(n_142),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_248),
.B1(n_206),
.B2(n_163),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_156),
.B1(n_144),
.B2(n_137),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_192),
.A2(n_137),
.B1(n_156),
.B2(n_153),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_178),
.A2(n_150),
.B1(n_42),
.B2(n_129),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_164),
.A2(n_42),
.B1(n_25),
.B2(n_41),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_162),
.A2(n_42),
.B1(n_59),
.B2(n_43),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_163),
.B1(n_172),
.B2(n_210),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_162),
.B(n_37),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_219),
.C(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_179),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_262),
.B(n_269),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_264),
.A2(n_279),
.B1(n_283),
.B2(n_287),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_227),
.B(n_169),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_265),
.B(n_302),
.Y(n_308)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_266),
.Y(n_328)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_190),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_277),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_244),
.B(n_233),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_166),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_273),
.B(n_282),
.Y(n_318)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_281),
.Y(n_310)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_222),
.A2(n_184),
.B1(n_194),
.B2(n_165),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

CKINVDCx12_ASAP7_75t_R g281 ( 
.A(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_196),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_173),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_285),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_180),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_232),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_297),
.C(n_225),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_222),
.A2(n_200),
.B1(n_201),
.B2(n_172),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_220),
.B(n_202),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_220),
.B(n_197),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_250),
.B(n_245),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_293),
.B(n_294),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_203),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_228),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_170),
.C(n_176),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_235),
.B(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_298),
.B(n_299),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_209),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_261),
.B(n_13),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_271),
.A2(n_241),
.B1(n_236),
.B2(n_248),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_303),
.A2(n_313),
.B1(n_316),
.B2(n_322),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_241),
.B(n_240),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_305),
.A2(n_309),
.B(n_324),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_292),
.A2(n_240),
.B(n_239),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_296),
.A2(n_226),
.B1(n_239),
.B2(n_256),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_276),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_319),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_256),
.B1(n_174),
.B2(n_205),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_260),
.Y(n_319)
);

AO21x2_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_239),
.B(n_221),
.Y(n_321)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_277),
.A2(n_204),
.B1(n_217),
.B2(n_228),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_238),
.B1(n_257),
.B2(n_255),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_323),
.A2(n_339),
.B1(n_280),
.B2(n_301),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_284),
.A2(n_238),
.B(n_237),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_286),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_288),
.A2(n_225),
.B(n_103),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_330),
.A2(n_335),
.B(n_270),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_263),
.A2(n_295),
.B1(n_267),
.B2(n_289),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_272),
.B(n_237),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_268),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_263),
.A2(n_208),
.B1(n_234),
.B2(n_218),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_328),
.Y(n_341)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_365),
.C(n_326),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_343),
.B(n_346),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_333),
.B(n_285),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_344),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_333),
.B(n_266),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_308),
.B(n_279),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_349),
.B(n_352),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_274),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_355),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_311),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_351),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_334),
.B(n_297),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_275),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_356),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_332),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_364),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_278),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_359),
.B(n_361),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_290),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g388 ( 
.A1(n_360),
.A2(n_371),
.B(n_337),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_307),
.B(n_300),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_313),
.B1(n_316),
.B2(n_303),
.Y(n_378)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_291),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_368),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_367),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_370),
.Y(n_387)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_317),
.B(n_264),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_372),
.B(n_353),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_388),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_378),
.A2(n_384),
.B1(n_390),
.B2(n_344),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_365),
.C(n_360),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_343),
.C(n_358),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_322),
.B1(n_304),
.B2(n_321),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_373),
.A2(n_306),
.B1(n_317),
.B2(n_305),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_385),
.A2(n_394),
.B1(n_397),
.B2(n_363),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_321),
.B(n_336),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_403),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_368),
.A2(n_304),
.B1(n_321),
.B2(n_306),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_321),
.B1(n_323),
.B2(n_304),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_312),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_395),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_312),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_396),
.B(n_338),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_324),
.B1(n_338),
.B2(n_314),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_401),
.A2(n_383),
.B1(n_400),
.B2(n_390),
.Y(n_413)
);

NOR2x1_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_381),
.Y(n_405)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_405),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_406),
.A2(n_410),
.B1(n_421),
.B2(n_426),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_407),
.A2(n_408),
.B1(n_414),
.B2(n_419),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_345),
.B1(n_360),
.B2(n_353),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_384),
.A2(n_359),
.B1(n_361),
.B2(n_345),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_417),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_397),
.A2(n_357),
.B1(n_372),
.B2(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_418),
.Y(n_431)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_385),
.A2(n_357),
.B1(n_341),
.B2(n_356),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_382),
.A2(n_378),
.B1(n_391),
.B2(n_399),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_422),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_357),
.B1(n_347),
.B2(n_364),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_369),
.C(n_366),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_376),
.C(n_402),
.Y(n_442)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_425),
.Y(n_436)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_380),
.A2(n_362),
.B1(n_354),
.B2(n_320),
.Y(n_426)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_428),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_382),
.B(n_327),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_407),
.A2(n_392),
.B1(n_389),
.B2(n_398),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_437),
.B1(n_410),
.B2(n_429),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_374),
.B1(n_392),
.B2(n_401),
.Y(n_434)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_414),
.A2(n_389),
.B1(n_398),
.B2(n_403),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_406),
.A2(n_401),
.B1(n_403),
.B2(n_389),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_438),
.A2(n_430),
.B1(n_435),
.B2(n_429),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_379),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_415),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_446),
.C(n_415),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_393),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_445),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_421),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_402),
.C(n_315),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_409),
.A2(n_375),
.B(n_327),
.Y(n_447)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_448),
.A2(n_419),
.B1(n_408),
.B2(n_409),
.Y(n_449)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_450),
.B(n_451),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_452),
.A2(n_447),
.B1(n_431),
.B2(n_439),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_426),
.C(n_424),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_454),
.C(n_431),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_418),
.C(n_416),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_405),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_457),
.A2(n_463),
.B(n_443),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_427),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_459),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_404),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_432),
.B(n_375),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_430),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_442),
.B(n_234),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_465),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_438),
.A2(n_229),
.B(n_223),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_229),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_469),
.B(n_37),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_435),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_472),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_474),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_433),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_456),
.B(n_440),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_476),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_42),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_453),
.C(n_450),
.Y(n_481)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_480),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_490)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_483),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_473),
.A2(n_451),
.B(n_455),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_452),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_486),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_37),
.C(n_48),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_15),
.C(n_14),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_490),
.A2(n_471),
.B1(n_477),
.B2(n_2),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_480),
.A2(n_11),
.B(n_1),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_478),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_493),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_491),
.A2(n_474),
.B1(n_476),
.B2(n_479),
.Y(n_494)
);

AOI322xp5_ASAP7_75t_L g504 ( 
.A1(n_494),
.A2(n_493),
.A3(n_499),
.B1(n_500),
.B2(n_50),
.C1(n_6),
.C2(n_7),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_467),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_497),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_0),
.C(n_1),
.Y(n_503)
);

AOI321xp33_ASAP7_75t_L g501 ( 
.A1(n_496),
.A2(n_482),
.A3(n_481),
.B1(n_488),
.B2(n_486),
.C(n_492),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_503),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_504),
.B(n_4),
.C(n_5),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_505),
.A2(n_2),
.B(n_3),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_506),
.B(n_507),
.Y(n_509)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_508),
.A2(n_502),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_4),
.C2(n_10),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_4),
.C(n_8),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_509),
.B(n_9),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_512),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_48),
.B(n_502),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_514),
.A2(n_48),
.B(n_239),
.Y(n_515)
);


endmodule