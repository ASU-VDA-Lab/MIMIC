module fake_jpeg_17768_n_183 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_1),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_19),
.B(n_30),
.Y(n_44)
);

OR2x4_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_40),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_15),
.B1(n_16),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_51),
.B1(n_56),
.B2(n_17),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_57),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_24),
.B1(n_16),
.B2(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_30),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_29),
.B(n_26),
.C(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_68),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_31),
.B1(n_17),
.B2(n_21),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_72),
.B1(n_73),
.B2(n_1),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_75),
.Y(n_80)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_59),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_21),
.B1(n_25),
.B2(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_95),
.B1(n_72),
.B2(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_28),
.B(n_27),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_70),
.A3(n_62),
.B1(n_60),
.B2(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_46),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_109),
.B1(n_94),
.B2(n_85),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_5),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_106),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_28),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_113),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_95),
.B1(n_87),
.B2(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_48),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_81),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_127),
.B1(n_101),
.B2(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_125),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_93),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_27),
.B(n_26),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_79),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_105),
.B1(n_110),
.B2(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_112),
.C(n_97),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_97),
.B(n_108),
.C(n_104),
.D(n_107),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_135),
.A2(n_142),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_125),
.C(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_115),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_127),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_129),
.C(n_28),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_122),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_146),
.C(n_152),
.Y(n_160)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_6),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_7),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_7),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_135),
.B1(n_142),
.B2(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_148),
.B(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_158),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_8),
.C(n_9),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_146),
.C(n_152),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_149),
.B(n_151),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_12),
.B1(n_14),
.B2(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_160),
.B(n_9),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_174),
.B(n_12),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_8),
.C(n_10),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_177),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_178),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_166),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_170),
.Y(n_183)
);


endmodule