module real_jpeg_490_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_13),
.C(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_16),
.B1(n_33),
.B2(n_39),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_41),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_27),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_22),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_20),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_17),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_18),
.Y(n_19)
);

AO22x1_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_13),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_13),
.B(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

OA21x2_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_37),
.B(n_40),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_38),
.Y(n_37)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_26),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);


endmodule