module real_jpeg_32451_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_0),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_0),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_0),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_2),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_2),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_2),
.B(n_161),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_2),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_2),
.B(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_2),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_2),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_3),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_3),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_472),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_4),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_5),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_9),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_9),
.B(n_136),
.Y(n_135)
);

NAND2x1_ASAP7_75t_L g160 ( 
.A(n_9),
.B(n_161),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_10),
.B(n_49),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_10),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_10),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_10),
.B(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_10),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_10),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_11),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_11),
.B(n_103),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_11),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_11),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_11),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_11),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_11),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_12),
.B(n_86),
.Y(n_237)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_12),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_12),
.B(n_379),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_12),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_13),
.Y(n_310)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_16),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_17),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_17),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_17),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_17),
.B(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_202),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_200),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_22),
.B(n_166),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_94),
.C(n_127),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_24),
.B(n_95),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_65),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_25),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_39),
.B(n_64),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_26),
.B(n_40),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_35),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_29),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_34),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_34),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_34),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_35),
.B(n_99),
.C(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_35),
.A2(n_36),
.B1(n_236),
.B2(n_237),
.Y(n_339)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_36),
.B(n_193),
.C(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_38),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_38),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_53),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_53),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_52),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_42),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_42),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_42),
.A2(n_145),
.B1(n_275),
.B2(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_44),
.Y(n_367)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_44),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_54),
.B1(n_55),
.B2(n_63),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_91),
.C(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_63),
.Y(n_144)
);

AO22x1_ASAP7_75t_SL g448 ( 
.A1(n_45),
.A2(n_63),
.B1(n_365),
.B2(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_46),
.Y(n_438)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_51),
.Y(n_153)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_52),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_53),
.Y(n_254)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_60),
.B(n_154),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_62),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_63),
.B(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_83),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_66),
.B(n_168),
.C(n_169),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_78),
.C(n_79),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_67),
.B(n_164),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.C(n_74),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_74),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_68),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_68),
.A2(n_132),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_70),
.B(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_72),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_77),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_88),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_80),
.B(n_85),
.C(n_89),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_91),
.B(n_118),
.C(n_121),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_115),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_114),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_97),
.B(n_114),
.C(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_105),
.C(n_108),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_104)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_135),
.C(n_139),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_105),
.A2(n_113),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_112),
.Y(n_286)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_118),
.A2(n_191),
.B1(n_192),
.B2(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_118),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_118),
.B(n_279),
.C(n_282),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_118),
.A2(n_195),
.B1(n_282),
.B2(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_119),
.Y(n_385)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_120),
.Y(n_242)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_120),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_123),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_127),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_146),
.C(n_162),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_129),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_142),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_130),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_134),
.A2(n_142),
.B1(n_143),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_134),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_135),
.B(n_139),
.Y(n_290)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_146),
.A2(n_147),
.B1(n_162),
.B2(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.C(n_160),
.Y(n_147)
);

XOR2x2_ASAP7_75t_L g250 ( 
.A(n_148),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_154),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_150),
.Y(n_231)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_154),
.B(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g277 ( 
.A(n_155),
.Y(n_277)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_155),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_157),
.B(n_160),
.Y(n_251)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_184),
.Y(n_171)
);

XOR2x1_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_183),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_192),
.B(n_339),
.Y(n_338)
);

BUFx4f_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_466),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_295),
.C(n_460),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_258),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g466 ( 
.A1(n_206),
.A2(n_259),
.B(n_467),
.C(n_470),
.D(n_471),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_256),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_207),
.B(n_256),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_252),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_209),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g294 ( 
.A(n_212),
.B(n_253),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_232),
.C(n_248),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_267),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_222),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g343 ( 
.A(n_214),
.B(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_216),
.A2(n_217),
.B1(n_222),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_217),
.A2(n_218),
.B(n_219),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_222),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_229),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_223),
.A2(n_224),
.B1(n_229),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_234),
.B1(n_249),
.B2(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.C(n_243),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_242),
.Y(n_414)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_293),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_260),
.B(n_293),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.C(n_268),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_262),
.B(n_266),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_268),
.B(n_465),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_287),
.C(n_291),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_269),
.B(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_278),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_274),
.B1(n_278),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_286),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_288),
.B(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2x1p5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_351),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_341),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_297),
.B(n_341),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.C(n_324),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_325),
.Y(n_354)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_321),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_303),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_321),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_311),
.C(n_318),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_307),
.B(n_389),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_310),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_311),
.A2(n_312),
.B1(n_318),
.B2(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_313),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_337),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_347),
.C(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.C(n_333),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_334),
.Y(n_370)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_349),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_343),
.B(n_349),
.C(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_346),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_371),
.B(n_459),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_353),
.B(n_355),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.C(n_368),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_369),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.C(n_364),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_360),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_361),
.B(n_406),
.Y(n_417)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

BUFx4f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_392),
.B(n_458),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_390),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_373),
.B(n_390),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.C(n_386),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_455),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_377),
.A2(n_387),
.B1(n_388),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_377),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_381),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_383),
.B(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_452),
.B(n_457),
.Y(n_392)
);

OAI21x1_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_440),
.B(n_451),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_421),
.B(n_439),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_407),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_407),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_403),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_398),
.A2(n_399),
.B1(n_403),
.B2(n_404),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_398),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_415),
.B2(n_416),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_413),
.C(n_415),
.Y(n_450)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_418),
.Y(n_446)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_433),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_432),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_432),
.B(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_437),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx8_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_450),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_450),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_445),
.C(n_448),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_454),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_468),
.B(n_469),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_462),
.B(n_464),
.Y(n_468)
);


endmodule