module fake_jpeg_20348_n_206 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_10),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_17),
.B1(n_21),
.B2(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_17),
.B1(n_15),
.B2(n_13),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_13),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_22),
.B1(n_20),
.B2(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_23),
.B1(n_28),
.B2(n_31),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_36),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_23),
.B1(n_28),
.B2(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_67),
.B(n_46),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_38),
.A3(n_39),
.B1(n_40),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_19),
.B1(n_32),
.B2(n_39),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_68),
.B1(n_40),
.B2(n_49),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_29),
.C(n_27),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_46),
.C(n_42),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_86),
.B(n_69),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_43),
.B1(n_54),
.B2(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_46),
.B1(n_55),
.B2(n_52),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_59),
.B(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_46),
.B1(n_40),
.B2(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_29),
.B(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_88),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_49),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_78),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_95),
.B(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_68),
.C(n_57),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_24),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_68),
.B1(n_64),
.B2(n_70),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_84),
.B1(n_70),
.B2(n_71),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_88),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_86),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_112),
.Y(n_131)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_116),
.Y(n_142)
);

XNOR2x2_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_84),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_102),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_99),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_84),
.B(n_82),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_100),
.B1(n_96),
.B2(n_90),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_94),
.C(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_143),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_96),
.B1(n_108),
.B2(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_135),
.B1(n_140),
.B2(n_144),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_101),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_145),
.B(n_144),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_94),
.B1(n_71),
.B2(n_73),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_65),
.C(n_29),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_123),
.C(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_24),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_151),
.Y(n_160)
);

OA21x2_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_109),
.B(n_114),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_155),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_118),
.B(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_107),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_27),
.C(n_26),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_159),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_27),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_27),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_141),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_162),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_140),
.B1(n_129),
.B2(n_138),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_139),
.B1(n_133),
.B2(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_148),
.B1(n_147),
.B2(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_158),
.B1(n_143),
.B2(n_44),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_164),
.B1(n_169),
.B2(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_159),
.C(n_146),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_146),
.B(n_157),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_9),
.B(n_8),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_131),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_41),
.C(n_26),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_170),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_177),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_167),
.B1(n_44),
.B2(n_41),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_26),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_24),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_12),
.B1(n_18),
.B2(n_3),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_174),
.B(n_171),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_193),
.A3(n_7),
.B1(n_18),
.B2(n_12),
.C1(n_4),
.C2(n_0),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_194),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_178),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_185),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_18),
.B1(n_12),
.B2(n_3),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_0),
.C(n_1),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_198),
.C(n_188),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_6),
.B(n_4),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_4),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_199),
.B(n_5),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_204),
.B1(n_201),
.B2(n_5),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_4),
.C(n_6),
.Y(n_206)
);


endmodule