module real_aes_21_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g92 ( .A1(n_0), .A2(n_52), .B1(n_89), .B2(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g189 ( .A(n_1), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_2), .A2(n_48), .B1(n_141), .B2(n_144), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_3), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g246 ( .A(n_4), .Y(n_246) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_5), .A2(n_15), .B1(n_89), .B2(n_90), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_6), .Y(n_261) );
INVx2_ASAP7_75t_L g209 ( .A(n_7), .Y(n_209) );
INVx1_ASAP7_75t_L g280 ( .A(n_8), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_9), .A2(n_77), .B1(n_134), .B2(n_138), .Y(n_133) );
INVx1_ASAP7_75t_L g277 ( .A(n_10), .Y(n_277) );
INVx1_ASAP7_75t_SL g331 ( .A(n_11), .Y(n_331) );
OAI22xp5_ASAP7_75t_SL g164 ( .A1(n_12), .A2(n_30), .B1(n_165), .B2(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g166 ( .A(n_12), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_12), .B(n_229), .Y(n_293) );
AOI33xp33_ASAP7_75t_L g317 ( .A1(n_13), .A2(n_33), .A3(n_214), .B1(n_222), .B2(n_318), .B3(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g254 ( .A(n_14), .Y(n_254) );
OAI221xp5_ASAP7_75t_L g181 ( .A1(n_15), .A2(n_52), .B1(n_57), .B2(n_182), .C(n_184), .Y(n_181) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_16), .A2(n_68), .B(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g239 ( .A(n_16), .B(n_68), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_17), .A2(n_81), .B1(n_82), .B2(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_17), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_18), .B(n_212), .Y(n_328) );
INVx1_ASAP7_75t_L g583 ( .A(n_18), .Y(n_583) );
INVx3_ASAP7_75t_L g89 ( .A(n_19), .Y(n_89) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_20), .A2(n_55), .B1(n_85), .B2(n_102), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_21), .B(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g100 ( .A(n_22), .Y(n_100) );
INVx1_ASAP7_75t_L g191 ( .A(n_23), .Y(n_191) );
AND2x2_ASAP7_75t_L g217 ( .A(n_23), .B(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g235 ( .A(n_23), .B(n_189), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_24), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_25), .B(n_212), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_26), .A2(n_207), .B1(n_271), .B2(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_27), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_28), .B(n_229), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_28), .A2(n_81), .B1(n_82), .B2(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_28), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_29), .B(n_243), .Y(n_248) );
INVx1_ASAP7_75t_L g165 ( .A(n_30), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_30), .B(n_229), .Y(n_247) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_31), .A2(n_57), .B1(n_89), .B2(n_96), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_32), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_34), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g215 ( .A(n_35), .Y(n_215) );
INVx1_ASAP7_75t_L g231 ( .A(n_35), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_36), .A2(n_73), .B1(n_108), .B2(n_114), .Y(n_107) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_37), .A2(n_47), .B1(n_148), .B2(n_151), .Y(n_147) );
AND2x2_ASAP7_75t_L g236 ( .A(n_38), .B(n_237), .Y(n_236) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_39), .A2(n_58), .B1(n_212), .B2(n_220), .C(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_40), .B(n_212), .Y(n_305) );
INVx1_ASAP7_75t_L g101 ( .A(n_41), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_42), .B(n_207), .Y(n_263) );
AOI21xp5_ASAP7_75t_SL g301 ( .A1(n_43), .A2(n_220), .B(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_44), .A2(n_170), .B1(n_171), .B2(n_175), .Y(n_169) );
INVx1_ASAP7_75t_L g175 ( .A(n_44), .Y(n_175) );
INVx1_ASAP7_75t_L g274 ( .A(n_45), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_46), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_46), .Y(n_174) );
INVx1_ASAP7_75t_L g226 ( .A(n_49), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_50), .A2(n_67), .B1(n_155), .B2(n_157), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_51), .A2(n_220), .B(n_225), .Y(n_219) );
INVxp33_ASAP7_75t_L g186 ( .A(n_52), .Y(n_186) );
INVx1_ASAP7_75t_L g218 ( .A(n_53), .Y(n_218) );
INVx1_ASAP7_75t_L g233 ( .A(n_53), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_54), .A2(n_62), .B1(n_126), .B2(n_128), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_56), .B(n_212), .Y(n_320) );
INVxp67_ASAP7_75t_L g185 ( .A(n_57), .Y(n_185) );
AND2x2_ASAP7_75t_L g333 ( .A(n_59), .B(n_206), .Y(n_333) );
INVx1_ASAP7_75t_L g275 ( .A(n_60), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_61), .A2(n_220), .B(n_330), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_63), .A2(n_220), .B(n_292), .C(n_296), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_64), .A2(n_168), .B1(n_169), .B2(n_176), .Y(n_167) );
INVx1_ASAP7_75t_L g176 ( .A(n_64), .Y(n_176) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_65), .B(n_206), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_66), .A2(n_220), .B1(n_315), .B2(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g303 ( .A(n_69), .Y(n_303) );
INVx1_ASAP7_75t_L g172 ( .A(n_70), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_71), .A2(n_81), .B1(n_82), .B2(n_161), .Y(n_80) );
INVx1_ASAP7_75t_L g161 ( .A(n_71), .Y(n_161) );
AND2x2_ASAP7_75t_L g321 ( .A(n_72), .B(n_206), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_74), .A2(n_252), .B(n_253), .C(n_256), .Y(n_251) );
BUFx2_ASAP7_75t_SL g183 ( .A(n_75), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_76), .B(n_229), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_178), .B1(n_192), .B2(n_563), .C(n_565), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_162), .Y(n_79) );
INVx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OR2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_132), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_107), .C(n_119), .D(n_125), .Y(n_83) );
BUFx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x4_ASAP7_75t_L g86 ( .A(n_87), .B(n_94), .Y(n_86) );
AND2x2_ASAP7_75t_L g127 ( .A(n_87), .B(n_112), .Y(n_127) );
AND2x4_ASAP7_75t_L g139 ( .A(n_87), .B(n_137), .Y(n_139) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
INVx1_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
INVx1_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
AND2x2_ASAP7_75t_L g130 ( .A(n_88), .B(n_92), .Y(n_130) );
INVx2_ASAP7_75t_L g90 ( .A(n_89), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_89), .Y(n_96) );
OAI22x1_ASAP7_75t_L g98 ( .A1(n_89), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
INVxp67_ASAP7_75t_L g105 ( .A(n_91), .Y(n_105) );
AND2x4_ASAP7_75t_L g123 ( .A(n_91), .B(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g110 ( .A(n_92), .B(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g143 ( .A(n_94), .B(n_123), .Y(n_143) );
AND2x2_ASAP7_75t_L g156 ( .A(n_94), .B(n_110), .Y(n_156) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_97), .Y(n_94) );
AND2x2_ASAP7_75t_L g106 ( .A(n_95), .B(n_98), .Y(n_106) );
INVx2_ASAP7_75t_L g113 ( .A(n_95), .Y(n_113) );
BUFx2_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
AND2x4_ASAP7_75t_L g137 ( .A(n_97), .B(n_113), .Y(n_137) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx6_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x4_ASAP7_75t_L g116 ( .A(n_106), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g122 ( .A(n_106), .B(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
AND2x4_ASAP7_75t_L g146 ( .A(n_110), .B(n_137), .Y(n_146) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_111), .Y(n_118) );
AND2x4_ASAP7_75t_L g150 ( .A(n_112), .B(n_123), .Y(n_150) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx6_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g136 ( .A(n_123), .B(n_137), .Y(n_136) );
BUFx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx12f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x4_ASAP7_75t_L g153 ( .A(n_130), .B(n_137), .Y(n_153) );
AND2x4_ASAP7_75t_L g159 ( .A(n_130), .B(n_160), .Y(n_159) );
NAND4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_140), .C(n_147), .D(n_154), .Y(n_132) );
INVx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx8_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx8_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx6_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx5_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B1(n_167), .B2(n_177), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_167), .Y(n_177) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
CKINVDCx14_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g173 ( .A(n_172), .Y(n_173) );
INVx1_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
AND3x1_ASAP7_75t_SL g180 ( .A(n_181), .B(n_187), .C(n_190), .Y(n_180) );
INVxp67_ASAP7_75t_L g573 ( .A(n_181), .Y(n_573) );
CKINVDCx8_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_187), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_187), .A2(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g213 ( .A(n_188), .B(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_SL g578 ( .A(n_188), .B(n_190), .Y(n_578) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g224 ( .A(n_189), .B(n_215), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_190), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2x1p5_ASAP7_75t_L g221 ( .A(n_191), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND4xp75_ASAP7_75t_L g195 ( .A(n_196), .B(n_435), .C(n_480), .D(n_549), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2x1_ASAP7_75t_L g197 ( .A(n_198), .B(n_395), .Y(n_197) );
NOR3xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_351), .C(n_376), .Y(n_198) );
OAI222xp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_265), .B1(n_306), .B2(n_322), .C1(n_338), .C2(n_345), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_240), .Y(n_201) );
AND2x2_ASAP7_75t_L g560 ( .A(n_202), .B(n_374), .Y(n_560) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_204), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_204), .B(n_249), .Y(n_350) );
INVx3_ASAP7_75t_L g365 ( .A(n_204), .Y(n_365) );
AND2x2_ASAP7_75t_L g498 ( .A(n_204), .B(n_499), .Y(n_498) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_210), .B(n_236), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_205), .A2(n_206), .B1(n_251), .B2(n_257), .Y(n_250) );
AO21x2_ASAP7_75t_L g383 ( .A1(n_205), .A2(n_210), .B(n_236), .Y(n_383) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_207), .B(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx4f_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_209), .B(n_239), .Y(n_238) );
AND2x4_ASAP7_75t_L g271 ( .A(n_209), .B(n_239), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_219), .Y(n_210) );
INVx1_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_216), .Y(n_212) );
INVx1_ASAP7_75t_L g288 ( .A(n_213), .Y(n_288) );
OR2x6_ASAP7_75t_L g227 ( .A(n_214), .B(n_223), .Y(n_227) );
INVxp33_ASAP7_75t_L g318 ( .A(n_214), .Y(n_318) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_214), .Y(n_581) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g282 ( .A(n_215), .B(n_232), .Y(n_282) );
INVx1_ASAP7_75t_L g289 ( .A(n_216), .Y(n_289) );
BUFx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g223 ( .A(n_218), .Y(n_223) );
AND2x6_ASAP7_75t_L g279 ( .A(n_218), .B(n_230), .Y(n_279) );
INVxp67_ASAP7_75t_L g262 ( .A(n_220), .Y(n_262) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_224), .Y(n_220) );
INVx1_ASAP7_75t_L g319 ( .A(n_222), .Y(n_319) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .C(n_234), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g245 ( .A1(n_227), .A2(n_234), .B(n_246), .C(n_247), .Y(n_245) );
INVxp67_ASAP7_75t_L g252 ( .A(n_227), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_227), .A2(n_255), .B1(n_274), .B2(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g295 ( .A(n_227), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_227), .A2(n_234), .B(n_303), .C(n_304), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_SL g330 ( .A1(n_227), .A2(n_234), .B(n_331), .C(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g255 ( .A(n_229), .Y(n_255) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_234), .B(n_271), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_234), .A2(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g315 ( .A(n_234), .Y(n_315) );
INVx5_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_235), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_237), .Y(n_326) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g428 ( .A(n_240), .B(n_381), .Y(n_428) );
AND2x2_ASAP7_75t_L g430 ( .A(n_240), .B(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g465 ( .A(n_240), .Y(n_465) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_249), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g348 ( .A(n_242), .Y(n_348) );
INVx1_ASAP7_75t_L g367 ( .A(n_242), .Y(n_367) );
AND2x4_ASAP7_75t_L g374 ( .A(n_242), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_242), .B(n_312), .Y(n_390) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_242), .Y(n_499) );
INVx1_ASAP7_75t_L g509 ( .A(n_242), .Y(n_509) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_248), .Y(n_242) );
INVx2_ASAP7_75t_SL g296 ( .A(n_243), .Y(n_296) );
INVx1_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
INVx2_ASAP7_75t_L g362 ( .A(n_249), .Y(n_362) );
INVx1_ASAP7_75t_L g443 ( .A(n_249), .Y(n_443) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_258), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B1(n_263), .B2(n_264), .Y(n_258) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_264), .Y(n_564) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_267), .B(n_297), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_267), .B(n_324), .Y(n_418) );
INVx2_ASAP7_75t_L g439 ( .A(n_267), .Y(n_439) );
AND2x2_ASAP7_75t_L g447 ( .A(n_267), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_284), .Y(n_267) );
AND2x4_ASAP7_75t_L g337 ( .A(n_268), .B(n_285), .Y(n_337) );
INVx1_ASAP7_75t_L g344 ( .A(n_268), .Y(n_344) );
AND2x2_ASAP7_75t_L g520 ( .A(n_268), .B(n_325), .Y(n_520) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g358 ( .A(n_269), .B(n_285), .Y(n_358) );
INVx2_ASAP7_75t_L g394 ( .A(n_269), .Y(n_394) );
AND2x2_ASAP7_75t_L g473 ( .A(n_269), .B(n_325), .Y(n_473) );
NOR2x1_ASAP7_75t_SL g516 ( .A(n_269), .B(n_298), .Y(n_516) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_301), .B(n_305), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_283), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B1(n_280), .B2(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g356 ( .A(n_284), .Y(n_356) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g370 ( .A(n_285), .B(n_298), .Y(n_370) );
INVx1_ASAP7_75t_L g386 ( .A(n_285), .Y(n_386) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_285), .Y(n_494) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
NOR3xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .C(n_290), .Y(n_287) );
INVxp67_ASAP7_75t_L g582 ( .A(n_289), .Y(n_582) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_296), .A2(n_313), .B(n_321), .Y(n_312) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_296), .A2(n_313), .B(n_321), .Y(n_363) );
AND2x2_ASAP7_75t_L g357 ( .A(n_297), .B(n_358), .Y(n_357) );
OR2x6_ASAP7_75t_L g438 ( .A(n_297), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g476 ( .A(n_297), .B(n_473), .Y(n_476) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_298), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g405 ( .A(n_298), .Y(n_405) );
OR2x2_ASAP7_75t_L g411 ( .A(n_298), .B(n_325), .Y(n_411) );
AND2x4_ASAP7_75t_L g425 ( .A(n_298), .B(n_386), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_298), .B(n_394), .Y(n_426) );
OR2x6_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g470 ( .A(n_309), .B(n_389), .Y(n_470) );
BUFx2_ASAP7_75t_L g522 ( .A(n_309), .Y(n_522) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g553 ( .A(n_311), .B(n_465), .Y(n_553) );
INVx2_ASAP7_75t_L g347 ( .A(n_312), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_314), .B(n_320), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_334), .Y(n_322) );
AND2x2_ASAP7_75t_L g369 ( .A(n_323), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_SL g354 ( .A(n_324), .B(n_344), .Y(n_354) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g342 ( .A(n_325), .Y(n_342) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_325), .Y(n_448) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_325), .Y(n_515) );
INVx1_ASAP7_75t_L g555 ( .A(n_325), .Y(n_555) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_333), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
BUFx2_ASAP7_75t_L g469 ( .A(n_334), .Y(n_469) );
NOR2x1_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x4_ASAP7_75t_L g385 ( .A(n_335), .B(n_386), .Y(n_385) );
NOR2xp67_ASAP7_75t_SL g417 ( .A(n_335), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g490 ( .A(n_335), .B(n_473), .Y(n_490) );
AND2x4_ASAP7_75t_SL g493 ( .A(n_335), .B(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g542 ( .A(n_335), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g409 ( .A(n_336), .Y(n_409) );
INVx4_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g404 ( .A(n_337), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_337), .B(n_402), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_337), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_337), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g487 ( .A(n_341), .B(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g403 ( .A(n_342), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AND2x2_ASAP7_75t_L g521 ( .A(n_346), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g529 ( .A(n_346), .B(n_458), .Y(n_529) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g398 ( .A(n_347), .B(n_383), .Y(n_398) );
AND2x4_ASAP7_75t_L g431 ( .A(n_347), .B(n_365), .Y(n_431) );
INVx1_ASAP7_75t_L g548 ( .A(n_347), .Y(n_548) );
AND2x2_ASAP7_75t_L g434 ( .A(n_349), .B(n_374), .Y(n_434) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g455 ( .A(n_350), .B(n_390), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_359), .B1(n_368), .B2(n_371), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_357), .Y(n_352) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_353), .A2(n_422), .B1(n_530), .B2(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_354), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g423 ( .A(n_354), .B(n_355), .Y(n_423) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_354), .B(n_425), .Y(n_453) );
AOI211xp5_ASAP7_75t_SL g541 ( .A1(n_354), .A2(n_542), .B(n_544), .C(n_545), .Y(n_541) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_355), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_355), .B(n_401), .Y(n_527) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g432 ( .A(n_357), .Y(n_432) );
INVx2_ASAP7_75t_L g488 ( .A(n_358), .Y(n_488) );
AND2x2_ASAP7_75t_L g562 ( .A(n_358), .B(n_555), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_359), .A2(n_511), .B(n_517), .Y(n_510) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g497 ( .A(n_361), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g507 ( .A(n_361), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g414 ( .A(n_362), .B(n_367), .Y(n_414) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_362), .B(n_383), .Y(n_416) );
AND2x2_ASAP7_75t_L g458 ( .A(n_362), .B(n_383), .Y(n_458) );
INVx2_ASAP7_75t_L g375 ( .A(n_363), .Y(n_375) );
AND2x4_ASAP7_75t_L g381 ( .A(n_363), .B(n_382), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx3_ASAP7_75t_L g373 ( .A(n_365), .Y(n_373) );
INVx3_ASAP7_75t_L g379 ( .A(n_366), .Y(n_379) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_370), .A2(n_476), .B(n_552), .Y(n_556) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_373), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_373), .B(n_448), .Y(n_463) );
OR2x2_ASAP7_75t_L g478 ( .A(n_373), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g485 ( .A(n_373), .B(n_389), .Y(n_485) );
AND2x2_ASAP7_75t_L g441 ( .A(n_374), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g457 ( .A(n_374), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g474 ( .A(n_374), .B(n_443), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_384), .B1(n_387), .B2(n_391), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_379), .B(n_380), .Y(n_451) );
NOR2xp67_ASAP7_75t_SL g489 ( .A(n_379), .B(n_397), .Y(n_489) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_383), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g392 ( .A(n_385), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g456 ( .A(n_385), .B(n_402), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_385), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g559 ( .A(n_393), .B(n_425), .Y(n_559) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_394), .B(n_505), .Y(n_504) );
NOR2xp67_ASAP7_75t_SL g395 ( .A(n_396), .B(n_419), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_406), .C(n_415), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_397), .A2(n_450), .B(n_460), .C(n_464), .Y(n_459) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g539 ( .A(n_398), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g450 ( .A(n_402), .B(n_426), .Y(n_450) );
AND2x2_ASAP7_75t_L g537 ( .A(n_402), .B(n_516), .Y(n_537) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g505 ( .A(n_405), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_409), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g479 ( .A(n_414), .Y(n_479) );
NAND2xp33_ASAP7_75t_SL g415 ( .A(n_416), .B(n_417), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_427), .B1(n_429), .B2(n_432), .C(n_433), .Y(n_419) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .C(n_424), .D(n_426), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g538 ( .A(n_425), .B(n_501), .Y(n_538) );
INVx2_ASAP7_75t_L g544 ( .A(n_425), .Y(n_544) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_428), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g531 ( .A(n_431), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND4xp75_ASAP7_75t_L g436 ( .A(n_437), .B(n_459), .C(n_466), .D(n_475), .Y(n_436) );
OA211x2_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_444), .C(n_452), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_438), .B(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g532 ( .A(n_442), .Y(n_532) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g540 ( .A(n_443), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_445), .B(n_451), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g501 ( .A(n_448), .Y(n_501) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_456), .B2(n_457), .Y(n_452) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_456), .A2(n_507), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g535 ( .A(n_457), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_458), .B(n_548), .Y(n_547) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g533 ( .A(n_469), .Y(n_533) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_473), .B(n_493), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_474), .A2(n_537), .B1(n_559), .B2(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND3x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_523), .C(n_536), .Y(n_481) );
NOR3x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .C(n_510), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_491), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_489), .B2(n_490), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_500), .B1(n_502), .B2(n_506), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g554 ( .A(n_504), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_SL g543 ( .A(n_520), .Y(n_543) );
OAI21xp5_ASAP7_75t_SL g551 ( .A1(n_521), .A2(n_552), .B(n_554), .Y(n_551) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_534), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_528), .B1(n_530), .B2(n_533), .Y(n_524) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
O2A1O1Ixp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .C(n_541), .Y(n_536) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR2x1_ASAP7_75t_SL g549 ( .A(n_550), .B(n_557), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_556), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_558), .B(n_561), .Y(n_557) );
CKINVDCx16_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B1(n_574), .B2(n_576), .C1(n_579), .C2(n_583), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
endmodule