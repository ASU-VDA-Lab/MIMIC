module fake_netlist_1_814_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx3_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_6), .B(n_9), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_0), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_11), .B(n_0), .Y(n_18) );
INVxp67_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_17), .B(n_7), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_11), .B(n_1), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_14), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
NOR2x1p5_ASAP7_75t_L g25 ( .A(n_20), .B(n_12), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_19), .A2(n_16), .B1(n_15), .B2(n_13), .C(n_11), .Y(n_26) );
AND2x6_ASAP7_75t_L g27 ( .A(n_18), .B(n_13), .Y(n_27) );
OAI33xp33_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_19), .A3(n_22), .B1(n_23), .B2(n_15), .B3(n_21), .Y(n_28) );
NAND2xp33_ASAP7_75t_R g29 ( .A(n_24), .B(n_13), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_13), .B1(n_11), .B2(n_4), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_30), .B(n_26), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_28), .B(n_27), .Y(n_32) );
NAND2x1_ASAP7_75t_SL g33 ( .A(n_31), .B(n_29), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_27), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
BUFx12f_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AOI211xp5_ASAP7_75t_SL g37 ( .A1(n_35), .A2(n_2), .B(n_3), .C(n_10), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_33), .B(n_3), .Y(n_38) );
AND2x2_ASAP7_75t_L g39 ( .A(n_36), .B(n_34), .Y(n_39) );
INVx2_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
AOI22xp33_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_38), .B1(n_33), .B2(n_37), .Y(n_41) );
endmodule