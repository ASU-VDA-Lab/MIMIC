module fake_jpeg_3956_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_34),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_15),
.B1(n_28),
.B2(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_50),
.B1(n_63),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_18),
.B1(n_15),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_57),
.B1(n_31),
.B2(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_15),
.B1(n_28),
.B2(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_22),
.B(n_21),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_22),
.CON(n_63),
.SN(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_80),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_19),
.B1(n_31),
.B2(n_17),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_61),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_22),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_77),
.B(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_24),
.B1(n_17),
.B2(n_23),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_54),
.B(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_64),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_59),
.B1(n_54),
.B2(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_43),
.B1(n_56),
.B2(n_60),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_80),
.B1(n_29),
.B2(n_25),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_21),
.B(n_29),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_106),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_60),
.C(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_52),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_113),
.B1(n_122),
.B2(n_127),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_81),
.B1(n_82),
.B2(n_67),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_76),
.B1(n_81),
.B2(n_69),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_126),
.B1(n_107),
.B2(n_108),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_81),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_133),
.B(n_92),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_82),
.B1(n_56),
.B2(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_127),
.B1(n_91),
.B2(n_102),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_125),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_88),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_77),
.B1(n_56),
.B2(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_21),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_139),
.B(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_98),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_124),
.B(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_133),
.A2(n_117),
.B(n_130),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_122),
.C(n_118),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_145),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_146),
.B(n_156),
.C(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_88),
.B1(n_102),
.B2(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_157),
.B1(n_122),
.B2(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_95),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_95),
.B(n_103),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_101),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_112),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_167),
.C(n_180),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_115),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_169),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_113),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_113),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_155),
.CI(n_157),
.CON(n_171),
.SN(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_177),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_131),
.B1(n_121),
.B2(n_128),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_176),
.B(n_101),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

XOR2x1_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_128),
.Y(n_176)
);

AOI22x1_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_126),
.B1(n_120),
.B2(n_121),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_142),
.B1(n_141),
.B2(n_158),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_101),
.B1(n_29),
.B2(n_25),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_182),
.A2(n_151),
.B1(n_153),
.B2(n_148),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_188),
.B1(n_203),
.B2(n_168),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_149),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_198),
.B(n_182),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_138),
.B1(n_146),
.B2(n_137),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_202),
.B(n_171),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_141),
.C(n_152),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_142),
.C(n_116),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.C(n_160),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_132),
.C(n_99),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_177),
.B(n_10),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_64),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_201),
.B(n_199),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_29),
.B1(n_25),
.B2(n_65),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_64),
.B1(n_58),
.B2(n_65),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_213),
.B(n_14),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_208),
.C(n_212),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_178),
.C(n_170),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_185),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_173),
.C(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_174),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_190),
.A2(n_168),
.B(n_162),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_214),
.A2(n_218),
.B1(n_7),
.B2(n_13),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_221),
.B1(n_202),
.B2(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_221),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_65),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_65),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_228),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_185),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_232),
.C(n_233),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_186),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_58),
.C(n_1),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_58),
.C(n_1),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_206),
.C(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_247),
.C(n_11),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_212),
.B1(n_210),
.B2(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_243),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_7),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_8),
.B(n_13),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_8),
.Y(n_247)
);

NAND4xp25_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_0),
.C(n_2),
.D(n_3),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_226),
.B1(n_225),
.B2(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_222),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_252),
.B(n_254),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_0),
.C(n_2),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_256),
.C(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_3),
.C(n_4),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_237),
.B(n_245),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_259),
.B(n_262),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_248),
.C(n_11),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_12),
.C(n_13),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_9),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_3),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_4),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_256),
.B(n_12),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_263),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_265),
.B(n_14),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_14),
.B(n_4),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_271),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_5),
.Y(n_278)
);


endmodule