module fake_jpeg_22393_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_41),
.CON(n_50),
.SN(n_50)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_21),
.B1(n_23),
.B2(n_35),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_40),
.B1(n_36),
.B2(n_31),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_40),
.B1(n_23),
.B2(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_83),
.B1(n_36),
.B2(n_31),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_23),
.B1(n_21),
.B2(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_74),
.B1(n_53),
.B2(n_60),
.Y(n_98)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_23),
.B1(n_21),
.B2(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_34),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_43),
.B1(n_57),
.B2(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_102),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_52),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_0),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_99),
.B1(n_107),
.B2(n_110),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_109),
.B1(n_112),
.B2(n_24),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_50),
.B(n_52),
.C(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_38),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_24),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_67),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_38),
.C(n_22),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_113),
.C(n_24),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_43),
.B1(n_22),
.B2(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_85),
.B1(n_70),
.B2(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_55),
.B1(n_58),
.B2(n_37),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_80),
.B1(n_82),
.B2(n_76),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_117),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_100),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_34),
.B(n_41),
.C(n_18),
.Y(n_160)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_12),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_27),
.B(n_30),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_66),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_26),
.C(n_102),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_66),
.Y(n_136)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_29),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_33),
.Y(n_158)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_92),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_117),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_164),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_106),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_158),
.B(n_160),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_96),
.A3(n_105),
.B1(n_114),
.B2(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_163),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_108),
.B1(n_93),
.B2(n_91),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_134),
.B1(n_140),
.B2(n_122),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_19),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_135),
.C(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_153),
.C(n_158),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

AOI22x1_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_126),
.B1(n_121),
.B2(n_115),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_147),
.B1(n_33),
.B2(n_32),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_118),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_126),
.B1(n_129),
.B2(n_116),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_181),
.B1(n_188),
.B2(n_191),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_182),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_143),
.Y(n_182)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_219)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_142),
.B1(n_145),
.B2(n_164),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_128),
.B(n_127),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_190),
.B(n_192),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_118),
.C(n_128),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_141),
.B1(n_139),
.B2(n_133),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_144),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_141),
.C(n_139),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_167),
.B(n_161),
.Y(n_206)
);

BUFx4f_ASAP7_75t_SL g194 ( 
.A(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_154),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_195),
.B(n_201),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_165),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_197),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_171),
.B(n_154),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_159),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_204),
.B(n_210),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_203),
.C(n_214),
.Y(n_224)
);

XOR2x2_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_153),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_181),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_187),
.B(n_186),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_172),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_167),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_152),
.B(n_166),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_27),
.B(n_30),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_183),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_147),
.B1(n_133),
.B2(n_130),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_101),
.B1(n_93),
.B2(n_86),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_241),
.B1(n_216),
.B2(n_30),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_172),
.C(n_91),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_239),
.C(n_197),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_230),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_193),
.C(n_184),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_84),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_240),
.B1(n_242),
.B2(n_216),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

AOI21x1_ASAP7_75t_SL g234 ( 
.A1(n_198),
.A2(n_1),
.B(n_2),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_101),
.C(n_86),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_237),
.B(n_215),
.CI(n_203),
.CON(n_243),
.SN(n_243)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_250),
.C(n_261),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_212),
.B1(n_216),
.B2(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_245),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_196),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_249),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_205),
.C(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_20),
.B(n_32),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_79),
.B1(n_27),
.B2(n_15),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_260),
.B1(n_262),
.B2(n_28),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_226),
.A2(n_79),
.B1(n_15),
.B2(n_19),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_33),
.C(n_32),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_271),
.B(n_278),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_269),
.B1(n_275),
.B2(n_276),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_223),
.B(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_222),
.B1(n_241),
.B2(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_224),
.C(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.C(n_243),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_238),
.C(n_25),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_25),
.B1(n_20),
.B2(n_18),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_243),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_293),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_246),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_285),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_249),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_286),
.B(n_14),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_251),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_6),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_290),
.B(n_291),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_257),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_7),
.B(n_9),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_6),
.B(n_9),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_280),
.B1(n_292),
.B2(n_271),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_276),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_299),
.B(n_304),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_270),
.B1(n_265),
.B2(n_274),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_7),
.B1(n_9),
.B2(n_8),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_266),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_2),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_6),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_7),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_8),
.C(n_14),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_314),
.C(n_296),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_8),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_311),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_14),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_315),
.B(n_300),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_4),
.B(n_5),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_306),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_3),
.B(n_4),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_322),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_325),
.C(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_320),
.C(n_308),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_324),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_5),
.B1(n_323),
.B2(n_325),
.Y(n_332)
);


endmodule