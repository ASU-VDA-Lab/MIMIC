module fake_aes_3800_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI22xp33_ASAP7_75t_R g11 ( .A1(n_6), .A2(n_4), .B1(n_2), .B2(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_7), .B(n_0), .Y(n_14) );
NOR2xp67_ASAP7_75t_L g15 ( .A(n_5), .B(n_1), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_10), .B(n_4), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_12), .B(n_2), .Y(n_17) );
BUFx12f_ASAP7_75t_SL g18 ( .A(n_14), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_14), .B(n_3), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx6_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_23), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_19), .B1(n_16), .B2(n_14), .Y(n_27) );
NAND2xp33_ASAP7_75t_SL g28 ( .A(n_26), .B(n_25), .Y(n_28) );
AOI211xp5_ASAP7_75t_SL g29 ( .A1(n_27), .A2(n_15), .B(n_16), .C(n_11), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_13), .Y(n_30) );
NOR2xp67_ASAP7_75t_SL g31 ( .A(n_28), .B(n_21), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_28), .B(n_12), .Y(n_32) );
NAND2xp5_ASAP7_75t_SL g33 ( .A(n_32), .B(n_16), .Y(n_33) );
INVxp67_ASAP7_75t_SL g34 ( .A(n_31), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_34), .B(n_30), .Y(n_35) );
AOI322xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_33), .A3(n_11), .B1(n_5), .B2(n_3), .C1(n_8), .C2(n_21), .Y(n_36) );
endmodule