module fake_jpeg_2957_n_128 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_43),
.Y(n_61)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_27),
.Y(n_58)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_12),
.B(n_23),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_12),
.B1(n_16),
.B2(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_48),
.B1(n_27),
.B2(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_17),
.B1(n_27),
.B2(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_17),
.B1(n_22),
.B2(n_25),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_37),
.B1(n_29),
.B2(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_70),
.B1(n_78),
.B2(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_8),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_6),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_79),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_10),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_51),
.B(n_11),
.C(n_54),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_90),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_72),
.B1(n_63),
.B2(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_53),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_60),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_60),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_87),
.B(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_98),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_77),
.B1(n_67),
.B2(n_52),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_100),
.B1(n_82),
.B2(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_71),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_52),
.B1(n_47),
.B2(n_3),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_96),
.B1(n_97),
.B2(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_109),
.B1(n_108),
.B2(n_105),
.Y(n_114)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_103),
.A3(n_93),
.B1(n_86),
.B2(n_107),
.C(n_84),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_117),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_86),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_112),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_110),
.C(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_124),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_120),
.B(n_3),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_47),
.Y(n_128)
);


endmodule