module fake_jpeg_13436_n_64 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

AND2x2_ASAP7_75t_SL g9 ( 
.A(n_0),
.B(n_7),
.Y(n_9)
);

BUFx4f_ASAP7_75t_SL g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_1),
.B1(n_3),
.B2(n_8),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_11),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_16),
.B1(n_14),
.B2(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_15),
.B2(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_11),
.B(n_22),
.C(n_20),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_29),
.C(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_10),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_20),
.B(n_22),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_32),
.C(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_38),
.C(n_25),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_36),
.B(n_40),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

OAI211xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_53),
.B(n_43),
.C(n_33),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_46),
.B2(n_40),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_53),
.B(n_51),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.C(n_34),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B(n_5),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_4),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_6),
.B(n_7),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_1),
.B1(n_10),
.B2(n_62),
.C(n_61),
.Y(n_64)
);


endmodule