module fake_jpeg_2504_n_196 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_82),
.Y(n_97)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_74),
.Y(n_92)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_54),
.B1(n_57),
.B2(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_96),
.B1(n_99),
.B2(n_73),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_59),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_55),
.C(n_53),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_1),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_59),
.B1(n_61),
.B2(n_52),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_59),
.B1(n_61),
.B2(n_73),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_74),
.A3(n_56),
.B1(n_73),
.B2(n_81),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_108),
.B(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_113),
.B1(n_58),
.B2(n_94),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_80),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_66),
.B(n_67),
.C(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_57),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_94),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_80),
.B1(n_76),
.B2(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_1),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_2),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_6),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_107),
.B1(n_101),
.B2(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_136),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_98),
.B1(n_84),
.B2(n_58),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_129),
.B1(n_130),
.B2(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_137),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_107),
.B1(n_100),
.B2(n_108),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_70),
.CI(n_5),
.CON(n_132),
.SN(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_65),
.C(n_23),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_135),
.C(n_14),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_22),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_9),
.B(n_10),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_13),
.B(n_14),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_26),
.C(n_27),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_157),
.B(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_154),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_15),
.B(n_16),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_48),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_15),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_17),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_19),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_24),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_161),
.A2(n_34),
.B(n_35),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_167),
.C(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_47),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_39),
.C(n_40),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_43),
.B(n_46),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_168),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_167),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_145),
.B1(n_159),
.B2(n_169),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_181),
.B1(n_159),
.B2(n_171),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_149),
.B(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_172),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_185),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_186),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_148),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_182),
.B1(n_162),
.B2(n_179),
.Y(n_190)
);

AOI31xp33_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_191),
.A3(n_163),
.B(n_162),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_180),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_189),
.B(n_165),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_151),
.Y(n_196)
);


endmodule