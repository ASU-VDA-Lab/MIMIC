module fake_jpeg_17344_n_126 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_27),
.B(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_3),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.C(n_18),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_3),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_6),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_53),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_34),
.B1(n_29),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_24),
.B(n_23),
.C(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_64),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_16),
.B1(n_19),
.B2(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_26),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_26),
.B1(n_11),
.B2(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_55),
.B1(n_62),
.B2(n_47),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_42),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_51),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_52),
.B(n_50),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_72),
.C(n_67),
.Y(n_102)
);

OAI31xp33_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_59),
.A3(n_56),
.B(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_96),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_48),
.B1(n_55),
.B2(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_62),
.B1(n_69),
.B2(n_77),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_107),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_78),
.B1(n_68),
.B2(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_103),
.B(n_95),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_96),
.C(n_85),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_88),
.B1(n_84),
.B2(n_87),
.Y(n_119)
);

FAx1_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_93),
.CI(n_88),
.CON(n_109),
.SN(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_81),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_92),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_107),
.C(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_117),
.B1(n_83),
.B2(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_106),
.Y(n_117)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_112),
.B(n_109),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_75),
.B(n_83),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_122),
.C(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_121),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_124),
.Y(n_126)
);


endmodule