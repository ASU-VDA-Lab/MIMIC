module fake_jpeg_23699_n_32 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_32);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_0),
.B1(n_5),
.B2(n_10),
.Y(n_19)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_7),
.A3(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_18),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_6),
.A3(n_15),
.B1(n_2),
.B2(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_23),
.B(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_27),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_25),
.C(n_26),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_29),
.C(n_2),
.Y(n_32)
);


endmodule