module fake_jpeg_9204_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_16),
.B(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_52),
.B1(n_34),
.B2(n_38),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_25),
.C(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_16),
.B1(n_15),
.B2(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_23),
.B1(n_22),
.B2(n_31),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_63),
.B1(n_74),
.B2(n_75),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_73),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_40),
.B1(n_37),
.B2(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_42),
.B1(n_22),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_77)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_57),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_11),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_45),
.C(n_30),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_29),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_45),
.B1(n_55),
.B2(n_50),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_85),
.B1(n_90),
.B2(n_97),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_61),
.B(n_57),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_50),
.B1(n_40),
.B2(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_43),
.B1(n_49),
.B2(n_47),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_93),
.B(n_14),
.Y(n_107)
);

AOI22x1_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_67),
.B1(n_36),
.B2(n_29),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_36),
.B1(n_49),
.B2(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_102),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_83),
.B(n_84),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_68),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_80),
.C(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_70),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_9),
.B(n_13),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_71),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_36),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_87),
.B1(n_98),
.B2(n_84),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_114),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_10),
.C(n_14),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_98),
.B1(n_81),
.B2(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_122),
.B1(n_65),
.B2(n_28),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_111),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_89),
.B(n_36),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_125),
.B(n_8),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_110),
.B1(n_109),
.B2(n_102),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_47),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_103),
.B1(n_112),
.B2(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_128),
.B1(n_65),
.B2(n_124),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_137),
.B(n_139),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_1),
.B(n_2),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_120),
.C(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.C(n_138),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_140),
.Y(n_156)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_122),
.B1(n_125),
.B2(n_7),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_150),
.C(n_147),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_155),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_131),
.B1(n_8),
.B2(n_9),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_159),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_147),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_4),
.B(n_5),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_150),
.B(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_152),
.B(n_10),
.C(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_4),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_159),
.B(n_160),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_168),
.C(n_158),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_172),
.Y(n_174)
);


endmodule