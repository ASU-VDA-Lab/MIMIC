module fake_netlist_6_599_n_3833 (n_992, n_52, n_591, n_435, n_1115, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_1202, n_881, n_1199, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_1189, n_223, n_278, n_1079, n_341, n_362, n_1212, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_1103, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_1061, n_384, n_297, n_595, n_627, n_1203, n_524, n_342, n_77, n_820, n_1044, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_1217, n_160, n_751, n_449, n_131, n_749, n_1208, n_798, n_188, n_1164, n_310, n_509, n_186, n_245, n_1209, n_0, n_368, n_575, n_994, n_1072, n_677, n_969, n_988, n_805, n_1151, n_396, n_495, n_1065, n_815, n_350, n_1100, n_1214, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_1128, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_1071, n_628, n_1067, n_1204, n_1160, n_883, n_557, n_823, n_1132, n_349, n_643, n_233, n_617, n_698, n_898, n_1074, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_1138, n_893, n_214, n_925, n_485, n_1099, n_67, n_15, n_1026, n_443, n_1101, n_246, n_892, n_768, n_1097, n_38, n_471, n_289, n_935, n_1192, n_421, n_781, n_424, n_789, n_615, n_1130, n_59, n_181, n_1127, n_182, n_238, n_1095, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_1120, n_597, n_685, n_280, n_287, n_832, n_353, n_1187, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_1139, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_1172, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_1105, n_1206, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_1140, n_378, n_413, n_1196, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_1114, n_56, n_763, n_1057, n_1147, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_1143, n_536, n_895, n_1126, n_866, n_622, n_147, n_191, n_340, n_710, n_1108, n_387, n_1182, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_1119, n_73, n_581, n_428, n_761, n_785, n_746, n_1205, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_1056, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_1163, n_1173, n_1180, n_1116, n_611, n_943, n_156, n_1168, n_491, n_1219, n_1216, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_1174, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_1221, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_1094, n_1176, n_1190, n_494, n_539, n_493, n_397, n_155, n_1022, n_1083, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_1112, n_454, n_34, n_218, n_1213, n_638, n_70, n_234, n_1181, n_910, n_1211, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_1117, n_1087, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_1049, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1043, n_1011, n_118, n_224, n_48, n_926, n_927, n_1215, n_25, n_93, n_839, n_986, n_80, n_734, n_1088, n_708, n_196, n_919, n_1081, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_1084, n_107, n_1171, n_1104, n_907, n_854, n_6, n_1058, n_417, n_14, n_446, n_498, n_662, n_1122, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_1109, n_921, n_185, n_712, n_1183, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_1193, n_1148, n_293, n_1054, n_31, n_334, n_559, n_53, n_370, n_1161, n_44, n_458, n_1070, n_1085, n_232, n_650, n_998, n_16, n_1046, n_163, n_717, n_46, n_1145, n_330, n_771, n_1121, n_1152, n_470, n_475, n_924, n_1102, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_1149, n_564, n_1178, n_98, n_260, n_265, n_313, n_451, n_624, n_1184, n_824, n_962, n_1073, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_1195, n_356, n_577, n_166, n_936, n_184, n_552, n_1186, n_1062, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_1090, n_745, n_654, n_323, n_829, n_1156, n_606, n_393, n_818, n_984, n_411, n_1142, n_503, n_716, n_152, n_623, n_1048, n_1123, n_92, n_884, n_1201, n_599, n_1222, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_1078, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_1137, n_433, n_500, n_1218, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_1144, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_1162, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_1068, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_1075, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_1198, n_237, n_584, n_1110, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_1155, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_1133, n_635, n_95, n_787, n_1194, n_311, n_10, n_1064, n_403, n_1080, n_723, n_253, n_634, n_1051, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_1141, n_1146, n_249, n_201, n_386, n_764, n_1039, n_1220, n_556, n_159, n_1034, n_1086, n_1066, n_157, n_162, n_692, n_733, n_1158, n_754, n_1136, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_1125, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_1107, n_560, n_1014, n_753, n_642, n_995, n_276, n_1159, n_569, n_1092, n_441, n_221, n_811, n_882, n_1060, n_444, n_586, n_423, n_146, n_737, n_318, n_1207, n_1111, n_303, n_1223, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_1053, n_530, n_277, n_520, n_1029, n_418, n_1093, n_113, n_618, n_1055, n_790, n_1106, n_582, n_4, n_199, n_1167, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_1153, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_1210, n_679, n_1069, n_5, n_1185, n_453, n_612, n_633, n_1170, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1047, n_1010, n_355, n_1165, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_1166, n_431, n_90, n_347, n_812, n_24, n_459, n_1131, n_54, n_1052, n_502, n_1175, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_1045, n_786, n_670, n_203, n_286, n_1224, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_1089, n_1135, n_1169, n_1179, n_75, n_401, n_324, n_743, n_766, n_816, n_1157, n_335, n_430, n_1002, n_463, n_1188, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_1096, n_1063, n_729, n_1091, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_1124, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_1200, n_1059, n_1197, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_1077, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_1082, n_259, n_1154, n_177, n_1113, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_1098, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_1050, n_379, n_170, n_778, n_1025, n_1134, n_1177, n_332, n_891, n_336, n_1150, n_12, n_398, n_410, n_1129, n_1191, n_566, n_554, n_602, n_1013, n_1023, n_1076, n_1118, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_3833);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1115;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_881;
input n_1199;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_1189;
input n_223;
input n_278;
input n_1079;
input n_341;
input n_362;
input n_1212;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_1103;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_1061;
input n_384;
input n_297;
input n_595;
input n_627;
input n_1203;
input n_524;
input n_342;
input n_77;
input n_820;
input n_1044;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1217;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_1208;
input n_798;
input n_188;
input n_1164;
input n_310;
input n_509;
input n_186;
input n_245;
input n_1209;
input n_0;
input n_368;
input n_575;
input n_994;
input n_1072;
input n_677;
input n_969;
input n_988;
input n_805;
input n_1151;
input n_396;
input n_495;
input n_1065;
input n_815;
input n_350;
input n_1100;
input n_1214;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_1128;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_1071;
input n_628;
input n_1067;
input n_1204;
input n_1160;
input n_883;
input n_557;
input n_823;
input n_1132;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1074;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_1138;
input n_893;
input n_214;
input n_925;
input n_485;
input n_1099;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_1101;
input n_246;
input n_892;
input n_768;
input n_1097;
input n_38;
input n_471;
input n_289;
input n_935;
input n_1192;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_1130;
input n_59;
input n_181;
input n_1127;
input n_182;
input n_238;
input n_1095;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_1120;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_1187;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_1139;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_1172;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_1105;
input n_1206;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_1140;
input n_378;
input n_413;
input n_1196;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1057;
input n_1147;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_1143;
input n_536;
input n_895;
input n_1126;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_1108;
input n_387;
input n_1182;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_1119;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_1205;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_1163;
input n_1173;
input n_1180;
input n_1116;
input n_611;
input n_943;
input n_156;
input n_1168;
input n_491;
input n_1219;
input n_1216;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_1174;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_1221;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_1094;
input n_1176;
input n_1190;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_1083;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_1112;
input n_454;
input n_34;
input n_218;
input n_1213;
input n_638;
input n_70;
input n_234;
input n_1181;
input n_910;
input n_1211;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_1117;
input n_1087;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_1049;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1043;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_1088;
input n_708;
input n_196;
input n_919;
input n_1081;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_1084;
input n_107;
input n_1171;
input n_1104;
input n_907;
input n_854;
input n_6;
input n_1058;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_1122;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_1109;
input n_921;
input n_185;
input n_712;
input n_1183;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_1193;
input n_1148;
input n_293;
input n_1054;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_1161;
input n_44;
input n_458;
input n_1070;
input n_1085;
input n_232;
input n_650;
input n_998;
input n_16;
input n_1046;
input n_163;
input n_717;
input n_46;
input n_1145;
input n_330;
input n_771;
input n_1121;
input n_1152;
input n_470;
input n_475;
input n_924;
input n_1102;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_1149;
input n_564;
input n_1178;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_1184;
input n_824;
input n_962;
input n_1073;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_1195;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_1186;
input n_1062;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_1090;
input n_745;
input n_654;
input n_323;
input n_829;
input n_1156;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_1142;
input n_503;
input n_716;
input n_152;
input n_623;
input n_1048;
input n_1123;
input n_92;
input n_884;
input n_1201;
input n_599;
input n_1222;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_1078;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_1137;
input n_433;
input n_500;
input n_1218;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_1144;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_1162;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_1068;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_1075;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_1198;
input n_237;
input n_584;
input n_1110;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_1155;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_787;
input n_1194;
input n_311;
input n_10;
input n_1064;
input n_403;
input n_1080;
input n_723;
input n_253;
input n_634;
input n_1051;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_1141;
input n_1146;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_1220;
input n_556;
input n_159;
input n_1034;
input n_1086;
input n_1066;
input n_157;
input n_162;
input n_692;
input n_733;
input n_1158;
input n_754;
input n_1136;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_1125;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_1107;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_569;
input n_1092;
input n_441;
input n_221;
input n_811;
input n_882;
input n_1060;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_1207;
input n_1111;
input n_303;
input n_1223;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_1053;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_1093;
input n_113;
input n_618;
input n_1055;
input n_790;
input n_1106;
input n_582;
input n_4;
input n_199;
input n_1167;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_1153;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_1210;
input n_679;
input n_1069;
input n_5;
input n_1185;
input n_453;
input n_612;
input n_633;
input n_1170;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1047;
input n_1010;
input n_355;
input n_1165;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_1166;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_1131;
input n_54;
input n_1052;
input n_502;
input n_1175;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_1045;
input n_786;
input n_670;
input n_203;
input n_286;
input n_1224;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_1089;
input n_1135;
input n_1169;
input n_1179;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_1157;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_1188;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_1096;
input n_1063;
input n_729;
input n_1091;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_1124;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_1200;
input n_1059;
input n_1197;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_1077;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_1082;
input n_259;
input n_1154;
input n_177;
input n_1113;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_1098;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_1050;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_1134;
input n_1177;
input n_332;
input n_891;
input n_336;
input n_1150;
input n_12;
input n_398;
input n_410;
input n_1129;
input n_1191;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_3833;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_3392;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_3152;
wire n_3579;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1581;
wire n_1237;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1348;
wire n_2260;
wire n_1387;
wire n_3222;
wire n_1708;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_2647;
wire n_2997;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_1555;
wire n_2211;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_3106;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_3316;
wire n_2212;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_2729;
wire n_3063;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1471;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_1658;
wire n_2593;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_1967;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_1441;
wire n_3373;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_3732;
wire n_1302;
wire n_1599;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_3716;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_2068;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1950;
wire n_1726;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_3273;
wire n_2311;
wire n_1386;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_3691;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_2347;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_3415;
wire n_1588;
wire n_3785;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_3510;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_2271;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3337;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3431;
wire n_3450;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1627;
wire n_1295;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_1952;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_1932;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_2316;
wire n_1771;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_2239;
wire n_1707;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_2134;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_2424;
wire n_2296;
wire n_1604;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_1398;
wire n_2682;
wire n_3032;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_1837;
wire n_2218;
wire n_1314;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_3755;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_2329;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_2250;
wire n_1951;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_2990;
wire n_1775;
wire n_1286;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_2928;
wire n_2249;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_2315;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_3663;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1832;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_2201;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_3276;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_3548;
wire n_3767;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_3230;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_2404;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_3238;
wire n_3529;
wire n_2235;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_3819;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_2699;
wire n_2046;
wire n_2272;
wire n_1828;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_2258;
wire n_1485;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_3712;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_2533;
wire n_1672;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_3506;
wire n_2398;
wire n_1559;
wire n_1928;
wire n_1725;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3818;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2923;
wire n_2888;
wire n_2715;
wire n_2793;
wire n_1804;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_3308;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_2358;
wire n_1401;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_3034;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3567;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_1848;
wire n_1785;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1570;
wire n_1702;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_3573;
wire n_1944;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_3494;
wire n_1737;
wire n_2430;
wire n_1464;
wire n_1414;
wire n_3486;
wire n_2649;
wire n_2721;
wire n_3556;
wire n_2034;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_2437;
wire n_2444;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_2609;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_2071;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_3374;
wire n_3786;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_2909;
wire n_2248;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_2221;
wire n_1629;
wire n_2055;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_3444;
wire n_2553;
wire n_3059;
wire n_2038;
wire n_2891;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_2477;
wire n_1805;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3433;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3815;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_3504;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1097),
.Y(n_1225)
);

BUFx10_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

CKINVDCx16_ASAP7_75t_R g1227 ( 
.A(n_1076),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_602),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1162),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_315),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1119),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1112),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1078),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_381),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1004),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1218),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_988),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_968),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1047),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1080),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_230),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_941),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1037),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_462),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_784),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_180),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1045),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1082),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_424),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1140),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1085),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_584),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_717),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_709),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1004),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1053),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_624),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1111),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_185),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_674),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_242),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_942),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_915),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_446),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_236),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_123),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1167),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1064),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_667),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1083),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1127),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_129),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_667),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_154),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_25),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_563),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_15),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_488),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1172),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_828),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_144),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1151),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_857),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_605),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_249),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_967),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_238),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_768),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_48),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_529),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_435),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1052),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_924),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_685),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1175),
.Y(n_1295)
);

BUFx8_ASAP7_75t_SL g1296 ( 
.A(n_811),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_488),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1101),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_534),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1040),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_14),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1063),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_869),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1165),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_865),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_810),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_836),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_837),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1166),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_286),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1161),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_993),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_864),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_552),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_986),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1003),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_262),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_427),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_733),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1125),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_278),
.Y(n_1321)
);

BUFx5_ASAP7_75t_L g1322 ( 
.A(n_1147),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_961),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_743),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_1104),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1143),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1157),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_436),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1149),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_786),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_971),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_901),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_462),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_504),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1067),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1122),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_629),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1219),
.Y(n_1338)
);

CKINVDCx14_ASAP7_75t_R g1339 ( 
.A(n_1055),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1176),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_117),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_625),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_197),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_877),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_904),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_616),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_854),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1173),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_969),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_835),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_770),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1120),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_655),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_23),
.Y(n_1354)
);

CKINVDCx16_ASAP7_75t_R g1355 ( 
.A(n_65),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_497),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1114),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1178),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1193),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_959),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_607),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_630),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_32),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1168),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_773),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1138),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_785),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_898),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_516),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_220),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1099),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1058),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1125),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_104),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_332),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_819),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_925),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_927),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_148),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_958),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1040),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_255),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_876),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_442),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_291),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1164),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_933),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1058),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_552),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_454),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_731),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_179),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_894),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_469),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1195),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_931),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1222),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1072),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_418),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1044),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_838),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_919),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_226),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_345),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_63),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_448),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1114),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_772),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_897),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_899),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_217),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1117),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1092),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1153),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_515),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_190),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_708),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_321),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_845),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_280),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_180),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_961),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_366),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_510),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_852),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_896),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_503),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1154),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_944),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_827),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_665),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_757),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_607),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1098),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_609),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_345),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_271),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_991),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_839),
.Y(n_1439)
);

BUFx5_ASAP7_75t_L g1440 ( 
.A(n_509),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_742),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1119),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1059),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1014),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_808),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_328),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_700),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_129),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1009),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_979),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1073),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_579),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_837),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_266),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_602),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_913),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_895),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_980),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_976),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_851),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_487),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1198),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1209),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_984),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_209),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1215),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_770),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1146),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_146),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_218),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_303),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1126),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_812),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_22),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1057),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1131),
.Y(n_1476)
);

BUFx5_ASAP7_75t_L g1477 ( 
.A(n_791),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_176),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_370),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1105),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_779),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1001),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_666),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_194),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_564),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_908),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1096),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1203),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1038),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1214),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_368),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_717),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_599),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_336),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1191),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_912),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1113),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_735),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_789),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_584),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1136),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1145),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_995),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_185),
.Y(n_1504)
);

BUFx10_ASAP7_75t_L g1505 ( 
.A(n_455),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_489),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_983),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1068),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_625),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1023),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_509),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1072),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_626),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1188),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_741),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_876),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_890),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_853),
.Y(n_1518)
);

BUFx10_ASAP7_75t_L g1519 ( 
.A(n_1171),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_305),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_154),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_180),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_960),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_640),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_856),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_484),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_366),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_829),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_642),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1212),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_502),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_990),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_795),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1051),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_841),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_756),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_872),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_699),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_545),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_714),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1055),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1014),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_793),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_909),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1005),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1090),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1161),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_589),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1118),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_279),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_718),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1196),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1223),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1089),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_874),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_235),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_951),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_764),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1042),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_242),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_969),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_809),
.B(n_146),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1205),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1130),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_769),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1088),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1010),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_815),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_1033),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_575),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1150),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_954),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_940),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1093),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1163),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_457),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_606),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1159),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_58),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1170),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_873),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1138),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_937),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_140),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_677),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1074),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1211),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_248),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1169),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_875),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_26),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_269),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_515),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_505),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_415),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_504),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_191),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_994),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1141),
.Y(n_1599)
);

BUFx10_ASAP7_75t_L g1600 ( 
.A(n_1142),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_251),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_211),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_865),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_763),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1220),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_71),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1086),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_759),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_805),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_299),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_262),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1124),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_547),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_663),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1020),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_481),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_996),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_106),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_393),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_847),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_537),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_780),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_224),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_855),
.Y(n_1624)
);

BUFx10_ASAP7_75t_L g1625 ( 
.A(n_457),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1148),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_37),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_781),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_981),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_479),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_902),
.Y(n_1631)
);

BUFx10_ASAP7_75t_L g1632 ( 
.A(n_824),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_45),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_451),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_765),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_985),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_223),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_914),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1077),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_794),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_600),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1156),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1106),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_881),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_771),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1174),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1034),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1062),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_788),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_208),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_847),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_885),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1135),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_232),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_722),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_450),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1108),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_712),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1075),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_167),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_964),
.Y(n_1661)
);

BUFx10_ASAP7_75t_L g1662 ( 
.A(n_1026),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1197),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_365),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_707),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_758),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_479),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1110),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1183),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1066),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_900),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1070),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1180),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_987),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_893),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1123),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_3),
.Y(n_1677)
);

CKINVDCx14_ASAP7_75t_R g1678 ( 
.A(n_955),
.Y(n_1678)
);

CKINVDCx16_ASAP7_75t_R g1679 ( 
.A(n_1139),
.Y(n_1679)
);

CKINVDCx14_ASAP7_75t_R g1680 ( 
.A(n_1141),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_356),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_498),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_734),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_938),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_378),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_937),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1155),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1061),
.Y(n_1688)
);

CKINVDCx16_ASAP7_75t_R g1689 ( 
.A(n_804),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_653),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1049),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_681),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_697),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1158),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_895),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_824),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_957),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1137),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_473),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1094),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1107),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1100),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_882),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_728),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1212),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_58),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_966),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_112),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_189),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1039),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_870),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_869),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_421),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_982),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_652),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_784),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_965),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_608),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1085),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1091),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_840),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_221),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1094),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1069),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1084),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1144),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1087),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1221),
.Y(n_1728)
);

BUFx2_ASAP7_75t_R g1729 ( 
.A(n_548),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1056),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_520),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_671),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1054),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1115),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1124),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_996),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_95),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1048),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_338),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1177),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_243),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1152),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_705),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_482),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1116),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_83),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_542),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_930),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1137),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1062),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_952),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_54),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1060),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_410),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1132),
.Y(n_1755)
);

BUFx10_ASAP7_75t_L g1756 ( 
.A(n_528),
.Y(n_1756)
);

CKINVDCx14_ASAP7_75t_R g1757 ( 
.A(n_1146),
.Y(n_1757)
);

CKINVDCx14_ASAP7_75t_R g1758 ( 
.A(n_787),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_850),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1179),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_20),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_715),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_456),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1129),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_958),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1184),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_963),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_817),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_343),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1109),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_689),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1143),
.Y(n_1772)
);

BUFx10_ASAP7_75t_L g1773 ( 
.A(n_1041),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_1070),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_434),
.Y(n_1775)
);

CKINVDCx16_ASAP7_75t_R g1776 ( 
.A(n_915),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1090),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_571),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_689),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1122),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1046),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1133),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_277),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1194),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_903),
.Y(n_1786)
);

CKINVDCx16_ASAP7_75t_R g1787 ( 
.A(n_1169),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_385),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_525),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1071),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_873),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1206),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_256),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_696),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_955),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_289),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_529),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1024),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_997),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1185),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_402),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1102),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_814),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_225),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_834),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1101),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_48),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_166),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1216),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_747),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_397),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_871),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_27),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_685),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1017),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_104),
.Y(n_1816)
);

CKINVDCx20_ASAP7_75t_R g1817 ( 
.A(n_766),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1103),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_624),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_792),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_950),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_53),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1224),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1079),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1081),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_735),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_986),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1095),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_52),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1134),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1121),
.Y(n_1831)
);

CKINVDCx20_ASAP7_75t_R g1832 ( 
.A(n_718),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1223),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1065),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_33),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_199),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_19),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_268),
.Y(n_1838)
);

BUFx10_ASAP7_75t_L g1839 ( 
.A(n_1128),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_175),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_342),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_344),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1103),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_522),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_566),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1139),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_949),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_820),
.Y(n_1848)
);

BUFx10_ASAP7_75t_L g1849 ( 
.A(n_997),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1022),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_58),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_962),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1160),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1050),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_799),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1322),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1322),
.Y(n_1857)
);

CKINVDCx20_ASAP7_75t_R g1858 ( 
.A(n_1339),
.Y(n_1858)
);

INVxp33_ASAP7_75t_SL g1859 ( 
.A(n_1677),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1322),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1322),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1440),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1440),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1440),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1440),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1440),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1296),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1477),
.Y(n_1868)
);

INVxp33_ASAP7_75t_SL g1869 ( 
.A(n_1298),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1650),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1477),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1477),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1477),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1477),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1230),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1265),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1266),
.Y(n_1877)
);

INVxp33_ASAP7_75t_SL g1878 ( 
.A(n_1319),
.Y(n_1878)
);

INVxp33_ASAP7_75t_L g1879 ( 
.A(n_1358),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1355),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1287),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1498),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1678),
.Y(n_1883)
);

NOR2xp67_ASAP7_75t_L g1884 ( 
.A(n_1498),
.B(n_0),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1341),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1343),
.Y(n_1886)
);

INVxp33_ASAP7_75t_SL g1887 ( 
.A(n_1436),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1379),
.Y(n_1888)
);

INVxp33_ASAP7_75t_SL g1889 ( 
.A(n_1473),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1277),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1277),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1277),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1680),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1757),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1257),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1416),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1310),
.Y(n_1897)
);

CKINVDCx20_ASAP7_75t_R g1898 ( 
.A(n_1758),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1454),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1227),
.Y(n_1900)
);

CKINVDCx16_ASAP7_75t_R g1901 ( 
.A(n_1453),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1469),
.Y(n_1902)
);

CKINVDCx20_ASAP7_75t_R g1903 ( 
.A(n_1569),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1448),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1679),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1689),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1775),
.Y(n_1907)
);

CKINVDCx20_ASAP7_75t_R g1908 ( 
.A(n_1776),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1560),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1584),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1611),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1623),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1708),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1709),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1722),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_1787),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1737),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1741),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1746),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1456),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1752),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1761),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1546),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1241),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_1228),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1796),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1804),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1461),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1813),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1840),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1448),
.Y(n_1931)
);

INVxp33_ASAP7_75t_L g1932 ( 
.A(n_1499),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1403),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1246),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1807),
.Y(n_1935)
);

INVxp67_ASAP7_75t_SL g1936 ( 
.A(n_1807),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1633),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1654),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_1253),
.Y(n_1939)
);

INVxp33_ASAP7_75t_SL g1940 ( 
.A(n_1772),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1660),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1846),
.Y(n_1942)
);

INVxp67_ASAP7_75t_SL g1943 ( 
.A(n_1807),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1783),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1620),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1837),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1465),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1478),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1504),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1627),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1706),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1850),
.Y(n_1952)
);

CKINVDCx20_ASAP7_75t_R g1953 ( 
.A(n_1316),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1261),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1326),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1237),
.Y(n_1956)
);

CKINVDCx20_ASAP7_75t_R g1957 ( 
.A(n_1338),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1280),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1280),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_1346),
.Y(n_1960)
);

INVxp33_ASAP7_75t_SL g1961 ( 
.A(n_1272),
.Y(n_1961)
);

INVxp67_ASAP7_75t_SL g1962 ( 
.A(n_1303),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1274),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1307),
.Y(n_1964)
);

INVxp33_ASAP7_75t_SL g1965 ( 
.A(n_1275),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1226),
.Y(n_1966)
);

CKINVDCx20_ASAP7_75t_R g1967 ( 
.A(n_1349),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1307),
.Y(n_1968)
);

CKINVDCx20_ASAP7_75t_R g1969 ( 
.A(n_1352),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1342),
.Y(n_1970)
);

BUFx2_ASAP7_75t_SL g1971 ( 
.A(n_1233),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1342),
.Y(n_1972)
);

CKINVDCx16_ASAP7_75t_R g1973 ( 
.A(n_1325),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1359),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1359),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1359),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1366),
.Y(n_1977)
);

INVxp67_ASAP7_75t_SL g1978 ( 
.A(n_1375),
.Y(n_1978)
);

INVxp33_ASAP7_75t_SL g1979 ( 
.A(n_1285),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1850),
.Y(n_1980)
);

CKINVDCx16_ASAP7_75t_R g1981 ( 
.A(n_1849),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1391),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1356),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1412),
.Y(n_1984)
);

INVxp33_ASAP7_75t_L g1985 ( 
.A(n_1562),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1289),
.Y(n_1986)
);

INVxp67_ASAP7_75t_SL g1987 ( 
.A(n_1441),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1460),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1488),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1488),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1357),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1488),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1489),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1362),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1489),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1509),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1317),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1321),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1509),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1850),
.Y(n_2000)
);

CKINVDCx20_ASAP7_75t_R g2001 ( 
.A(n_1364),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1851),
.Y(n_2002)
);

INVxp33_ASAP7_75t_L g2003 ( 
.A(n_1225),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1509),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1570),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1575),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1575),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1674),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1674),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1674),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1766),
.Y(n_2011)
);

INVxp33_ASAP7_75t_SL g2012 ( 
.A(n_1354),
.Y(n_2012)
);

INVxp67_ASAP7_75t_SL g2013 ( 
.A(n_1795),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1795),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1396),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1363),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1370),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1423),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1525),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_1925),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1952),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1962),
.Y(n_2022)
);

INVx4_ASAP7_75t_L g2023 ( 
.A(n_1924),
.Y(n_2023)
);

INVx4_ASAP7_75t_L g2024 ( 
.A(n_1934),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1897),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1968),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_1903),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1980),
.Y(n_2028)
);

OA21x2_ASAP7_75t_L g2029 ( 
.A1(n_1857),
.A2(n_1263),
.B(n_1235),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1882),
.B(n_1350),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1890),
.Y(n_2031)
);

CKINVDCx11_ASAP7_75t_R g2032 ( 
.A(n_1939),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1891),
.B(n_1458),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1867),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1976),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1985),
.A2(n_1382),
.B1(n_1385),
.B2(n_1374),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1961),
.B(n_1405),
.Y(n_2037)
);

OAI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1856),
.A2(n_1308),
.B(n_1284),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1978),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1988),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1989),
.Y(n_2041)
);

OA21x2_ASAP7_75t_L g2042 ( 
.A1(n_1860),
.A2(n_1340),
.B(n_1313),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1965),
.B(n_1411),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1990),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1890),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1892),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1892),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1892),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1870),
.B(n_1895),
.Y(n_2049)
);

OA21x2_ASAP7_75t_L g2050 ( 
.A1(n_1861),
.A2(n_1367),
.B(n_1360),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1977),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1904),
.B(n_1472),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2000),
.Y(n_2053)
);

BUFx12f_ASAP7_75t_L g2054 ( 
.A(n_1900),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1977),
.Y(n_2055)
);

INVx4_ASAP7_75t_L g2056 ( 
.A(n_1954),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1920),
.B(n_1923),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1945),
.B(n_1641),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1886),
.Y(n_2059)
);

BUFx12f_ASAP7_75t_L g2060 ( 
.A(n_1905),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1906),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1869),
.A2(n_1878),
.B1(n_1889),
.B2(n_1887),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1940),
.A2(n_1420),
.B1(n_1437),
.B2(n_1421),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1946),
.Y(n_2064)
);

INVxp67_ASAP7_75t_SL g2065 ( 
.A(n_1987),
.Y(n_2065)
);

INVx6_ASAP7_75t_L g2066 ( 
.A(n_2019),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2013),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1859),
.A2(n_1471),
.B1(n_1474),
.B2(n_1470),
.Y(n_2068)
);

OA21x2_ASAP7_75t_L g2069 ( 
.A1(n_1863),
.A2(n_1427),
.B(n_1419),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1931),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_1880),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1935),
.Y(n_2072)
);

INVx4_ASAP7_75t_L g2073 ( 
.A(n_1963),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1902),
.Y(n_2074)
);

OA21x2_ASAP7_75t_L g2075 ( 
.A1(n_1864),
.A2(n_1866),
.B(n_1865),
.Y(n_2075)
);

NOR2x1_ASAP7_75t_L g2076 ( 
.A(n_1868),
.B(n_1682),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1998),
.B(n_1700),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1919),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1936),
.B(n_1555),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1930),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1956),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1958),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1943),
.B(n_1710),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1986),
.Y(n_2084)
);

INVx4_ASAP7_75t_L g2085 ( 
.A(n_1997),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1959),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1971),
.B(n_2016),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2017),
.B(n_1566),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2015),
.B(n_1701),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1964),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1979),
.B(n_2012),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2018),
.B(n_1716),
.Y(n_2092)
);

OA21x2_ASAP7_75t_L g2093 ( 
.A1(n_1871),
.A2(n_1503),
.B(n_1483),
.Y(n_2093)
);

INVx6_ASAP7_75t_L g2094 ( 
.A(n_1973),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1970),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1972),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1907),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1974),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_1975),
.Y(n_2099)
);

NOR2x1_ASAP7_75t_L g2100 ( 
.A(n_1872),
.B(n_1723),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1982),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_1901),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1984),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_L g2104 ( 
.A(n_2002),
.B(n_1484),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1879),
.B(n_1735),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1992),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1993),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1995),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1996),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1999),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2004),
.Y(n_2111)
);

AND2x6_ASAP7_75t_L g2112 ( 
.A(n_1933),
.B(n_1259),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2005),
.Y(n_2113)
);

INVx5_ASAP7_75t_L g2114 ( 
.A(n_1981),
.Y(n_2114)
);

BUFx2_ASAP7_75t_L g2115 ( 
.A(n_1908),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2006),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2007),
.Y(n_2117)
);

AOI22x1_ASAP7_75t_SL g2118 ( 
.A1(n_1916),
.A2(n_1392),
.B1(n_1418),
.B2(n_1281),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_1858),
.A2(n_1521),
.B1(n_1522),
.B2(n_1520),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_1862),
.A2(n_1534),
.B(n_1513),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2008),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_2009),
.Y(n_2122)
);

OAI21x1_ASAP7_75t_L g2123 ( 
.A1(n_1873),
.A2(n_1594),
.B(n_1573),
.Y(n_2123)
);

OA21x2_ASAP7_75t_L g2124 ( 
.A1(n_1874),
.A2(n_2011),
.B(n_2010),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_1932),
.B(n_1550),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1937),
.B(n_1556),
.Y(n_2126)
);

BUFx12f_ASAP7_75t_L g2127 ( 
.A(n_1883),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_1893),
.A2(n_1579),
.B1(n_1591),
.B2(n_1588),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_1894),
.A2(n_1592),
.B1(n_1601),
.B2(n_1597),
.Y(n_2129)
);

AND2x6_ASAP7_75t_L g2130 ( 
.A(n_1938),
.B(n_1301),
.Y(n_2130)
);

INVx2_ASAP7_75t_SL g2131 ( 
.A(n_1928),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_SL g2132 ( 
.A(n_1898),
.B(n_1729),
.Y(n_2132)
);

INVxp67_ASAP7_75t_L g2133 ( 
.A(n_1942),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2014),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1966),
.B(n_1602),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1875),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1941),
.B(n_1606),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1876),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1877),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2003),
.B(n_1823),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1944),
.B(n_1610),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1881),
.Y(n_2142)
);

OAI21x1_ASAP7_75t_L g2143 ( 
.A1(n_1885),
.A2(n_1621),
.B(n_1619),
.Y(n_2143)
);

NOR2x1_ASAP7_75t_L g2144 ( 
.A(n_1884),
.B(n_1847),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1888),
.B(n_1618),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1896),
.Y(n_2146)
);

OA21x2_ASAP7_75t_L g2147 ( 
.A1(n_1899),
.A2(n_1652),
.B(n_1647),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_2032),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_2020),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2136),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2140),
.B(n_2105),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2037),
.B(n_2043),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_2051),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_2127),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2021),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_2034),
.Y(n_2156)
);

CKINVDCx20_ASAP7_75t_R g2157 ( 
.A(n_2027),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_2054),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2026),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_2060),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2028),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_2023),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_2024),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_2056),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_2073),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2040),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2065),
.B(n_1909),
.Y(n_2167)
);

BUFx3_ASAP7_75t_L g2168 ( 
.A(n_2066),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_2085),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2041),
.Y(n_2170)
);

CKINVDCx20_ASAP7_75t_R g2171 ( 
.A(n_2061),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2044),
.Y(n_2172)
);

BUFx2_ASAP7_75t_L g2173 ( 
.A(n_2102),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_2055),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_2031),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_2045),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_2097),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2139),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_2115),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_2114),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_2091),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2142),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_2094),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_2071),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_R g2185 ( 
.A(n_2104),
.B(n_1953),
.Y(n_2185)
);

NAND2xp33_ASAP7_75t_R g2186 ( 
.A(n_2049),
.B(n_1637),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2053),
.Y(n_2187)
);

AND3x2_ASAP7_75t_L g2188 ( 
.A(n_2132),
.B(n_1430),
.C(n_1347),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_2087),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_2083),
.Y(n_2190)
);

OA21x2_ASAP7_75t_L g2191 ( 
.A1(n_2038),
.A2(n_1911),
.B(n_1910),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2088),
.B(n_2022),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2035),
.B(n_1912),
.Y(n_2193)
);

INVxp67_ASAP7_75t_L g2194 ( 
.A(n_2125),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_2128),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_R g2196 ( 
.A(n_2070),
.B(n_1955),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_2062),
.Y(n_2197)
);

INVxp67_ASAP7_75t_SL g2198 ( 
.A(n_2075),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2059),
.Y(n_2199)
);

CKINVDCx20_ASAP7_75t_R g2200 ( 
.A(n_2119),
.Y(n_2200)
);

AND2x6_ASAP7_75t_L g2201 ( 
.A(n_2144),
.B(n_1229),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_2046),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2074),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_R g2204 ( 
.A(n_2072),
.B(n_1957),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2078),
.Y(n_2205)
);

BUFx10_ASAP7_75t_L g2206 ( 
.A(n_2057),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2080),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_R g2208 ( 
.A(n_2039),
.B(n_1960),
.Y(n_2208)
);

BUFx3_ASAP7_75t_L g2209 ( 
.A(n_2029),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_2036),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2143),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_2118),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_2129),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2138),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_2063),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_2077),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_2135),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_2068),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_2131),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_2067),
.Y(n_2220)
);

CKINVDCx20_ASAP7_75t_R g2221 ( 
.A(n_2133),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2030),
.B(n_1913),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_R g2223 ( 
.A(n_2033),
.B(n_1967),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2112),
.Y(n_2224)
);

CKINVDCx20_ASAP7_75t_R g2225 ( 
.A(n_2126),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2146),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_R g2227 ( 
.A(n_2052),
.B(n_1969),
.Y(n_2227)
);

CKINVDCx20_ASAP7_75t_R g2228 ( 
.A(n_2137),
.Y(n_2228)
);

INVxp67_ASAP7_75t_SL g2229 ( 
.A(n_2124),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2058),
.Y(n_2230)
);

INVxp67_ASAP7_75t_L g2231 ( 
.A(n_2145),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2042),
.B(n_1914),
.Y(n_2232)
);

CKINVDCx20_ASAP7_75t_R g2233 ( 
.A(n_2141),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2064),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_2050),
.Y(n_2235)
);

AOI21x1_ASAP7_75t_L g2236 ( 
.A1(n_2120),
.A2(n_1917),
.B(n_1915),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2069),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2086),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_2130),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_2130),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2093),
.B(n_1918),
.Y(n_2241)
);

CKINVDCx20_ASAP7_75t_R g2242 ( 
.A(n_2079),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_2047),
.Y(n_2243)
);

BUFx2_ASAP7_75t_L g2244 ( 
.A(n_2076),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_2081),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_2082),
.Y(n_2246)
);

HB1xp67_ASAP7_75t_L g2247 ( 
.A(n_2048),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_2107),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_R g2249 ( 
.A(n_2089),
.B(n_1983),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_2108),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_2110),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_2122),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2092),
.B(n_1921),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2100),
.B(n_1922),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2123),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_2090),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_R g2257 ( 
.A(n_2099),
.B(n_1991),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_2095),
.Y(n_2258)
);

CKINVDCx20_ASAP7_75t_R g2259 ( 
.A(n_2147),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_R g2260 ( 
.A(n_2103),
.B(n_1994),
.Y(n_2260)
);

BUFx2_ASAP7_75t_L g2261 ( 
.A(n_2096),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_R g2262 ( 
.A(n_2098),
.B(n_2001),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2101),
.Y(n_2263)
);

BUFx6f_ASAP7_75t_L g2264 ( 
.A(n_2111),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_2113),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_2117),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2106),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_R g2268 ( 
.A(n_2109),
.B(n_1373),
.Y(n_2268)
);

BUFx10_ASAP7_75t_L g2269 ( 
.A(n_2116),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_2121),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2134),
.A2(n_1531),
.B1(n_1315),
.B2(n_1327),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2084),
.Y(n_2272)
);

BUFx10_ASAP7_75t_L g2273 ( 
.A(n_2094),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_2025),
.Y(n_2274)
);

CKINVDCx20_ASAP7_75t_R g2275 ( 
.A(n_2020),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2136),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2025),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2140),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2155),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2159),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_2231),
.B(n_1452),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2192),
.B(n_1926),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2191),
.Y(n_2283)
);

INVxp67_ASAP7_75t_SL g2284 ( 
.A(n_2209),
.Y(n_2284)
);

INVx5_ASAP7_75t_L g2285 ( 
.A(n_2273),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2168),
.B(n_1927),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2236),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2152),
.B(n_2217),
.Y(n_2288)
);

BUFx3_ASAP7_75t_L g2289 ( 
.A(n_2274),
.Y(n_2289)
);

INVx5_ASAP7_75t_L g2290 ( 
.A(n_2206),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2278),
.B(n_1929),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2198),
.B(n_1231),
.Y(n_2292)
);

AOI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_2232),
.A2(n_1667),
.B1(n_1688),
.B2(n_1655),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2161),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_2241),
.A2(n_2259),
.B1(n_2235),
.B2(n_2237),
.Y(n_2295)
);

BUFx3_ASAP7_75t_L g2296 ( 
.A(n_2246),
.Y(n_2296)
);

INVxp67_ASAP7_75t_L g2297 ( 
.A(n_2186),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2173),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2181),
.B(n_1468),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2220),
.B(n_2219),
.Y(n_2300)
);

CKINVDCx20_ASAP7_75t_R g2301 ( 
.A(n_2275),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_2242),
.B(n_1479),
.Y(n_2302)
);

BUFx10_ASAP7_75t_L g2303 ( 
.A(n_2158),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2150),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2175),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_2162),
.B(n_1234),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2229),
.B(n_1236),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_2269),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2163),
.B(n_1238),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2277),
.B(n_1947),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2166),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2170),
.Y(n_2312)
);

NAND2xp33_ASAP7_75t_SL g2313 ( 
.A(n_2224),
.B(n_1836),
.Y(n_2313)
);

NAND2x1p5_ASAP7_75t_L g2314 ( 
.A(n_2190),
.B(n_1948),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_2272),
.Y(n_2315)
);

BUFx4f_ASAP7_75t_L g2316 ( 
.A(n_2201),
.Y(n_2316)
);

INVx3_ASAP7_75t_L g2317 ( 
.A(n_2176),
.Y(n_2317)
);

INVx4_ASAP7_75t_L g2318 ( 
.A(n_2248),
.Y(n_2318)
);

BUFx4f_ASAP7_75t_L g2319 ( 
.A(n_2201),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2172),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2211),
.A2(n_2255),
.B1(n_2276),
.B2(n_2167),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_2202),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2202),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2187),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2267),
.Y(n_2325)
);

AND2x6_ASAP7_75t_L g2326 ( 
.A(n_2254),
.B(n_1232),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_2202),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_2164),
.B(n_1239),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2210),
.B(n_1528),
.Y(n_2329)
);

INVx5_ASAP7_75t_L g2330 ( 
.A(n_2243),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2214),
.Y(n_2331)
);

BUFx8_ASAP7_75t_SL g2332 ( 
.A(n_2148),
.Y(n_2332)
);

INVx5_ASAP7_75t_L g2333 ( 
.A(n_2243),
.Y(n_2333)
);

INVx2_ASAP7_75t_SL g2334 ( 
.A(n_2256),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2250),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2253),
.B(n_1505),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2165),
.B(n_1240),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_SL g2338 ( 
.A(n_2169),
.B(n_1242),
.Y(n_2338)
);

AND2x6_ASAP7_75t_L g2339 ( 
.A(n_2207),
.B(n_1251),
.Y(n_2339)
);

NAND2x1p5_ASAP7_75t_L g2340 ( 
.A(n_2178),
.B(n_1949),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2226),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2234),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2218),
.B(n_1544),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2222),
.B(n_1243),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2268),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2238),
.Y(n_2346)
);

BUFx6f_ASAP7_75t_L g2347 ( 
.A(n_2153),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2263),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2261),
.B(n_1505),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2215),
.B(n_1574),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2251),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2252),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2258),
.B(n_1244),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2199),
.B(n_2203),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2205),
.B(n_1950),
.Y(n_2355)
);

AND2x6_ASAP7_75t_L g2356 ( 
.A(n_2271),
.B(n_1255),
.Y(n_2356)
);

OR2x2_ASAP7_75t_SL g2357 ( 
.A(n_2213),
.B(n_1728),
.Y(n_2357)
);

NOR2xp33_ASAP7_75t_L g2358 ( 
.A(n_2265),
.B(n_1663),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2270),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_2182),
.B(n_1951),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2193),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2266),
.Y(n_2362)
);

CKINVDCx20_ASAP7_75t_R g2363 ( 
.A(n_2149),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2264),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2247),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2225),
.B(n_1687),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2239),
.B(n_2240),
.Y(n_2367)
);

INVx1_ASAP7_75t_SL g2368 ( 
.A(n_2260),
.Y(n_2368)
);

INVxp67_ASAP7_75t_SL g2369 ( 
.A(n_2244),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2230),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2184),
.B(n_1519),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2223),
.B(n_1245),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2228),
.B(n_1699),
.Y(n_2373)
);

BUFx4f_ASAP7_75t_L g2374 ( 
.A(n_2160),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2233),
.B(n_1247),
.Y(n_2375)
);

INVx4_ASAP7_75t_L g2376 ( 
.A(n_2183),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2227),
.B(n_1248),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2249),
.B(n_1249),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2188),
.Y(n_2379)
);

AND2x6_ASAP7_75t_L g2380 ( 
.A(n_2185),
.B(n_1258),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_2195),
.B(n_1736),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_2196),
.B(n_1250),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2204),
.B(n_1252),
.Y(n_2383)
);

INVx1_ASAP7_75t_SL g2384 ( 
.A(n_2221),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2208),
.B(n_1254),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2262),
.B(n_1256),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2177),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2179),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2157),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2180),
.B(n_1260),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2197),
.B(n_1742),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2200),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2171),
.B(n_1267),
.Y(n_2393)
);

INVx4_ASAP7_75t_L g2394 ( 
.A(n_2156),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2154),
.B(n_1262),
.Y(n_2395)
);

OAI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2212),
.A2(n_1475),
.B1(n_1646),
.B2(n_1443),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2191),
.Y(n_2397)
);

INVx4_ASAP7_75t_SL g2398 ( 
.A(n_2201),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2191),
.Y(n_2399)
);

BUFx4f_ASAP7_75t_L g2400 ( 
.A(n_2201),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2192),
.B(n_1264),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2189),
.B(n_1268),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2191),
.Y(n_2403)
);

AND2x6_ASAP7_75t_L g2404 ( 
.A(n_2151),
.B(n_1270),
.Y(n_2404)
);

OAI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2259),
.A2(n_1712),
.B1(n_1802),
.B2(n_1691),
.Y(n_2405)
);

AND2x6_ASAP7_75t_L g2406 ( 
.A(n_2151),
.B(n_1273),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2168),
.B(n_1276),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2151),
.B(n_1600),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2191),
.Y(n_2409)
);

AND2x6_ASAP7_75t_L g2410 ( 
.A(n_2151),
.B(n_1279),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2202),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_2194),
.B(n_1791),
.Y(n_2412)
);

INVxp67_ASAP7_75t_L g2413 ( 
.A(n_2186),
.Y(n_2413)
);

AND2x6_ASAP7_75t_L g2414 ( 
.A(n_2151),
.B(n_1288),
.Y(n_2414)
);

INVx4_ASAP7_75t_L g2415 ( 
.A(n_2245),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2191),
.Y(n_2416)
);

CKINVDCx16_ASAP7_75t_R g2417 ( 
.A(n_2275),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2192),
.B(n_1269),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_2202),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2189),
.B(n_1271),
.Y(n_2420)
);

INVxp33_ASAP7_75t_L g2421 ( 
.A(n_2257),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2151),
.B(n_1600),
.Y(n_2422)
);

INVx5_ASAP7_75t_L g2423 ( 
.A(n_2273),
.Y(n_2423)
);

INVxp33_ASAP7_75t_L g2424 ( 
.A(n_2257),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2191),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_2168),
.B(n_1290),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2151),
.B(n_1625),
.Y(n_2427)
);

INVx4_ASAP7_75t_L g2428 ( 
.A(n_2245),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2194),
.B(n_1794),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2151),
.B(n_1625),
.Y(n_2430)
);

BUFx4f_ASAP7_75t_L g2431 ( 
.A(n_2201),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2278),
.B(n_1803),
.Y(n_2432)
);

INVx1_ASAP7_75t_SL g2433 ( 
.A(n_2219),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2202),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2155),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2192),
.B(n_1278),
.Y(n_2436)
);

BUFx2_ASAP7_75t_L g2437 ( 
.A(n_2216),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2155),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2191),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2232),
.A2(n_1297),
.B1(n_1300),
.B2(n_1295),
.Y(n_2440)
);

BUFx6f_ASAP7_75t_L g2441 ( 
.A(n_2202),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2194),
.B(n_1826),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2191),
.Y(n_2443)
);

INVx3_ASAP7_75t_L g2444 ( 
.A(n_2174),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2151),
.B(n_1632),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2151),
.B(n_1632),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2151),
.B(n_1662),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2279),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2288),
.B(n_1480),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2322),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2334),
.B(n_1486),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2284),
.A2(n_1304),
.B(n_1302),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2280),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2294),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2401),
.B(n_1282),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2311),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2418),
.B(n_1283),
.Y(n_2457)
);

INVx5_ASAP7_75t_L g2458 ( 
.A(n_2351),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2299),
.B(n_1545),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2436),
.B(n_1286),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2381),
.B(n_1547),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2312),
.Y(n_2462)
);

NAND3xp33_ASAP7_75t_L g2463 ( 
.A(n_2329),
.B(n_1292),
.C(n_1291),
.Y(n_2463)
);

A2O1A1Ixp33_ASAP7_75t_L g2464 ( 
.A1(n_2281),
.A2(n_1306),
.B(n_1311),
.C(n_1305),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_SL g2465 ( 
.A(n_2303),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2320),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2343),
.B(n_1568),
.Y(n_2467)
);

INVx2_ASAP7_75t_SL g2468 ( 
.A(n_2298),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2412),
.B(n_1662),
.Y(n_2469)
);

NOR2xp33_ASAP7_75t_L g2470 ( 
.A(n_2391),
.B(n_2350),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2324),
.Y(n_2471)
);

NAND2x1_ASAP7_75t_L g2472 ( 
.A(n_2283),
.B(n_1312),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2282),
.B(n_2429),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2442),
.B(n_1293),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2297),
.B(n_1578),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_L g2476 ( 
.A(n_2413),
.B(n_1590),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2295),
.B(n_1294),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2321),
.A2(n_1616),
.B1(n_1629),
.B2(n_1603),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2435),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2300),
.B(n_1635),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_2322),
.Y(n_2481)
);

INVx8_ASAP7_75t_L g2482 ( 
.A(n_2423),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2344),
.B(n_1299),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2438),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2323),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2292),
.B(n_1309),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2358),
.B(n_1756),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_2327),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2325),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2307),
.B(n_1314),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_2362),
.B(n_1744),
.Y(n_2491)
);

AOI22xp33_ASAP7_75t_L g2492 ( 
.A1(n_2440),
.A2(n_1788),
.B1(n_1799),
.B2(n_1774),
.Y(n_2492)
);

O2A1O1Ixp33_ASAP7_75t_L g2493 ( 
.A1(n_2405),
.A2(n_1323),
.B(n_1328),
.C(n_1320),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2331),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2408),
.B(n_1318),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_2327),
.Y(n_2496)
);

A2O1A1Ixp33_ASAP7_75t_L g2497 ( 
.A1(n_2422),
.A2(n_1332),
.B(n_1335),
.C(n_1329),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2393),
.Y(n_2498)
);

O2A1O1Ixp5_ASAP7_75t_L g2499 ( 
.A1(n_2287),
.A2(n_1348),
.B(n_1351),
.C(n_1345),
.Y(n_2499)
);

AOI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2404),
.A2(n_1832),
.B1(n_1834),
.B2(n_1817),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2427),
.B(n_2430),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2445),
.B(n_1324),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2342),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2446),
.B(n_2447),
.Y(n_2504)
);

AOI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_2397),
.A2(n_1365),
.B(n_1361),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2336),
.B(n_2291),
.Y(n_2506)
);

NOR3x1_ASAP7_75t_L g2507 ( 
.A(n_2396),
.B(n_1377),
.C(n_1376),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2330),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2349),
.B(n_1773),
.Y(n_2509)
);

BUFx5_ASAP7_75t_L g2510 ( 
.A(n_2399),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2421),
.B(n_1330),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2406),
.A2(n_1393),
.B1(n_1395),
.B2(n_1387),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2424),
.B(n_1331),
.Y(n_2513)
);

AOI22xp33_ASAP7_75t_L g2514 ( 
.A1(n_2410),
.A2(n_1401),
.B1(n_1413),
.B2(n_1399),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2433),
.B(n_1333),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2410),
.A2(n_1417),
.B1(n_1424),
.B2(n_1415),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2302),
.B(n_2368),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2366),
.B(n_1334),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2346),
.B(n_1336),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2373),
.B(n_1337),
.Y(n_2520)
);

INVx2_ASAP7_75t_SL g2521 ( 
.A(n_2330),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_SL g2522 ( 
.A(n_2315),
.B(n_1839),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2375),
.B(n_1784),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2359),
.B(n_1344),
.Y(n_2524)
);

INVxp67_ASAP7_75t_L g2525 ( 
.A(n_2432),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2316),
.B(n_2319),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2400),
.B(n_1353),
.Y(n_2527)
);

NAND2xp33_ASAP7_75t_L g2528 ( 
.A(n_2414),
.B(n_1793),
.Y(n_2528)
);

BUFx6f_ASAP7_75t_L g2529 ( 
.A(n_2411),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2341),
.Y(n_2530)
);

OAI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_2348),
.A2(n_1816),
.B1(n_1822),
.B2(n_1808),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2355),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2403),
.A2(n_1429),
.B(n_1426),
.Y(n_2533)
);

BUFx3_ASAP7_75t_L g2534 ( 
.A(n_2296),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2360),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2409),
.B(n_1368),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2416),
.B(n_1369),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2364),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2425),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2371),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2431),
.B(n_1371),
.Y(n_2541)
);

NOR2x1p5_ASAP7_75t_L g2542 ( 
.A(n_2335),
.B(n_1829),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2439),
.B(n_1372),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2443),
.B(n_2293),
.Y(n_2544)
);

AOI22xp33_ASAP7_75t_L g2545 ( 
.A1(n_2326),
.A2(n_1433),
.B1(n_1435),
.B2(n_1432),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2345),
.B(n_2308),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2310),
.Y(n_2547)
);

AOI22xp33_ASAP7_75t_L g2548 ( 
.A1(n_2326),
.A2(n_1442),
.B1(n_1446),
.B2(n_1439),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2377),
.B(n_1378),
.Y(n_2549)
);

O2A1O1Ixp5_ASAP7_75t_L g2550 ( 
.A1(n_2402),
.A2(n_1449),
.B(n_1451),
.C(n_1447),
.Y(n_2550)
);

INVx2_ASAP7_75t_SL g2551 ( 
.A(n_2333),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2354),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2369),
.B(n_1835),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2318),
.B(n_1380),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2420),
.B(n_1381),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2378),
.B(n_1383),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2340),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2415),
.B(n_1384),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2419),
.Y(n_2559)
);

NAND2xp33_ASAP7_75t_L g2560 ( 
.A(n_2380),
.B(n_1838),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2380),
.B(n_1386),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2365),
.Y(n_2562)
);

O2A1O1Ixp5_ASAP7_75t_L g2563 ( 
.A1(n_2372),
.A2(n_1462),
.B(n_1463),
.C(n_1455),
.Y(n_2563)
);

INVx4_ASAP7_75t_L g2564 ( 
.A(n_2352),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2419),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2379),
.B(n_1388),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_2428),
.B(n_1389),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2306),
.B(n_2309),
.Y(n_2568)
);

A2O1A1Ixp33_ASAP7_75t_L g2569 ( 
.A1(n_2313),
.A2(n_2353),
.B(n_2337),
.C(n_2338),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2328),
.B(n_1390),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2434),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2437),
.B(n_1394),
.Y(n_2572)
);

OAI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2387),
.A2(n_1398),
.B1(n_1400),
.B2(n_1397),
.Y(n_2573)
);

NAND3xp33_ASAP7_75t_L g2574 ( 
.A(n_2388),
.B(n_1404),
.C(n_1402),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2367),
.A2(n_1407),
.B1(n_1408),
.B2(n_1406),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2441),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2441),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2314),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_2384),
.B(n_1409),
.Y(n_2579)
);

NOR3xp33_ASAP7_75t_L g2580 ( 
.A(n_2382),
.B(n_1414),
.C(n_1410),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2357),
.Y(n_2581)
);

INVx2_ASAP7_75t_SL g2582 ( 
.A(n_2286),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2290),
.B(n_1422),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2395),
.B(n_1425),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2407),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2290),
.B(n_1428),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2426),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2383),
.B(n_1431),
.Y(n_2588)
);

BUFx5_ASAP7_75t_L g2589 ( 
.A(n_2289),
.Y(n_2589)
);

OR2x6_ASAP7_75t_L g2590 ( 
.A(n_2376),
.B(n_1464),
.Y(n_2590)
);

NOR2xp67_ASAP7_75t_L g2591 ( 
.A(n_2394),
.B(n_1434),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2385),
.B(n_1438),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2386),
.B(n_1444),
.Y(n_2593)
);

AND2x2_ASAP7_75t_SL g2594 ( 
.A(n_2417),
.B(n_1466),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2389),
.B(n_1445),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2305),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2392),
.B(n_1450),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2398),
.B(n_1457),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2317),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2356),
.B(n_1459),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2347),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2444),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2370),
.B(n_1467),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2390),
.A2(n_1492),
.B(n_1481),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2374),
.B(n_1476),
.Y(n_2605)
);

INVx4_ASAP7_75t_L g2606 ( 
.A(n_2332),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_L g2607 ( 
.A(n_2363),
.B(n_1482),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2339),
.B(n_1485),
.Y(n_2608)
);

OAI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2301),
.A2(n_1490),
.B1(n_1491),
.B2(n_1487),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2304),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2285),
.B(n_1493),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_L g2612 ( 
.A(n_2299),
.B(n_1494),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2361),
.B(n_1495),
.Y(n_2613)
);

NAND3xp33_ASAP7_75t_L g2614 ( 
.A(n_2299),
.B(n_1497),
.C(n_1496),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2361),
.B(n_1500),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2299),
.B(n_1501),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2304),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2361),
.B(n_1502),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2304),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2412),
.B(n_1507),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2361),
.B(n_1511),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2299),
.B(n_1512),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2304),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_L g2624 ( 
.A1(n_2361),
.A2(n_1508),
.B1(n_1510),
.B2(n_1506),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_L g2625 ( 
.A(n_2299),
.B(n_1523),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2412),
.B(n_1524),
.Y(n_2626)
);

OAI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2295),
.A2(n_1529),
.B1(n_1530),
.B2(n_1526),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2412),
.B(n_1532),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2288),
.B(n_1533),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2304),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2304),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2361),
.A2(n_1515),
.B1(n_1516),
.B2(n_1514),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2288),
.B(n_1535),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2288),
.A2(n_1518),
.B(n_1527),
.C(n_1517),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2299),
.B(n_1536),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2279),
.Y(n_2636)
);

BUFx6f_ASAP7_75t_L g2637 ( 
.A(n_2322),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2361),
.B(n_1539),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2470),
.A2(n_1541),
.B1(n_1542),
.B2(n_1540),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2473),
.B(n_1543),
.Y(n_2640)
);

OAI21xp33_ASAP7_75t_L g2641 ( 
.A1(n_2467),
.A2(n_2459),
.B(n_2461),
.Y(n_2641)
);

AOI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2544),
.A2(n_1538),
.B(n_1537),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2564),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2568),
.A2(n_2539),
.B(n_2504),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2612),
.B(n_1548),
.Y(n_2645)
);

A2O1A1Ixp33_ASAP7_75t_L g2646 ( 
.A1(n_2616),
.A2(n_1557),
.B(n_1567),
.C(n_1553),
.Y(n_2646)
);

AOI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2501),
.A2(n_1577),
.B(n_1572),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2530),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2622),
.B(n_1549),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2448),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2453),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_L g2652 ( 
.A(n_2517),
.B(n_1551),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2625),
.B(n_1552),
.Y(n_2653)
);

OR2x2_ASAP7_75t_L g2654 ( 
.A(n_2506),
.B(n_1554),
.Y(n_2654)
);

AOI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2486),
.A2(n_1582),
.B(n_1581),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2635),
.B(n_1558),
.Y(n_2656)
);

OAI21xp33_ASAP7_75t_L g2657 ( 
.A1(n_2518),
.A2(n_1561),
.B(n_1559),
.Y(n_2657)
);

HB1xp67_ASAP7_75t_L g2658 ( 
.A(n_2468),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2454),
.Y(n_2659)
);

AOI21xp5_ASAP7_75t_L g2660 ( 
.A1(n_2490),
.A2(n_1589),
.B(n_1587),
.Y(n_2660)
);

O2A1O1Ixp33_ASAP7_75t_L g2661 ( 
.A1(n_2474),
.A2(n_1598),
.B(n_1599),
.C(n_1595),
.Y(n_2661)
);

OAI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2536),
.A2(n_2543),
.B(n_2537),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2456),
.Y(n_2663)
);

OAI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2505),
.A2(n_1614),
.B(n_1613),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2620),
.B(n_1563),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2569),
.A2(n_1624),
.B(n_1622),
.Y(n_2666)
);

O2A1O1Ixp33_ASAP7_75t_L g2667 ( 
.A1(n_2497),
.A2(n_1630),
.B(n_1634),
.C(n_1626),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2462),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2626),
.B(n_1564),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2628),
.B(n_1565),
.Y(n_2670)
);

OAI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2533),
.A2(n_1642),
.B(n_1640),
.Y(n_2671)
);

OAI21xp33_ASAP7_75t_L g2672 ( 
.A1(n_2520),
.A2(n_1576),
.B(n_1571),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2455),
.B(n_1580),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2457),
.A2(n_1651),
.B(n_1644),
.Y(n_2674)
);

NOR3xp33_ASAP7_75t_L g2675 ( 
.A(n_2449),
.B(n_1585),
.C(n_1583),
.Y(n_2675)
);

OAI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2499),
.A2(n_1659),
.B(n_1653),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2460),
.B(n_1586),
.Y(n_2677)
);

AOI22xp33_ASAP7_75t_L g2678 ( 
.A1(n_2581),
.A2(n_1664),
.B1(n_1666),
.B2(n_1661),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2534),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2458),
.B(n_1593),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2465),
.Y(n_2681)
);

AOI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_2483),
.A2(n_1681),
.B(n_1675),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2466),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2584),
.B(n_1596),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2556),
.A2(n_1686),
.B(n_1685),
.Y(n_2685)
);

O2A1O1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2629),
.A2(n_2633),
.B(n_2464),
.C(n_2493),
.Y(n_2686)
);

INVx4_ASAP7_75t_L g2687 ( 
.A(n_2482),
.Y(n_2687)
);

CKINVDCx10_ASAP7_75t_R g2688 ( 
.A(n_2590),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2469),
.A2(n_1696),
.B1(n_1697),
.B2(n_1692),
.Y(n_2689)
);

OAI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2477),
.A2(n_1703),
.B(n_1698),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2489),
.B(n_1604),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2450),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2610),
.B(n_1605),
.Y(n_2693)
);

O2A1O1Ixp33_ASAP7_75t_L g2694 ( 
.A1(n_2634),
.A2(n_1713),
.B(n_1714),
.C(n_1711),
.Y(n_2694)
);

OAI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2617),
.A2(n_1608),
.B1(n_1609),
.B2(n_1607),
.Y(n_2695)
);

INVx3_ASAP7_75t_L g2696 ( 
.A(n_2450),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2619),
.B(n_1612),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2623),
.B(n_1615),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2475),
.B(n_1617),
.Y(n_2699)
);

NAND2x1_ASAP7_75t_L g2700 ( 
.A(n_2471),
.B(n_1717),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2630),
.Y(n_2701)
);

A2O1A1Ixp33_ASAP7_75t_L g2702 ( 
.A1(n_2555),
.A2(n_1719),
.B(n_1725),
.C(n_1718),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2613),
.A2(n_1734),
.B(n_1733),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2631),
.B(n_1628),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2615),
.A2(n_1743),
.B(n_1738),
.Y(n_2705)
);

OAI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2472),
.A2(n_2621),
.B(n_2618),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2589),
.B(n_2525),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2487),
.B(n_1631),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2638),
.B(n_1636),
.Y(n_2709)
);

BUFx12f_ASAP7_75t_L g2710 ( 
.A(n_2606),
.Y(n_2710)
);

O2A1O1Ixp33_ASAP7_75t_L g2711 ( 
.A1(n_2495),
.A2(n_1748),
.B(n_1749),
.C(n_1747),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2494),
.B(n_1638),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2476),
.B(n_1639),
.Y(n_2713)
);

INVx3_ASAP7_75t_L g2714 ( 
.A(n_2481),
.Y(n_2714)
);

BUFx4f_ASAP7_75t_L g2715 ( 
.A(n_2488),
.Y(n_2715)
);

OAI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2540),
.A2(n_1645),
.B1(n_1648),
.B2(n_1643),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2502),
.B(n_1649),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2479),
.Y(n_2718)
);

NAND2xp33_ASAP7_75t_SL g2719 ( 
.A(n_2526),
.B(n_1656),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2484),
.A2(n_1760),
.B(n_1753),
.Y(n_2720)
);

AOI21x1_ASAP7_75t_L g2721 ( 
.A1(n_2527),
.A2(n_1765),
.B(n_1764),
.Y(n_2721)
);

INVx5_ASAP7_75t_L g2722 ( 
.A(n_2529),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2593),
.B(n_1657),
.Y(n_2723)
);

AOI21xp5_ASAP7_75t_L g2724 ( 
.A1(n_2503),
.A2(n_1771),
.B(n_1769),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2553),
.B(n_1658),
.Y(n_2725)
);

OAI21xp33_ASAP7_75t_L g2726 ( 
.A1(n_2492),
.A2(n_1668),
.B(n_1665),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2589),
.B(n_1669),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2511),
.B(n_1670),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2513),
.B(n_1671),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2523),
.B(n_1672),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2636),
.A2(n_1778),
.B1(n_1779),
.B2(n_1777),
.Y(n_2731)
);

NAND2x1_ASAP7_75t_L g2732 ( 
.A(n_2485),
.B(n_1780),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2624),
.B(n_1673),
.Y(n_2733)
);

AOI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2524),
.A2(n_2519),
.B(n_2549),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2632),
.B(n_1676),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2541),
.A2(n_1801),
.B(n_1800),
.Y(n_2736)
);

O2A1O1Ixp5_ASAP7_75t_L g2737 ( 
.A1(n_2588),
.A2(n_1806),
.B(n_1809),
.C(n_1805),
.Y(n_2737)
);

INVx2_ASAP7_75t_SL g2738 ( 
.A(n_2498),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2582),
.B(n_1811),
.Y(n_2739)
);

BUFx12f_ASAP7_75t_L g2740 ( 
.A(n_2529),
.Y(n_2740)
);

NAND3xp33_ASAP7_75t_L g2741 ( 
.A(n_2579),
.B(n_1684),
.C(n_1683),
.Y(n_2741)
);

AOI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2592),
.A2(n_1819),
.B(n_1815),
.Y(n_2742)
);

BUFx2_ASAP7_75t_SL g2743 ( 
.A(n_2508),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2562),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2597),
.B(n_1690),
.Y(n_2745)
);

OAI21xp33_ASAP7_75t_L g2746 ( 
.A1(n_2478),
.A2(n_1694),
.B(n_1693),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2452),
.B(n_1695),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2509),
.B(n_1702),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2538),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2480),
.B(n_1704),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2637),
.Y(n_2751)
);

AOI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2570),
.A2(n_1844),
.B(n_1843),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2559),
.Y(n_2753)
);

AOI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2578),
.A2(n_1848),
.B(n_1845),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2572),
.B(n_1705),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2491),
.B(n_2451),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2565),
.Y(n_2757)
);

BUFx6f_ASAP7_75t_L g2758 ( 
.A(n_2521),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2463),
.B(n_1707),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2510),
.B(n_1715),
.Y(n_2760)
);

OAI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2614),
.A2(n_1721),
.B(n_1720),
.Y(n_2761)
);

OAI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2566),
.A2(n_1726),
.B(n_1724),
.Y(n_2762)
);

A2O1A1Ixp33_ASAP7_75t_L g2763 ( 
.A1(n_2603),
.A2(n_1730),
.B(n_1731),
.C(n_1727),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2522),
.B(n_1732),
.Y(n_2764)
);

INVxp67_ASAP7_75t_L g2765 ( 
.A(n_2595),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2607),
.B(n_1739),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2594),
.B(n_1740),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2571),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2580),
.A2(n_1750),
.B1(n_1751),
.B2(n_1745),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2547),
.A2(n_1755),
.B(n_1754),
.Y(n_2770)
);

OAI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2550),
.A2(n_2563),
.B(n_2627),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2500),
.B(n_1759),
.Y(n_2772)
);

NOR3xp33_ASAP7_75t_L g2773 ( 
.A(n_2609),
.B(n_1763),
.C(n_1762),
.Y(n_2773)
);

OAI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2574),
.A2(n_1768),
.B(n_1767),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2512),
.B(n_1770),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2514),
.B(n_2516),
.Y(n_2776)
);

BUFx2_ASAP7_75t_L g2777 ( 
.A(n_2496),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2545),
.B(n_1781),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2548),
.B(n_1782),
.Y(n_2779)
);

OAI21x1_ASAP7_75t_L g2780 ( 
.A1(n_2557),
.A2(n_324),
.B(n_323),
.Y(n_2780)
);

OAI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2600),
.A2(n_1786),
.B(n_1785),
.Y(n_2781)
);

INVx11_ASAP7_75t_L g2782 ( 
.A(n_2551),
.Y(n_2782)
);

O2A1O1Ixp33_ASAP7_75t_L g2783 ( 
.A1(n_2560),
.A2(n_1790),
.B(n_1792),
.C(n_1789),
.Y(n_2783)
);

O2A1O1Ixp33_ASAP7_75t_SL g2784 ( 
.A1(n_2561),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2601),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2744),
.Y(n_2786)
);

AOI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_2662),
.A2(n_2706),
.B(n_2734),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2679),
.B(n_2643),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2644),
.A2(n_2546),
.B(n_2528),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2656),
.A2(n_2552),
.B1(n_2577),
.B2(n_2576),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2652),
.B(n_2515),
.Y(n_2791)
);

AOI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2673),
.A2(n_2598),
.B(n_2558),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2677),
.A2(n_2567),
.B(n_2554),
.Y(n_2793)
);

BUFx2_ASAP7_75t_L g2794 ( 
.A(n_2740),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2640),
.B(n_2591),
.Y(n_2795)
);

AOI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2686),
.A2(n_2605),
.B(n_2586),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2645),
.B(n_2531),
.Y(n_2797)
);

AOI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2760),
.A2(n_2583),
.B(n_2608),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2649),
.B(n_2573),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2725),
.B(n_2507),
.Y(n_2800)
);

BUFx8_ASAP7_75t_L g2801 ( 
.A(n_2710),
.Y(n_2801)
);

OAI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2699),
.A2(n_2604),
.B(n_2575),
.Y(n_2802)
);

INVx3_ASAP7_75t_SL g2803 ( 
.A(n_2681),
.Y(n_2803)
);

OR2x6_ASAP7_75t_L g2804 ( 
.A(n_2687),
.B(n_2585),
.Y(n_2804)
);

OR2x6_ASAP7_75t_L g2805 ( 
.A(n_2743),
.B(n_2587),
.Y(n_2805)
);

HB1xp67_ASAP7_75t_L g2806 ( 
.A(n_2658),
.Y(n_2806)
);

AOI22xp33_ASAP7_75t_L g2807 ( 
.A1(n_2772),
.A2(n_2713),
.B1(n_2773),
.B2(n_2756),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2653),
.B(n_2532),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2684),
.B(n_2535),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2701),
.Y(n_2810)
);

A2O1A1Ixp33_ASAP7_75t_L g2811 ( 
.A1(n_2690),
.A2(n_2542),
.B(n_2599),
.C(n_2596),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2648),
.Y(n_2812)
);

AOI22xp33_ASAP7_75t_L g2813 ( 
.A1(n_2746),
.A2(n_2602),
.B1(n_2611),
.B2(n_1798),
.Y(n_2813)
);

BUFx3_ASAP7_75t_L g2814 ( 
.A(n_2715),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2766),
.B(n_1797),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_SL g2816 ( 
.A(n_2738),
.B(n_1810),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2723),
.B(n_1812),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2728),
.B(n_1814),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2729),
.B(n_1818),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2745),
.B(n_1820),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2755),
.B(n_1821),
.Y(n_2821)
);

INVx5_ASAP7_75t_L g2822 ( 
.A(n_2692),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2709),
.B(n_2665),
.Y(n_2823)
);

CKINVDCx6p67_ASAP7_75t_R g2824 ( 
.A(n_2722),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2727),
.A2(n_1825),
.B(n_1824),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2669),
.B(n_1827),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_R g2827 ( 
.A(n_2696),
.B(n_1828),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_2767),
.B(n_1830),
.Y(n_2828)
);

INVx3_ASAP7_75t_SL g2829 ( 
.A(n_2758),
.Y(n_2829)
);

OAI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2771),
.A2(n_1833),
.B(n_1831),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2670),
.B(n_1841),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2722),
.B(n_2675),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2748),
.B(n_1842),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2650),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2651),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2717),
.B(n_1852),
.Y(n_2836)
);

BUFx6f_ASAP7_75t_L g2837 ( 
.A(n_2692),
.Y(n_2837)
);

AO32x2_ASAP7_75t_L g2838 ( 
.A1(n_2695),
.A2(n_6),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2708),
.B(n_1853),
.Y(n_2839)
);

A2O1A1Ixp33_ASAP7_75t_SL g2840 ( 
.A1(n_2750),
.A2(n_1855),
.B(n_1854),
.C(n_6),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_SL g2841 ( 
.A(n_2689),
.B(n_325),
.Y(n_2841)
);

A2O1A1Ixp33_ASAP7_75t_L g2842 ( 
.A1(n_2657),
.A2(n_7),
.B(n_4),
.C(n_5),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2659),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2730),
.B(n_5),
.Y(n_2844)
);

BUFx2_ASAP7_75t_L g2845 ( 
.A(n_2714),
.Y(n_2845)
);

OR2x2_ASAP7_75t_L g2846 ( 
.A(n_2654),
.B(n_8),
.Y(n_2846)
);

A2O1A1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2672),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_2847)
);

AOI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2776),
.A2(n_327),
.B(n_326),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2663),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2741),
.B(n_326),
.Y(n_2850)
);

AOI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2707),
.A2(n_328),
.B(n_327),
.Y(n_2851)
);

OAI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2749),
.A2(n_330),
.B1(n_331),
.B2(n_329),
.Y(n_2852)
);

BUFx2_ASAP7_75t_SL g2853 ( 
.A(n_2758),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_R g2854 ( 
.A(n_2751),
.B(n_2719),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2762),
.B(n_2781),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2668),
.Y(n_2856)
);

INVxp67_ASAP7_75t_SL g2857 ( 
.A(n_2757),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2683),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2666),
.A2(n_334),
.B(n_333),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2691),
.B(n_11),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2754),
.A2(n_2642),
.B(n_2770),
.Y(n_2861)
);

NAND2x1p5_ASAP7_75t_L g2862 ( 
.A(n_2777),
.B(n_335),
.Y(n_2862)
);

INVxp67_ASAP7_75t_L g2863 ( 
.A(n_2739),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2693),
.B(n_12),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2718),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_2697),
.B(n_13),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2698),
.B(n_13),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_L g2868 ( 
.A(n_2726),
.B(n_337),
.Y(n_2868)
);

CKINVDCx14_ASAP7_75t_R g2869 ( 
.A(n_2716),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2704),
.B(n_14),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2747),
.A2(n_340),
.B(n_339),
.Y(n_2871)
);

AO21x1_ASAP7_75t_L g2872 ( 
.A1(n_2676),
.A2(n_340),
.B(n_339),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2759),
.A2(n_344),
.B(n_341),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2785),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2712),
.A2(n_347),
.B(n_346),
.Y(n_2875)
);

OAI22x1_ASAP7_75t_L g2876 ( 
.A1(n_2639),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2647),
.B(n_16),
.Y(n_2877)
);

AOI22xp33_ASAP7_75t_L g2878 ( 
.A1(n_2761),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2674),
.B(n_19),
.Y(n_2879)
);

A2O1A1Ixp33_ASAP7_75t_L g2880 ( 
.A1(n_2711),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_2880)
);

O2A1O1Ixp33_ASAP7_75t_L g2881 ( 
.A1(n_2763),
.A2(n_349),
.B(n_350),
.C(n_348),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2753),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2768),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2769),
.B(n_349),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2655),
.A2(n_351),
.B(n_350),
.Y(n_2885)
);

CKINVDCx8_ASAP7_75t_R g2886 ( 
.A(n_2688),
.Y(n_2886)
);

O2A1O1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_2646),
.A2(n_353),
.B(n_354),
.C(n_352),
.Y(n_2887)
);

OAI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2775),
.A2(n_2779),
.B1(n_2778),
.B2(n_2733),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2774),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2783),
.B(n_355),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2700),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2780),
.Y(n_2892)
);

AOI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2680),
.A2(n_357),
.B1(n_358),
.B2(n_356),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2732),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_SL g2895 ( 
.A(n_2764),
.B(n_357),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2660),
.A2(n_359),
.B(n_358),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2737),
.Y(n_2897)
);

O2A1O1Ixp5_ASAP7_75t_L g2898 ( 
.A1(n_2721),
.A2(n_2671),
.B(n_2664),
.C(n_2682),
.Y(n_2898)
);

O2A1O1Ixp33_ASAP7_75t_L g2899 ( 
.A1(n_2702),
.A2(n_360),
.B(n_361),
.C(n_359),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2678),
.B(n_24),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2782),
.Y(n_2901)
);

AOI21x1_ASAP7_75t_L g2902 ( 
.A1(n_2685),
.A2(n_361),
.B(n_360),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_L g2903 ( 
.A1(n_2735),
.A2(n_363),
.B1(n_364),
.B2(n_362),
.Y(n_2903)
);

OR2x6_ASAP7_75t_SL g2904 ( 
.A(n_2784),
.B(n_2661),
.Y(n_2904)
);

O2A1O1Ixp33_ASAP7_75t_L g2905 ( 
.A1(n_2667),
.A2(n_368),
.B(n_369),
.C(n_367),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2720),
.A2(n_369),
.B(n_367),
.Y(n_2906)
);

AOI22xp5_ASAP7_75t_L g2907 ( 
.A1(n_2731),
.A2(n_372),
.B1(n_373),
.B2(n_371),
.Y(n_2907)
);

INVx4_ASAP7_75t_L g2908 ( 
.A(n_2724),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2752),
.B(n_2742),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2703),
.B(n_371),
.Y(n_2910)
);

INVx3_ASAP7_75t_L g2911 ( 
.A(n_2736),
.Y(n_2911)
);

BUFx10_ASAP7_75t_L g2912 ( 
.A(n_2705),
.Y(n_2912)
);

O2A1O1Ixp33_ASAP7_75t_L g2913 ( 
.A1(n_2694),
.A2(n_375),
.B(n_376),
.C(n_374),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2641),
.A2(n_379),
.B1(n_380),
.B2(n_377),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2641),
.B(n_28),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2641),
.B(n_29),
.Y(n_2916)
);

A2O1A1Ixp33_ASAP7_75t_L g2917 ( 
.A1(n_2641),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2765),
.B(n_381),
.Y(n_2918)
);

BUFx6f_ASAP7_75t_L g2919 ( 
.A(n_2740),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_2740),
.Y(n_2920)
);

BUFx6f_ASAP7_75t_L g2921 ( 
.A(n_2740),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2641),
.B(n_29),
.Y(n_2922)
);

OR2x6_ASAP7_75t_L g2923 ( 
.A(n_2740),
.B(n_382),
.Y(n_2923)
);

AOI21x1_ASAP7_75t_L g2924 ( 
.A1(n_2644),
.A2(n_384),
.B(n_383),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2765),
.B(n_383),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2641),
.B(n_384),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2641),
.A2(n_387),
.B1(n_388),
.B2(n_386),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2765),
.B(n_389),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2662),
.A2(n_391),
.B(n_390),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2662),
.A2(n_392),
.B(n_391),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2740),
.Y(n_2931)
);

INVxp67_ASAP7_75t_SL g2932 ( 
.A(n_2806),
.Y(n_2932)
);

AO31x2_ASAP7_75t_L g2933 ( 
.A1(n_2787),
.A2(n_36),
.A3(n_34),
.B(n_35),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2807),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2823),
.B(n_35),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2791),
.B(n_37),
.Y(n_2936)
);

OAI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2855),
.A2(n_38),
.B(n_39),
.Y(n_2937)
);

OA21x2_ASAP7_75t_L g2938 ( 
.A1(n_2892),
.A2(n_38),
.B(n_39),
.Y(n_2938)
);

AOI211x1_ASAP7_75t_L g2939 ( 
.A1(n_2929),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2829),
.Y(n_2940)
);

INVx3_ASAP7_75t_L g2941 ( 
.A(n_2814),
.Y(n_2941)
);

A2O1A1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2802),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_2942)
);

OAI21xp5_ASAP7_75t_SL g2943 ( 
.A1(n_2821),
.A2(n_43),
.B(n_45),
.Y(n_2943)
);

AOI221xp5_ASAP7_75t_L g2944 ( 
.A1(n_2926),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_2944)
);

OAI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2869),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_2945)
);

INVx4_ASAP7_75t_L g2946 ( 
.A(n_2822),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_2886),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2799),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_2948)
);

CKINVDCx8_ASAP7_75t_R g2949 ( 
.A(n_2853),
.Y(n_2949)
);

OAI21x1_ASAP7_75t_SL g2950 ( 
.A1(n_2796),
.A2(n_50),
.B(n_51),
.Y(n_2950)
);

NOR3xp33_ASAP7_75t_L g2951 ( 
.A(n_2795),
.B(n_50),
.C(n_51),
.Y(n_2951)
);

AOI21xp33_ASAP7_75t_L g2952 ( 
.A1(n_2830),
.A2(n_50),
.B(n_51),
.Y(n_2952)
);

O2A1O1Ixp5_ASAP7_75t_L g2953 ( 
.A1(n_2890),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_2953)
);

AOI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2884),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.Y(n_2954)
);

OAI21x1_ASAP7_75t_SL g2955 ( 
.A1(n_2872),
.A2(n_56),
.B(n_57),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2808),
.B(n_57),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2797),
.B(n_394),
.Y(n_2957)
);

OA22x2_ASAP7_75t_L g2958 ( 
.A1(n_2923),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2958)
);

BUFx12f_ASAP7_75t_L g2959 ( 
.A(n_2801),
.Y(n_2959)
);

OAI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2813),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2960)
);

A2O1A1Ixp33_ASAP7_75t_L g2961 ( 
.A1(n_2909),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2809),
.B(n_395),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2818),
.B(n_63),
.Y(n_2963)
);

OR2x2_ASAP7_75t_L g2964 ( 
.A(n_2915),
.B(n_2916),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2819),
.B(n_64),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2789),
.A2(n_64),
.B(n_65),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_SL g2967 ( 
.A1(n_2923),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2817),
.B(n_2820),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2833),
.B(n_66),
.Y(n_2969)
);

AOI211x1_ASAP7_75t_L g2970 ( 
.A1(n_2930),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_2970)
);

AO21x2_ASAP7_75t_L g2971 ( 
.A1(n_2924),
.A2(n_67),
.B(n_68),
.Y(n_2971)
);

AOI22xp33_ASAP7_75t_L g2972 ( 
.A1(n_2868),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_2803),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2844),
.B(n_71),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2836),
.B(n_72),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_SL g2976 ( 
.A(n_2790),
.B(n_396),
.Y(n_2976)
);

OAI21x1_ASAP7_75t_L g2977 ( 
.A1(n_2861),
.A2(n_73),
.B(n_74),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2860),
.B(n_74),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2922),
.B(n_397),
.Y(n_2979)
);

OAI21x1_ASAP7_75t_L g2980 ( 
.A1(n_2798),
.A2(n_74),
.B(n_75),
.Y(n_2980)
);

BUFx6f_ASAP7_75t_L g2981 ( 
.A(n_2837),
.Y(n_2981)
);

OAI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2898),
.A2(n_75),
.B(n_76),
.Y(n_2982)
);

OR2x6_ASAP7_75t_L g2983 ( 
.A(n_2919),
.B(n_398),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2864),
.B(n_75),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2822),
.Y(n_2985)
);

AOI21xp33_ASAP7_75t_L g2986 ( 
.A1(n_2888),
.A2(n_76),
.B(n_77),
.Y(n_2986)
);

NAND3xp33_ASAP7_75t_L g2987 ( 
.A(n_2910),
.B(n_77),
.C(n_78),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2786),
.Y(n_2988)
);

OAI21x1_ASAP7_75t_L g2989 ( 
.A1(n_2897),
.A2(n_77),
.B(n_78),
.Y(n_2989)
);

INVxp67_ASAP7_75t_SL g2990 ( 
.A(n_2883),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2793),
.A2(n_400),
.B(n_399),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_SL g2992 ( 
.A1(n_2811),
.A2(n_403),
.B(n_401),
.Y(n_2992)
);

OAI22x1_ASAP7_75t_L g2993 ( 
.A1(n_2927),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2993)
);

OAI21x1_ASAP7_75t_L g2994 ( 
.A1(n_2911),
.A2(n_79),
.B(n_81),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2849),
.Y(n_2995)
);

AO32x2_ASAP7_75t_L g2996 ( 
.A1(n_2914),
.A2(n_84),
.A3(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2867),
.B(n_82),
.Y(n_2997)
);

OAI21xp33_ASAP7_75t_L g2998 ( 
.A1(n_2878),
.A2(n_84),
.B(n_85),
.Y(n_2998)
);

INVx3_ASAP7_75t_SL g2999 ( 
.A(n_2919),
.Y(n_2999)
);

O2A1O1Ixp33_ASAP7_75t_L g3000 ( 
.A1(n_2840),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_3000)
);

OAI21x1_ASAP7_75t_SL g3001 ( 
.A1(n_2881),
.A2(n_86),
.B(n_87),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2792),
.A2(n_405),
.B(n_404),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2870),
.B(n_86),
.Y(n_3003)
);

NAND2x1p5_ASAP7_75t_L g3004 ( 
.A(n_2822),
.B(n_406),
.Y(n_3004)
);

BUFx3_ASAP7_75t_L g3005 ( 
.A(n_2920),
.Y(n_3005)
);

OAI22x1_ASAP7_75t_L g3006 ( 
.A1(n_2893),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_3006)
);

INVx3_ASAP7_75t_L g3007 ( 
.A(n_2788),
.Y(n_3007)
);

OAI21x1_ASAP7_75t_SL g3008 ( 
.A1(n_2902),
.A2(n_91),
.B(n_92),
.Y(n_3008)
);

OAI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2826),
.A2(n_93),
.B(n_94),
.Y(n_3009)
);

OA21x2_ASAP7_75t_L g3010 ( 
.A1(n_2851),
.A2(n_94),
.B(n_95),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2831),
.A2(n_96),
.B(n_97),
.Y(n_3011)
);

AO31x2_ASAP7_75t_L g3012 ( 
.A1(n_2908),
.A2(n_98),
.A3(n_96),
.B(n_97),
.Y(n_3012)
);

O2A1O1Ixp33_ASAP7_75t_SL g3013 ( 
.A1(n_2842),
.A2(n_408),
.B(n_409),
.C(n_407),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2839),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2900),
.B(n_98),
.Y(n_3015)
);

INVx3_ASAP7_75t_L g3016 ( 
.A(n_2824),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2856),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2863),
.B(n_101),
.Y(n_3018)
);

INVx4_ASAP7_75t_SL g3019 ( 
.A(n_2921),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2845),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2846),
.B(n_102),
.Y(n_3021)
);

INVx8_ASAP7_75t_L g3022 ( 
.A(n_2921),
.Y(n_3022)
);

NAND3x1_ASAP7_75t_L g3023 ( 
.A(n_2800),
.B(n_103),
.C(n_104),
.Y(n_3023)
);

CKINVDCx20_ASAP7_75t_R g3024 ( 
.A(n_2901),
.Y(n_3024)
);

OAI21x1_ASAP7_75t_L g3025 ( 
.A1(n_2891),
.A2(n_103),
.B(n_105),
.Y(n_3025)
);

BUFx8_ASAP7_75t_L g3026 ( 
.A(n_2794),
.Y(n_3026)
);

BUFx2_ASAP7_75t_L g3027 ( 
.A(n_2857),
.Y(n_3027)
);

O2A1O1Ixp33_ASAP7_75t_SL g3028 ( 
.A1(n_2847),
.A2(n_412),
.B(n_413),
.C(n_411),
.Y(n_3028)
);

NOR2x1_ASAP7_75t_SL g3029 ( 
.A(n_2832),
.B(n_411),
.Y(n_3029)
);

NAND3xp33_ASAP7_75t_L g3030 ( 
.A(n_2889),
.B(n_105),
.C(n_106),
.Y(n_3030)
);

AOI21x1_ASAP7_75t_SL g3031 ( 
.A1(n_2877),
.A2(n_105),
.B(n_106),
.Y(n_3031)
);

OAI21x1_ASAP7_75t_L g3032 ( 
.A1(n_2859),
.A2(n_2894),
.B(n_2848),
.Y(n_3032)
);

OA22x2_ASAP7_75t_L g3033 ( 
.A1(n_2876),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3033)
);

A2O1A1Ixp33_ASAP7_75t_L g3034 ( 
.A1(n_2873),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2815),
.B(n_412),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2810),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2866),
.B(n_110),
.Y(n_3037)
);

INVxp67_ASAP7_75t_L g3038 ( 
.A(n_2874),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2812),
.B(n_110),
.Y(n_3039)
);

AOI221x1_ASAP7_75t_L g3040 ( 
.A1(n_2880),
.A2(n_416),
.B1(n_417),
.B2(n_415),
.C(n_414),
.Y(n_3040)
);

NOR4xp25_ASAP7_75t_L g3041 ( 
.A(n_2887),
.B(n_2899),
.C(n_2913),
.D(n_2905),
.Y(n_3041)
);

AOI21x1_ASAP7_75t_SL g3042 ( 
.A1(n_2879),
.A2(n_111),
.B(n_112),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2850),
.A2(n_417),
.B(n_416),
.Y(n_3043)
);

AO31x2_ASAP7_75t_L g3044 ( 
.A1(n_2917),
.A2(n_114),
.A3(n_111),
.B(n_113),
.Y(n_3044)
);

INVx6_ASAP7_75t_L g3045 ( 
.A(n_2931),
.Y(n_3045)
);

O2A1O1Ixp5_ASAP7_75t_SL g3046 ( 
.A1(n_2903),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_3046)
);

OAI21x1_ASAP7_75t_L g3047 ( 
.A1(n_2871),
.A2(n_116),
.B(n_117),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2834),
.B(n_116),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2835),
.B(n_2843),
.Y(n_3049)
);

OR2x6_ASAP7_75t_L g3050 ( 
.A(n_2805),
.B(n_419),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2858),
.B(n_118),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2865),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2841),
.B(n_119),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2828),
.A2(n_422),
.B(n_420),
.Y(n_3054)
);

AO22x2_ASAP7_75t_L g3055 ( 
.A1(n_2852),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2968),
.B(n_2912),
.Y(n_3056)
);

AO21x2_ASAP7_75t_L g3057 ( 
.A1(n_2982),
.A2(n_2875),
.B(n_2906),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_2964),
.B(n_2882),
.Y(n_3058)
);

AND2x4_ASAP7_75t_SL g3059 ( 
.A(n_2973),
.B(n_2804),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_L g3060 ( 
.A(n_2949),
.Y(n_3060)
);

OAI21x1_ASAP7_75t_L g3061 ( 
.A1(n_3032),
.A2(n_2896),
.B(n_2885),
.Y(n_3061)
);

OR2x6_ASAP7_75t_L g3062 ( 
.A(n_3022),
.B(n_2804),
.Y(n_3062)
);

BUFx12f_ASAP7_75t_L g3063 ( 
.A(n_2959),
.Y(n_3063)
);

OAI21x1_ASAP7_75t_L g3064 ( 
.A1(n_2977),
.A2(n_2966),
.B(n_2980),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2932),
.B(n_2918),
.Y(n_3065)
);

AO21x2_ASAP7_75t_L g3066 ( 
.A1(n_3008),
.A2(n_2825),
.B(n_2895),
.Y(n_3066)
);

OAI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_2936),
.A2(n_2904),
.B1(n_2907),
.B2(n_2925),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2940),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2957),
.B(n_2928),
.Y(n_3069)
);

OAI21x1_ASAP7_75t_L g3070 ( 
.A1(n_2994),
.A2(n_2816),
.B(n_2862),
.Y(n_3070)
);

OAI21x1_ASAP7_75t_L g3071 ( 
.A1(n_2989),
.A2(n_3002),
.B(n_3047),
.Y(n_3071)
);

OAI21x1_ASAP7_75t_L g3072 ( 
.A1(n_2991),
.A2(n_2838),
.B(n_2854),
.Y(n_3072)
);

INVx4_ASAP7_75t_SL g3073 ( 
.A(n_2999),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2935),
.B(n_2827),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2988),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2952),
.A2(n_424),
.B(n_423),
.Y(n_3076)
);

INVx1_ASAP7_75t_SL g3077 ( 
.A(n_3020),
.Y(n_3077)
);

O2A1O1Ixp33_ASAP7_75t_SL g3078 ( 
.A1(n_2942),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_3078)
);

BUFx8_ASAP7_75t_L g3079 ( 
.A(n_3005),
.Y(n_3079)
);

NAND3x1_ASAP7_75t_L g3080 ( 
.A(n_2951),
.B(n_124),
.C(n_125),
.Y(n_3080)
);

BUFx2_ASAP7_75t_R g3081 ( 
.A(n_2947),
.Y(n_3081)
);

HB1xp67_ASAP7_75t_L g3082 ( 
.A(n_3027),
.Y(n_3082)
);

AOI222xp33_ASAP7_75t_L g3083 ( 
.A1(n_2967),
.A2(n_2998),
.B1(n_2943),
.B2(n_3011),
.C1(n_3009),
.C2(n_2937),
.Y(n_3083)
);

OA21x2_ASAP7_75t_L g3084 ( 
.A1(n_3040),
.A2(n_126),
.B(n_127),
.Y(n_3084)
);

OAI221xp5_ASAP7_75t_L g3085 ( 
.A1(n_3035),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.C(n_130),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3036),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2990),
.B(n_425),
.Y(n_3087)
);

INVx3_ASAP7_75t_L g3088 ( 
.A(n_2941),
.Y(n_3088)
);

OAI221xp5_ASAP7_75t_L g3089 ( 
.A1(n_2934),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.C(n_134),
.Y(n_3089)
);

OAI21x1_ASAP7_75t_L g3090 ( 
.A1(n_3025),
.A2(n_131),
.B(n_132),
.Y(n_3090)
);

CKINVDCx20_ASAP7_75t_R g3091 ( 
.A(n_3024),
.Y(n_3091)
);

OAI21x1_ASAP7_75t_L g3092 ( 
.A1(n_2950),
.A2(n_132),
.B(n_133),
.Y(n_3092)
);

OAI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_3041),
.A2(n_134),
.B(n_135),
.Y(n_3093)
);

OR2x6_ASAP7_75t_L g3094 ( 
.A(n_3050),
.B(n_426),
.Y(n_3094)
);

OAI21x1_ASAP7_75t_L g3095 ( 
.A1(n_3031),
.A2(n_136),
.B(n_137),
.Y(n_3095)
);

OAI21x1_ASAP7_75t_L g3096 ( 
.A1(n_3042),
.A2(n_136),
.B(n_137),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2995),
.Y(n_3097)
);

INVx1_ASAP7_75t_SL g3098 ( 
.A(n_3007),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_2979),
.B(n_428),
.Y(n_3099)
);

AOI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2987),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_3017),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_SL g3102 ( 
.A(n_2956),
.B(n_429),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2962),
.B(n_429),
.Y(n_3103)
);

CKINVDCx20_ASAP7_75t_R g3104 ( 
.A(n_3026),
.Y(n_3104)
);

INVx4_ASAP7_75t_L g3105 ( 
.A(n_2985),
.Y(n_3105)
);

NAND2x1p5_ASAP7_75t_L g3106 ( 
.A(n_2946),
.B(n_430),
.Y(n_3106)
);

INVxp67_ASAP7_75t_SL g3107 ( 
.A(n_3049),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_SL g3108 ( 
.A1(n_3030),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_3033),
.B(n_431),
.Y(n_3109)
);

O2A1O1Ixp33_ASAP7_75t_SL g3110 ( 
.A1(n_2961),
.A2(n_3034),
.B(n_2976),
.C(n_2944),
.Y(n_3110)
);

OA21x2_ASAP7_75t_L g3111 ( 
.A1(n_2953),
.A2(n_144),
.B(n_145),
.Y(n_3111)
);

AO31x2_ASAP7_75t_L g3112 ( 
.A1(n_2993),
.A2(n_148),
.A3(n_145),
.B(n_147),
.Y(n_3112)
);

AOI22xp33_ASAP7_75t_L g3113 ( 
.A1(n_2960),
.A2(n_148),
.B1(n_145),
.B2(n_147),
.Y(n_3113)
);

INVxp67_ASAP7_75t_SL g3114 ( 
.A(n_3052),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2963),
.B(n_432),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_2965),
.B(n_3038),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2955),
.A2(n_149),
.B(n_150),
.Y(n_3117)
);

NAND3xp33_ASAP7_75t_L g3118 ( 
.A(n_2972),
.B(n_2954),
.C(n_2986),
.Y(n_3118)
);

OAI21x1_ASAP7_75t_L g3119 ( 
.A1(n_3001),
.A2(n_149),
.B(n_150),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_3015),
.B(n_433),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2933),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2981),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_3014),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_3123)
);

AO21x1_ASAP7_75t_L g3124 ( 
.A1(n_3000),
.A2(n_151),
.B(n_152),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2992),
.A2(n_434),
.B(n_433),
.Y(n_3125)
);

AO32x2_ASAP7_75t_L g3126 ( 
.A1(n_2948),
.A2(n_156),
.A3(n_153),
.B1(n_155),
.B2(n_157),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2933),
.Y(n_3127)
);

OAI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_3046),
.A2(n_153),
.B(n_155),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_3006),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2971),
.Y(n_3130)
);

AO31x2_ASAP7_75t_L g3131 ( 
.A1(n_3029),
.A2(n_159),
.A3(n_157),
.B(n_158),
.Y(n_3131)
);

AOI221xp5_ASAP7_75t_L g3132 ( 
.A1(n_3013),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.C(n_161),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3012),
.Y(n_3133)
);

AOI221xp5_ASAP7_75t_L g3134 ( 
.A1(n_3028),
.A2(n_2945),
.B1(n_2939),
.B2(n_2970),
.C(n_2974),
.Y(n_3134)
);

OAI21x1_ASAP7_75t_L g3135 ( 
.A1(n_3010),
.A2(n_159),
.B(n_160),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2938),
.Y(n_3136)
);

AO31x2_ASAP7_75t_L g3137 ( 
.A1(n_3043),
.A2(n_163),
.A3(n_161),
.B(n_162),
.Y(n_3137)
);

OAI221xp5_ASAP7_75t_L g3138 ( 
.A1(n_2975),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_3075),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_3107),
.B(n_2978),
.Y(n_3140)
);

OR2x6_ASAP7_75t_L g3141 ( 
.A(n_3060),
.B(n_3045),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_3114),
.B(n_2984),
.Y(n_3142)
);

OAI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_3125),
.A2(n_3054),
.B(n_2997),
.Y(n_3143)
);

OAI21x1_ASAP7_75t_L g3144 ( 
.A1(n_3061),
.A2(n_3048),
.B(n_3039),
.Y(n_3144)
);

OAI21x1_ASAP7_75t_L g3145 ( 
.A1(n_3064),
.A2(n_3051),
.B(n_3003),
.Y(n_3145)
);

AOI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_3056),
.A2(n_3055),
.B(n_3053),
.Y(n_3146)
);

NAND2x1p5_ASAP7_75t_L g3147 ( 
.A(n_3077),
.B(n_3016),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_3082),
.B(n_3019),
.Y(n_3148)
);

BUFx12f_ASAP7_75t_L g3149 ( 
.A(n_3063),
.Y(n_3149)
);

AOI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_3057),
.A2(n_3055),
.B(n_2969),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_3071),
.A2(n_3004),
.B(n_3023),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3086),
.Y(n_3152)
);

AO21x2_ASAP7_75t_L g3153 ( 
.A1(n_3121),
.A2(n_3127),
.B(n_3133),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_3058),
.B(n_3037),
.Y(n_3154)
);

OA21x2_ASAP7_75t_L g3155 ( 
.A1(n_3072),
.A2(n_3021),
.B(n_3018),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_3110),
.A2(n_2958),
.B(n_2996),
.Y(n_3156)
);

OR2x6_ASAP7_75t_L g3157 ( 
.A(n_3060),
.B(n_2983),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_3130),
.Y(n_3158)
);

OR2x2_ASAP7_75t_L g3159 ( 
.A(n_3065),
.B(n_3044),
.Y(n_3159)
);

INVxp67_ASAP7_75t_L g3160 ( 
.A(n_3116),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_3084),
.A2(n_165),
.B(n_166),
.Y(n_3161)
);

AOI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_3083),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_3162)
);

BUFx2_ASAP7_75t_L g3163 ( 
.A(n_3062),
.Y(n_3163)
);

OA21x2_ASAP7_75t_L g3164 ( 
.A1(n_3135),
.A2(n_169),
.B(n_170),
.Y(n_3164)
);

AO31x2_ASAP7_75t_L g3165 ( 
.A1(n_3136),
.A2(n_171),
.A3(n_169),
.B(n_170),
.Y(n_3165)
);

INVx2_ASAP7_75t_SL g3166 ( 
.A(n_3059),
.Y(n_3166)
);

OAI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_3076),
.A2(n_170),
.B(n_171),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_3078),
.A2(n_171),
.B(n_172),
.Y(n_3168)
);

AO31x2_ASAP7_75t_L g3169 ( 
.A1(n_3124),
.A2(n_3067),
.A3(n_3101),
.B(n_3097),
.Y(n_3169)
);

AO31x2_ASAP7_75t_L g3170 ( 
.A1(n_3087),
.A2(n_174),
.A3(n_172),
.B(n_173),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_L g3171 ( 
.A(n_3074),
.B(n_437),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3069),
.B(n_438),
.Y(n_3172)
);

OAI21x1_ASAP7_75t_L g3173 ( 
.A1(n_3090),
.A2(n_173),
.B(n_174),
.Y(n_3173)
);

BUFx2_ASAP7_75t_L g3174 ( 
.A(n_3062),
.Y(n_3174)
);

OA21x2_ASAP7_75t_L g3175 ( 
.A1(n_3095),
.A2(n_3096),
.B(n_3092),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_3109),
.B(n_439),
.Y(n_3176)
);

BUFx2_ASAP7_75t_SL g3177 ( 
.A(n_3091),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_3115),
.B(n_440),
.Y(n_3178)
);

AOI21xp5_ASAP7_75t_L g3179 ( 
.A1(n_3132),
.A2(n_177),
.B(n_178),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_3099),
.B(n_440),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_3102),
.B(n_441),
.Y(n_3181)
);

BUFx2_ASAP7_75t_L g3182 ( 
.A(n_3068),
.Y(n_3182)
);

INVx3_ASAP7_75t_L g3183 ( 
.A(n_3122),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_3120),
.B(n_441),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3137),
.Y(n_3185)
);

AO31x2_ASAP7_75t_L g3186 ( 
.A1(n_3103),
.A2(n_183),
.A3(n_181),
.B(n_182),
.Y(n_3186)
);

OAI21x1_ASAP7_75t_L g3187 ( 
.A1(n_3070),
.A2(n_181),
.B(n_182),
.Y(n_3187)
);

AO31x2_ASAP7_75t_L g3188 ( 
.A1(n_3105),
.A2(n_184),
.A3(n_182),
.B(n_183),
.Y(n_3188)
);

INVx5_ASAP7_75t_L g3189 ( 
.A(n_3094),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_3131),
.Y(n_3190)
);

OA21x2_ASAP7_75t_L g3191 ( 
.A1(n_3117),
.A2(n_184),
.B(n_185),
.Y(n_3191)
);

OA21x2_ASAP7_75t_L g3192 ( 
.A1(n_3093),
.A2(n_186),
.B(n_187),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_3098),
.B(n_443),
.Y(n_3193)
);

BUFx3_ASAP7_75t_L g3194 ( 
.A(n_3079),
.Y(n_3194)
);

OAI21x1_ASAP7_75t_L g3195 ( 
.A1(n_3119),
.A2(n_186),
.B(n_188),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_3134),
.B(n_444),
.Y(n_3196)
);

OAI21x1_ASAP7_75t_L g3197 ( 
.A1(n_3128),
.A2(n_188),
.B(n_189),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3111),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_3073),
.B(n_444),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3118),
.A2(n_188),
.B(n_189),
.Y(n_3200)
);

OA21x2_ASAP7_75t_L g3201 ( 
.A1(n_3100),
.A2(n_190),
.B(n_191),
.Y(n_3201)
);

OAI21x1_ASAP7_75t_L g3202 ( 
.A1(n_3106),
.A2(n_190),
.B(n_191),
.Y(n_3202)
);

OR2x2_ASAP7_75t_L g3203 ( 
.A(n_3112),
.B(n_445),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_3066),
.A2(n_192),
.B(n_193),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3129),
.B(n_445),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3089),
.A2(n_3080),
.B1(n_3108),
.B2(n_3085),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3088),
.B(n_446),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3126),
.Y(n_3208)
);

BUFx2_ASAP7_75t_L g3209 ( 
.A(n_3073),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3163),
.B(n_3174),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3139),
.Y(n_3211)
);

BUFx2_ASAP7_75t_L g3212 ( 
.A(n_3209),
.Y(n_3212)
);

OA21x2_ASAP7_75t_L g3213 ( 
.A1(n_3150),
.A2(n_3138),
.B(n_3123),
.Y(n_3213)
);

HB1xp67_ASAP7_75t_L g3214 ( 
.A(n_3159),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3152),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_3160),
.B(n_3081),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3140),
.B(n_3113),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3142),
.B(n_447),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3166),
.B(n_3104),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3158),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3190),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3153),
.Y(n_3222)
);

OR2x2_ASAP7_75t_L g3223 ( 
.A(n_3154),
.B(n_448),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3185),
.Y(n_3224)
);

BUFx3_ASAP7_75t_L g3225 ( 
.A(n_3149),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3198),
.Y(n_3226)
);

CKINVDCx5p33_ASAP7_75t_R g3227 ( 
.A(n_3177),
.Y(n_3227)
);

BUFx3_ASAP7_75t_L g3228 ( 
.A(n_3141),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3165),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3165),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3145),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3170),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3170),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_3144),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3208),
.Y(n_3235)
);

BUFx6f_ASAP7_75t_L g3236 ( 
.A(n_3183),
.Y(n_3236)
);

OR2x6_ASAP7_75t_L g3237 ( 
.A(n_3151),
.B(n_449),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3186),
.Y(n_3238)
);

INVx4_ASAP7_75t_L g3239 ( 
.A(n_3157),
.Y(n_3239)
);

INVx1_ASAP7_75t_SL g3240 ( 
.A(n_3189),
.Y(n_3240)
);

BUFx2_ASAP7_75t_L g3241 ( 
.A(n_3155),
.Y(n_3241)
);

INVx5_ASAP7_75t_L g3242 ( 
.A(n_3199),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3176),
.B(n_450),
.Y(n_3243)
);

INVx3_ASAP7_75t_L g3244 ( 
.A(n_3189),
.Y(n_3244)
);

AO21x2_ASAP7_75t_L g3245 ( 
.A1(n_3204),
.A2(n_195),
.B(n_196),
.Y(n_3245)
);

INVx4_ASAP7_75t_SL g3246 ( 
.A(n_3188),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3169),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3171),
.B(n_3193),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3187),
.Y(n_3249)
);

INVx3_ASAP7_75t_L g3250 ( 
.A(n_3207),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3146),
.B(n_452),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3175),
.Y(n_3252)
);

INVx1_ASAP7_75t_SL g3253 ( 
.A(n_3172),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3203),
.Y(n_3254)
);

HB1xp67_ASAP7_75t_L g3255 ( 
.A(n_3191),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3164),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_3180),
.Y(n_3257)
);

INVx3_ASAP7_75t_L g3258 ( 
.A(n_3202),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3173),
.Y(n_3259)
);

BUFx3_ASAP7_75t_L g3260 ( 
.A(n_3184),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3195),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3181),
.Y(n_3262)
);

CKINVDCx6p67_ASAP7_75t_R g3263 ( 
.A(n_3178),
.Y(n_3263)
);

HB1xp67_ASAP7_75t_L g3264 ( 
.A(n_3143),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_3156),
.B(n_453),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3192),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3197),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3161),
.Y(n_3268)
);

OAI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3200),
.A2(n_197),
.B(n_198),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3196),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3167),
.Y(n_3271)
);

INVx3_ASAP7_75t_L g3272 ( 
.A(n_3201),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3168),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3205),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3206),
.Y(n_3275)
);

OR2x2_ASAP7_75t_L g3276 ( 
.A(n_3179),
.B(n_455),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3162),
.B(n_456),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3182),
.B(n_458),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_3148),
.Y(n_3279)
);

INVxp33_ASAP7_75t_L g3280 ( 
.A(n_3147),
.Y(n_3280)
);

INVx4_ASAP7_75t_L g3281 ( 
.A(n_3194),
.Y(n_3281)
);

AOI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_3206),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_3282)
);

AOI22xp33_ASAP7_75t_L g3283 ( 
.A1(n_3213),
.A2(n_460),
.B1(n_461),
.B2(n_459),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3210),
.B(n_202),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3226),
.Y(n_3285)
);

AOI21xp33_ASAP7_75t_L g3286 ( 
.A1(n_3271),
.A2(n_3251),
.B(n_3268),
.Y(n_3286)
);

OR2x2_ASAP7_75t_L g3287 ( 
.A(n_3214),
.B(n_203),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_3211),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_3269),
.A2(n_464),
.B1(n_465),
.B2(n_463),
.Y(n_3289)
);

INVx4_ASAP7_75t_L g3290 ( 
.A(n_3227),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3273),
.A2(n_467),
.B1(n_468),
.B2(n_466),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3215),
.Y(n_3292)
);

AOI21xp33_ASAP7_75t_L g3293 ( 
.A1(n_3276),
.A2(n_3267),
.B(n_3266),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3254),
.B(n_469),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3279),
.B(n_204),
.Y(n_3295)
);

AOI211xp5_ASAP7_75t_SL g3296 ( 
.A1(n_3272),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_3296)
);

AO21x2_ASAP7_75t_L g3297 ( 
.A1(n_3222),
.A2(n_207),
.B(n_209),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3263),
.A2(n_471),
.B1(n_472),
.B2(n_470),
.Y(n_3298)
);

HB1xp67_ASAP7_75t_L g3299 ( 
.A(n_3241),
.Y(n_3299)
);

OAI21x1_ASAP7_75t_L g3300 ( 
.A1(n_3252),
.A2(n_210),
.B(n_211),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_3237),
.A2(n_3245),
.B1(n_3277),
.B2(n_3260),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3270),
.A2(n_213),
.B1(n_210),
.B2(n_212),
.Y(n_3302)
);

BUFx6f_ASAP7_75t_L g3303 ( 
.A(n_3236),
.Y(n_3303)
);

NAND3xp33_ASAP7_75t_L g3304 ( 
.A(n_3255),
.B(n_475),
.C(n_474),
.Y(n_3304)
);

OAI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_3240),
.A2(n_477),
.B1(n_478),
.B2(n_476),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_3280),
.B(n_3239),
.Y(n_3306)
);

AOI221xp5_ASAP7_75t_L g3307 ( 
.A1(n_3274),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_3307)
);

OAI22xp5_ASAP7_75t_SL g3308 ( 
.A1(n_3281),
.A2(n_3265),
.B1(n_3216),
.B2(n_3228),
.Y(n_3308)
);

INVx11_ASAP7_75t_L g3309 ( 
.A(n_3219),
.Y(n_3309)
);

AOI22xp33_ASAP7_75t_L g3310 ( 
.A1(n_3258),
.A2(n_482),
.B1(n_483),
.B2(n_480),
.Y(n_3310)
);

OAI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_3244),
.A2(n_484),
.B1(n_485),
.B2(n_483),
.Y(n_3311)
);

AOI221xp5_ASAP7_75t_L g3312 ( 
.A1(n_3232),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.C(n_222),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3262),
.B(n_486),
.Y(n_3313)
);

OAI22xp33_ASAP7_75t_L g3314 ( 
.A1(n_3253),
.A2(n_491),
.B1(n_492),
.B2(n_490),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_3257),
.A2(n_493),
.B1(n_494),
.B2(n_491),
.Y(n_3315)
);

OAI221xp5_ASAP7_75t_L g3316 ( 
.A1(n_3250),
.A2(n_3217),
.B1(n_3218),
.B2(n_3223),
.C(n_3233),
.Y(n_3316)
);

A2O1A1Ixp33_ASAP7_75t_L g3317 ( 
.A1(n_3256),
.A2(n_495),
.B(n_496),
.C(n_494),
.Y(n_3317)
);

OR2x2_ASAP7_75t_L g3318 ( 
.A(n_3235),
.B(n_223),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3224),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_3248),
.A2(n_500),
.B1(n_501),
.B2(n_499),
.Y(n_3320)
);

AO21x2_ASAP7_75t_L g3321 ( 
.A1(n_3247),
.A2(n_227),
.B(n_228),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_3261),
.A2(n_507),
.B1(n_508),
.B2(n_506),
.Y(n_3322)
);

CKINVDCx10_ASAP7_75t_R g3323 ( 
.A(n_3243),
.Y(n_3323)
);

OAI221xp5_ASAP7_75t_L g3324 ( 
.A1(n_3238),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.C(n_230),
.Y(n_3324)
);

HB1xp67_ASAP7_75t_L g3325 ( 
.A(n_3259),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3220),
.Y(n_3326)
);

AOI221xp5_ASAP7_75t_L g3327 ( 
.A1(n_3278),
.A2(n_232),
.B1(n_229),
.B2(n_231),
.C(n_233),
.Y(n_3327)
);

OAI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_3249),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3328)
);

AOI21x1_ASAP7_75t_L g3329 ( 
.A1(n_3221),
.A2(n_234),
.B(n_235),
.Y(n_3329)
);

OAI221xp5_ASAP7_75t_L g3330 ( 
.A1(n_3231),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3229),
.Y(n_3331)
);

AOI211xp5_ASAP7_75t_L g3332 ( 
.A1(n_3230),
.A2(n_3234),
.B(n_3246),
.C(n_240),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3226),
.Y(n_3333)
);

AOI221xp5_ASAP7_75t_L g3334 ( 
.A1(n_3264),
.A2(n_240),
.B1(n_237),
.B2(n_239),
.C(n_241),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3264),
.A2(n_511),
.B1(n_512),
.B2(n_510),
.Y(n_3335)
);

NAND3xp33_ASAP7_75t_L g3336 ( 
.A(n_3264),
.B(n_514),
.C(n_513),
.Y(n_3336)
);

BUFx2_ASAP7_75t_L g3337 ( 
.A(n_3212),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3210),
.B(n_241),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3264),
.B(n_514),
.Y(n_3339)
);

INVx4_ASAP7_75t_L g3340 ( 
.A(n_3227),
.Y(n_3340)
);

AOI221xp5_ASAP7_75t_L g3341 ( 
.A1(n_3264),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.C(n_246),
.Y(n_3341)
);

NOR2x1_ASAP7_75t_R g3342 ( 
.A(n_3242),
.B(n_245),
.Y(n_3342)
);

AOI22xp33_ASAP7_75t_L g3343 ( 
.A1(n_3264),
.A2(n_517),
.B1(n_518),
.B2(n_516),
.Y(n_3343)
);

NOR2x1_ASAP7_75t_SL g3344 ( 
.A(n_3237),
.B(n_246),
.Y(n_3344)
);

INVx4_ASAP7_75t_SL g3345 ( 
.A(n_3225),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3275),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3211),
.Y(n_3347)
);

NAND4xp25_ASAP7_75t_L g3348 ( 
.A(n_3282),
.B(n_250),
.C(n_248),
.D(n_249),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3264),
.B(n_519),
.Y(n_3349)
);

OA21x2_ASAP7_75t_L g3350 ( 
.A1(n_3241),
.A2(n_252),
.B(n_253),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3331),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3333),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3348),
.A2(n_522),
.B1(n_523),
.B2(n_521),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3286),
.B(n_521),
.Y(n_3354)
);

NOR2xp67_ASAP7_75t_L g3355 ( 
.A(n_3299),
.B(n_254),
.Y(n_3355)
);

INVx2_ASAP7_75t_SL g3356 ( 
.A(n_3309),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3306),
.B(n_256),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_3334),
.A2(n_526),
.B1(n_527),
.B2(n_524),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3293),
.B(n_527),
.Y(n_3359)
);

AOI22xp5_ASAP7_75t_L g3360 ( 
.A1(n_3341),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3288),
.Y(n_3361)
);

HB1xp67_ASAP7_75t_L g3362 ( 
.A(n_3325),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3326),
.B(n_530),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3292),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_3283),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_3365)
);

BUFx2_ASAP7_75t_L g3366 ( 
.A(n_3345),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_3345),
.B(n_530),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3332),
.B(n_531),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3347),
.B(n_261),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3319),
.Y(n_3370)
);

BUFx12f_ASAP7_75t_L g3371 ( 
.A(n_3290),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3318),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3350),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3339),
.B(n_532),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3303),
.B(n_3284),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3350),
.Y(n_3376)
);

INVxp67_ASAP7_75t_L g3377 ( 
.A(n_3342),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3287),
.Y(n_3378)
);

OAI22xp5_ASAP7_75t_L g3379 ( 
.A1(n_3301),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3329),
.Y(n_3380)
);

INVxp67_ASAP7_75t_SL g3381 ( 
.A(n_3349),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3338),
.B(n_264),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3295),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3294),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3313),
.Y(n_3385)
);

OAI21xp5_ASAP7_75t_SL g3386 ( 
.A1(n_3296),
.A2(n_266),
.B(n_267),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_3316),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3321),
.Y(n_3388)
);

INVx3_ASAP7_75t_L g3389 ( 
.A(n_3340),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3297),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3300),
.Y(n_3391)
);

AND2x4_ASAP7_75t_L g3392 ( 
.A(n_3344),
.B(n_533),
.Y(n_3392)
);

INVxp67_ASAP7_75t_SL g3393 ( 
.A(n_3308),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3304),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3336),
.Y(n_3395)
);

BUFx6f_ASAP7_75t_L g3396 ( 
.A(n_3323),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3324),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3328),
.Y(n_3398)
);

HB1xp67_ASAP7_75t_L g3399 ( 
.A(n_3302),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3327),
.B(n_535),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3298),
.B(n_270),
.Y(n_3401)
);

AND2x4_ASAP7_75t_L g3402 ( 
.A(n_3317),
.B(n_536),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3330),
.Y(n_3403)
);

CKINVDCx5p33_ASAP7_75t_R g3404 ( 
.A(n_3346),
.Y(n_3404)
);

AND2x4_ASAP7_75t_L g3405 ( 
.A(n_3310),
.B(n_537),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3315),
.B(n_272),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3311),
.Y(n_3407)
);

OR2x2_ASAP7_75t_L g3408 ( 
.A(n_3314),
.B(n_272),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3305),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3320),
.B(n_3289),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3291),
.B(n_3322),
.Y(n_3411)
);

BUFx2_ASAP7_75t_L g3412 ( 
.A(n_3312),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3307),
.B(n_538),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3335),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3343),
.Y(n_3415)
);

AND2x4_ASAP7_75t_L g3416 ( 
.A(n_3337),
.B(n_539),
.Y(n_3416)
);

AND2x2_ASAP7_75t_L g3417 ( 
.A(n_3337),
.B(n_273),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3285),
.Y(n_3418)
);

BUFx2_ASAP7_75t_L g3419 ( 
.A(n_3337),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3394),
.B(n_540),
.Y(n_3420)
);

OAI221xp5_ASAP7_75t_L g3421 ( 
.A1(n_3412),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3395),
.B(n_541),
.Y(n_3422)
);

OA211x2_ASAP7_75t_L g3423 ( 
.A1(n_3368),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3355),
.B(n_3389),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3385),
.B(n_543),
.Y(n_3425)
);

OR2x2_ASAP7_75t_L g3426 ( 
.A(n_3372),
.B(n_3378),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3383),
.B(n_278),
.Y(n_3427)
);

AOI22xp33_ASAP7_75t_SL g3428 ( 
.A1(n_3393),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3391),
.B(n_544),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3352),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3384),
.B(n_281),
.Y(n_3431)
);

NOR2x1_ASAP7_75t_L g3432 ( 
.A(n_3376),
.B(n_3390),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3375),
.B(n_282),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3361),
.Y(n_3434)
);

NAND2x1_ASAP7_75t_SL g3435 ( 
.A(n_3392),
.B(n_282),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3370),
.Y(n_3436)
);

OR2x2_ASAP7_75t_L g3437 ( 
.A(n_3388),
.B(n_283),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3364),
.Y(n_3438)
);

INVxp67_ASAP7_75t_SL g3439 ( 
.A(n_3362),
.Y(n_3439)
);

BUFx2_ASAP7_75t_SL g3440 ( 
.A(n_3396),
.Y(n_3440)
);

OR2x2_ASAP7_75t_L g3441 ( 
.A(n_3380),
.B(n_284),
.Y(n_3441)
);

NOR2xp67_ASAP7_75t_L g3442 ( 
.A(n_3377),
.B(n_285),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3418),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3359),
.B(n_546),
.Y(n_3444)
);

AND2x4_ASAP7_75t_L g3445 ( 
.A(n_3356),
.B(n_286),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3369),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3363),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3354),
.B(n_549),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_3399),
.B(n_287),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_3357),
.B(n_287),
.Y(n_3450)
);

HB1xp67_ASAP7_75t_SL g3451 ( 
.A(n_3367),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3398),
.B(n_550),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3416),
.Y(n_3453)
);

NAND2x1p5_ASAP7_75t_L g3454 ( 
.A(n_3417),
.B(n_288),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_3407),
.B(n_289),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3409),
.B(n_290),
.Y(n_3456)
);

OR2x2_ASAP7_75t_L g3457 ( 
.A(n_3397),
.B(n_290),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3382),
.B(n_291),
.Y(n_3458)
);

OR2x2_ASAP7_75t_L g3459 ( 
.A(n_3403),
.B(n_291),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3374),
.Y(n_3460)
);

NAND3xp33_ASAP7_75t_L g3461 ( 
.A(n_3360),
.B(n_292),
.C(n_293),
.Y(n_3461)
);

OR2x2_ASAP7_75t_L g3462 ( 
.A(n_3414),
.B(n_292),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3415),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_3404),
.B(n_293),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_3411),
.A2(n_553),
.B1(n_554),
.B2(n_551),
.Y(n_3465)
);

AOI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3410),
.A2(n_553),
.B1(n_555),
.B2(n_551),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3379),
.Y(n_3467)
);

AOI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3402),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.C(n_297),
.Y(n_3468)
);

OR2x2_ASAP7_75t_L g3469 ( 
.A(n_3408),
.B(n_295),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3400),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3413),
.Y(n_3471)
);

OR2x2_ASAP7_75t_L g3472 ( 
.A(n_3401),
.B(n_298),
.Y(n_3472)
);

INVxp67_ASAP7_75t_L g3473 ( 
.A(n_3406),
.Y(n_3473)
);

OR2x2_ASAP7_75t_L g3474 ( 
.A(n_3365),
.B(n_298),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3405),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3358),
.B(n_556),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3353),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3419),
.Y(n_3478)
);

INVx3_ASAP7_75t_L g3479 ( 
.A(n_3371),
.Y(n_3479)
);

HB1xp67_ASAP7_75t_L g3480 ( 
.A(n_3373),
.Y(n_3480)
);

OAI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3387),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_3481)
);

NOR3xp33_ASAP7_75t_L g3482 ( 
.A(n_3379),
.B(n_300),
.C(n_301),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3351),
.Y(n_3483)
);

AND2x4_ASAP7_75t_L g3484 ( 
.A(n_3366),
.B(n_302),
.Y(n_3484)
);

OR2x2_ASAP7_75t_L g3485 ( 
.A(n_3381),
.B(n_303),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3351),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3351),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3419),
.B(n_304),
.Y(n_3488)
);

OR2x6_ASAP7_75t_L g3489 ( 
.A(n_3366),
.B(n_557),
.Y(n_3489)
);

OR2x2_ASAP7_75t_L g3490 ( 
.A(n_3381),
.B(n_304),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3351),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3419),
.B(n_304),
.Y(n_3492)
);

CKINVDCx16_ASAP7_75t_R g3493 ( 
.A(n_3396),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3381),
.B(n_558),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3419),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3419),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3351),
.Y(n_3497)
);

OAI21xp5_ASAP7_75t_SL g3498 ( 
.A1(n_3386),
.A2(n_305),
.B(n_306),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3351),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3381),
.B(n_558),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3419),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3381),
.B(n_559),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3351),
.Y(n_3503)
);

OR2x2_ASAP7_75t_L g3504 ( 
.A(n_3381),
.B(n_307),
.Y(n_3504)
);

OR2x2_ASAP7_75t_L g3505 ( 
.A(n_3381),
.B(n_308),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3381),
.B(n_560),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3419),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_3381),
.B(n_309),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3366),
.B(n_309),
.Y(n_3509)
);

NAND3xp33_ASAP7_75t_SL g3510 ( 
.A(n_3498),
.B(n_318),
.C(n_310),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3478),
.Y(n_3511)
);

AOI33xp33_ASAP7_75t_L g3512 ( 
.A1(n_3428),
.A2(n_313),
.A3(n_315),
.B1(n_311),
.B2(n_312),
.B3(n_314),
.Y(n_3512)
);

NAND3xp33_ASAP7_75t_L g3513 ( 
.A(n_3468),
.B(n_312),
.C(n_313),
.Y(n_3513)
);

AND2x2_ASAP7_75t_SL g3514 ( 
.A(n_3493),
.B(n_313),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3426),
.B(n_314),
.Y(n_3515)
);

NAND2x1p5_ASAP7_75t_SL g3516 ( 
.A(n_3432),
.B(n_3424),
.Y(n_3516)
);

AOI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3482),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_3517)
);

AND2x4_ASAP7_75t_L g3518 ( 
.A(n_3479),
.B(n_316),
.Y(n_3518)
);

OR2x2_ASAP7_75t_L g3519 ( 
.A(n_3463),
.B(n_317),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3495),
.B(n_319),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3496),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3501),
.B(n_320),
.Y(n_3522)
);

AOI222xp33_ASAP7_75t_L g3523 ( 
.A1(n_3461),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C1(n_562),
.C2(n_561),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3507),
.B(n_322),
.Y(n_3524)
);

BUFx2_ASAP7_75t_L g3525 ( 
.A(n_3439),
.Y(n_3525)
);

AOI33xp33_ASAP7_75t_L g3526 ( 
.A1(n_3481),
.A2(n_3467),
.A3(n_3471),
.B1(n_3470),
.B2(n_3465),
.B3(n_3466),
.Y(n_3526)
);

HB1xp67_ASAP7_75t_L g3527 ( 
.A(n_3480),
.Y(n_3527)
);

INVx4_ASAP7_75t_L g3528 ( 
.A(n_3489),
.Y(n_3528)
);

AOI221xp5_ASAP7_75t_L g3529 ( 
.A1(n_3421),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.C(n_568),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3453),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_3440),
.B(n_569),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3451),
.Y(n_3532)
);

AOI22xp33_ASAP7_75t_L g3533 ( 
.A1(n_3477),
.A2(n_573),
.B1(n_570),
.B2(n_572),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3460),
.B(n_574),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3430),
.Y(n_3535)
);

INVxp67_ASAP7_75t_L g3536 ( 
.A(n_3442),
.Y(n_3536)
);

OR2x2_ASAP7_75t_SL g3537 ( 
.A(n_3485),
.B(n_576),
.Y(n_3537)
);

OAI221xp5_ASAP7_75t_L g3538 ( 
.A1(n_3474),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.C(n_580),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3447),
.B(n_580),
.Y(n_3539)
);

AOI22xp33_ASAP7_75t_L g3540 ( 
.A1(n_3473),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3476),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_3541)
);

AOI31xp33_ASAP7_75t_L g3542 ( 
.A1(n_3454),
.A2(n_589),
.A3(n_587),
.B(n_588),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3434),
.B(n_588),
.Y(n_3543)
);

NOR2x1_ASAP7_75t_L g3544 ( 
.A(n_3437),
.B(n_590),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3446),
.B(n_590),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3436),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_3438),
.B(n_591),
.Y(n_3547)
);

OAI221xp5_ASAP7_75t_SL g3548 ( 
.A1(n_3489),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.C(n_595),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3475),
.B(n_593),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3429),
.B(n_594),
.Y(n_3550)
);

INVx1_ASAP7_75t_SL g3551 ( 
.A(n_3435),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_L g3552 ( 
.A(n_3457),
.B(n_596),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3483),
.Y(n_3553)
);

OAI222xp33_ASAP7_75t_L g3554 ( 
.A1(n_3469),
.A2(n_598),
.B1(n_601),
.B2(n_603),
.C1(n_597),
.C2(n_600),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3431),
.B(n_596),
.Y(n_3555)
);

AOI22xp33_ASAP7_75t_L g3556 ( 
.A1(n_3464),
.A2(n_604),
.B1(n_601),
.B2(n_603),
.Y(n_3556)
);

NAND3xp33_ASAP7_75t_L g3557 ( 
.A(n_3422),
.B(n_604),
.C(n_605),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3486),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3487),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3491),
.Y(n_3560)
);

INVx2_ASAP7_75t_SL g3561 ( 
.A(n_3484),
.Y(n_3561)
);

BUFx2_ASAP7_75t_L g3562 ( 
.A(n_3509),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3497),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3443),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3449),
.B(n_610),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3499),
.Y(n_3566)
);

AOI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_3420),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3488),
.B(n_3492),
.Y(n_3568)
);

OR2x2_ASAP7_75t_L g3569 ( 
.A(n_3455),
.B(n_614),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3503),
.Y(n_3570)
);

OAI33xp33_ASAP7_75t_L g3571 ( 
.A1(n_3441),
.A2(n_618),
.A3(n_620),
.B1(n_615),
.B2(n_617),
.B3(n_619),
.Y(n_3571)
);

NOR2x1_ASAP7_75t_L g3572 ( 
.A(n_3490),
.B(n_615),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3452),
.B(n_621),
.Y(n_3573)
);

AND2x4_ASAP7_75t_L g3574 ( 
.A(n_3433),
.B(n_622),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3504),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3459),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3532),
.B(n_3456),
.Y(n_3577)
);

BUFx3_ASAP7_75t_L g3578 ( 
.A(n_3562),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3528),
.B(n_3462),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3561),
.Y(n_3580)
);

BUFx2_ASAP7_75t_L g3581 ( 
.A(n_3536),
.Y(n_3581)
);

OR2x4_ASAP7_75t_L g3582 ( 
.A(n_3510),
.B(n_3472),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3525),
.B(n_3505),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3530),
.B(n_3450),
.Y(n_3584)
);

INVx1_ASAP7_75t_SL g3585 ( 
.A(n_3514),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3551),
.B(n_3494),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3527),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3568),
.B(n_3500),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3576),
.B(n_3502),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3575),
.B(n_3508),
.Y(n_3590)
);

AND2x4_ASAP7_75t_SL g3591 ( 
.A(n_3518),
.B(n_3445),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3526),
.B(n_3506),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3515),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_3511),
.B(n_3458),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_3521),
.B(n_3427),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3543),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3552),
.B(n_3425),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3544),
.B(n_3448),
.Y(n_3598)
);

OR2x2_ASAP7_75t_L g3599 ( 
.A(n_3516),
.B(n_3444),
.Y(n_3599)
);

OAI211xp5_ASAP7_75t_L g3600 ( 
.A1(n_3523),
.A2(n_3423),
.B(n_631),
.C(n_639),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3547),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3545),
.B(n_623),
.Y(n_3602)
);

NOR2xp67_ASAP7_75t_L g3603 ( 
.A(n_3519),
.B(n_627),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3534),
.B(n_628),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3537),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3572),
.B(n_632),
.Y(n_3606)
);

AND3x1_ASAP7_75t_L g3607 ( 
.A(n_3512),
.B(n_633),
.C(n_634),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_SL g3608 ( 
.A(n_3557),
.B(n_634),
.Y(n_3608)
);

OAI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3513),
.A2(n_635),
.B(n_636),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3520),
.B(n_3522),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3524),
.B(n_3549),
.Y(n_3611)
);

INVxp67_ASAP7_75t_L g3612 ( 
.A(n_3531),
.Y(n_3612)
);

NAND4xp25_ASAP7_75t_L g3613 ( 
.A(n_3529),
.B(n_639),
.C(n_637),
.D(n_638),
.Y(n_3613)
);

OR2x2_ASAP7_75t_L g3614 ( 
.A(n_3564),
.B(n_1215),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3539),
.B(n_641),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_3574),
.B(n_1217),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3535),
.Y(n_3617)
);

AOI322xp5_ASAP7_75t_L g3618 ( 
.A1(n_3517),
.A2(n_648),
.A3(n_647),
.B1(n_645),
.B2(n_643),
.C1(n_644),
.C2(n_646),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3605),
.B(n_3542),
.Y(n_3619)
);

OAI33xp33_ASAP7_75t_L g3620 ( 
.A1(n_3592),
.A2(n_3558),
.A3(n_3546),
.B1(n_3560),
.B2(n_3559),
.B3(n_3553),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3578),
.B(n_3563),
.Y(n_3621)
);

OR2x2_ASAP7_75t_L g3622 ( 
.A(n_3583),
.B(n_3569),
.Y(n_3622)
);

OR2x2_ASAP7_75t_L g3623 ( 
.A(n_3581),
.B(n_3565),
.Y(n_3623)
);

AND3x2_ASAP7_75t_L g3624 ( 
.A(n_3612),
.B(n_3555),
.C(n_3573),
.Y(n_3624)
);

OR2x2_ASAP7_75t_L g3625 ( 
.A(n_3586),
.B(n_3566),
.Y(n_3625)
);

OR2x2_ASAP7_75t_L g3626 ( 
.A(n_3590),
.B(n_3570),
.Y(n_3626)
);

INVx1_ASAP7_75t_SL g3627 ( 
.A(n_3591),
.Y(n_3627)
);

AND2x2_ASAP7_75t_L g3628 ( 
.A(n_3577),
.B(n_3550),
.Y(n_3628)
);

OR2x2_ASAP7_75t_L g3629 ( 
.A(n_3580),
.B(n_3548),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3610),
.B(n_3541),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3611),
.B(n_3567),
.Y(n_3631)
);

OAI22xp5_ASAP7_75t_L g3632 ( 
.A1(n_3582),
.A2(n_3533),
.B1(n_3538),
.B2(n_3540),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3584),
.B(n_3556),
.Y(n_3633)
);

OR2x2_ASAP7_75t_L g3634 ( 
.A(n_3588),
.B(n_3554),
.Y(n_3634)
);

OR2x2_ASAP7_75t_L g3635 ( 
.A(n_3593),
.B(n_645),
.Y(n_3635)
);

NAND2x1p5_ASAP7_75t_L g3636 ( 
.A(n_3579),
.B(n_3571),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3587),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3594),
.B(n_649),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3614),
.Y(n_3639)
);

OAI211xp5_ASAP7_75t_L g3640 ( 
.A1(n_3600),
.A2(n_3609),
.B(n_3599),
.C(n_3618),
.Y(n_3640)
);

HB1xp67_ASAP7_75t_L g3641 ( 
.A(n_3603),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3596),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3601),
.Y(n_3643)
);

AND2x4_ASAP7_75t_L g3644 ( 
.A(n_3595),
.B(n_650),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3617),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3598),
.B(n_1213),
.Y(n_3646)
);

OR2x6_ASAP7_75t_L g3647 ( 
.A(n_3606),
.B(n_651),
.Y(n_3647)
);

OR2x2_ASAP7_75t_L g3648 ( 
.A(n_3589),
.B(n_654),
.Y(n_3648)
);

NOR2x1_ASAP7_75t_L g3649 ( 
.A(n_3608),
.B(n_654),
.Y(n_3649)
);

AOI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3607),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3602),
.B(n_656),
.Y(n_3651)
);

INVx2_ASAP7_75t_SL g3652 ( 
.A(n_3616),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3597),
.B(n_657),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3604),
.B(n_659),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3615),
.Y(n_3655)
);

NAND2x1p5_ASAP7_75t_L g3656 ( 
.A(n_3613),
.B(n_660),
.Y(n_3656)
);

INVx1_ASAP7_75t_SL g3657 ( 
.A(n_3585),
.Y(n_3657)
);

NAND4xp25_ASAP7_75t_SL g3658 ( 
.A(n_3640),
.B(n_662),
.C(n_660),
.D(n_661),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3629),
.B(n_664),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3652),
.B(n_3627),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3622),
.Y(n_3661)
);

OAI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3632),
.A2(n_668),
.B(n_669),
.Y(n_3662)
);

OAI22xp33_ASAP7_75t_L g3663 ( 
.A1(n_3650),
.A2(n_673),
.B1(n_670),
.B2(n_672),
.Y(n_3663)
);

INVxp67_ASAP7_75t_L g3664 ( 
.A(n_3619),
.Y(n_3664)
);

OAI21xp33_ASAP7_75t_SL g3665 ( 
.A1(n_3634),
.A2(n_675),
.B(n_676),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3626),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3635),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3624),
.B(n_678),
.Y(n_3668)
);

OR2x2_ASAP7_75t_L g3669 ( 
.A(n_3623),
.B(n_3636),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3630),
.B(n_679),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3631),
.B(n_680),
.Y(n_3671)
);

OAI32xp33_ASAP7_75t_L g3672 ( 
.A1(n_3656),
.A2(n_684),
.A3(n_682),
.B1(n_683),
.B2(n_686),
.Y(n_3672)
);

HB1xp67_ASAP7_75t_L g3673 ( 
.A(n_3647),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3633),
.B(n_3628),
.Y(n_3674)
);

OR2x2_ASAP7_75t_L g3675 ( 
.A(n_3625),
.B(n_683),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3638),
.Y(n_3676)
);

OAI221xp5_ASAP7_75t_L g3677 ( 
.A1(n_3649),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.C(n_690),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3639),
.Y(n_3678)
);

OAI21xp5_ASAP7_75t_SL g3679 ( 
.A1(n_3642),
.A2(n_3643),
.B(n_3646),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3644),
.Y(n_3680)
);

OAI221xp5_ASAP7_75t_L g3681 ( 
.A1(n_3621),
.A2(n_692),
.B1(n_690),
.B2(n_691),
.C(n_693),
.Y(n_3681)
);

AOI221xp5_ASAP7_75t_L g3682 ( 
.A1(n_3620),
.A2(n_694),
.B1(n_691),
.B2(n_693),
.C(n_695),
.Y(n_3682)
);

AOI22xp5_ASAP7_75t_L g3683 ( 
.A1(n_3655),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.Y(n_3683)
);

HB1xp67_ASAP7_75t_L g3684 ( 
.A(n_3648),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3637),
.Y(n_3685)
);

OR2x2_ASAP7_75t_L g3686 ( 
.A(n_3653),
.B(n_701),
.Y(n_3686)
);

AOI22xp5_ASAP7_75t_L g3687 ( 
.A1(n_3645),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3654),
.B(n_706),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3651),
.Y(n_3689)
);

INVx1_ASAP7_75t_SL g3690 ( 
.A(n_3657),
.Y(n_3690)
);

HB1xp67_ASAP7_75t_L g3691 ( 
.A(n_3641),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3641),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3641),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3641),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3673),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3665),
.B(n_710),
.Y(n_3696)
);

AOI222xp33_ASAP7_75t_L g3697 ( 
.A1(n_3682),
.A2(n_728),
.B1(n_716),
.B2(n_736),
.C1(n_722),
.C2(n_711),
.Y(n_3697)
);

OAI21xp33_ASAP7_75t_L g3698 ( 
.A1(n_3660),
.A2(n_713),
.B(n_714),
.Y(n_3698)
);

AOI222xp33_ASAP7_75t_L g3699 ( 
.A1(n_3662),
.A2(n_3668),
.B1(n_3664),
.B2(n_3694),
.C1(n_3693),
.C2(n_3692),
.Y(n_3699)
);

OAI21xp33_ASAP7_75t_L g3700 ( 
.A1(n_3674),
.A2(n_719),
.B(n_720),
.Y(n_3700)
);

AOI221xp5_ASAP7_75t_L g3701 ( 
.A1(n_3679),
.A2(n_736),
.B1(n_739),
.B2(n_727),
.C(n_721),
.Y(n_3701)
);

OR2x2_ASAP7_75t_L g3702 ( 
.A(n_3659),
.B(n_721),
.Y(n_3702)
);

NAND4xp25_ASAP7_75t_L g3703 ( 
.A(n_3661),
.B(n_725),
.C(n_723),
.D(n_724),
.Y(n_3703)
);

AOI21xp33_ASAP7_75t_SL g3704 ( 
.A1(n_3677),
.A2(n_3666),
.B(n_3667),
.Y(n_3704)
);

AOI32xp33_ASAP7_75t_L g3705 ( 
.A1(n_3663),
.A2(n_729),
.A3(n_726),
.B1(n_727),
.B2(n_730),
.Y(n_3705)
);

OR2x2_ASAP7_75t_L g3706 ( 
.A(n_3670),
.B(n_732),
.Y(n_3706)
);

HB1xp67_ASAP7_75t_L g3707 ( 
.A(n_3684),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3672),
.A2(n_737),
.B(n_738),
.Y(n_3708)
);

INVx2_ASAP7_75t_SL g3709 ( 
.A(n_3680),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3689),
.B(n_740),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3676),
.B(n_744),
.Y(n_3711)
);

A2O1A1O1Ixp25_ASAP7_75t_L g3712 ( 
.A1(n_3681),
.A2(n_747),
.B(n_745),
.C(n_746),
.D(n_748),
.Y(n_3712)
);

OAI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3671),
.A2(n_751),
.B1(n_749),
.B2(n_750),
.Y(n_3713)
);

OAI221xp5_ASAP7_75t_L g3714 ( 
.A1(n_3678),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.C(n_755),
.Y(n_3714)
);

NOR2xp67_ASAP7_75t_L g3715 ( 
.A(n_3675),
.B(n_760),
.Y(n_3715)
);

OAI32xp33_ASAP7_75t_L g3716 ( 
.A1(n_3685),
.A2(n_762),
.A3(n_764),
.B1(n_761),
.B2(n_763),
.Y(n_3716)
);

AND2x4_ASAP7_75t_L g3717 ( 
.A(n_3686),
.B(n_3688),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3687),
.B(n_767),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3683),
.B(n_767),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3691),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3690),
.B(n_773),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3691),
.Y(n_3722)
);

AOI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3658),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_3723)
);

OAI322xp33_ASAP7_75t_L g3724 ( 
.A1(n_3669),
.A2(n_783),
.A3(n_782),
.B1(n_779),
.B2(n_777),
.C1(n_778),
.C2(n_780),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3691),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3691),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3691),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3691),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3691),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3691),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3691),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3691),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3691),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3691),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_3690),
.B(n_790),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3707),
.Y(n_3736)
);

O2A1O1Ixp33_ASAP7_75t_L g3737 ( 
.A1(n_3712),
.A2(n_798),
.B(n_796),
.C(n_797),
.Y(n_3737)
);

OR2x2_ASAP7_75t_L g3738 ( 
.A(n_3709),
.B(n_800),
.Y(n_3738)
);

AOI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_3695),
.A2(n_1202),
.B1(n_1203),
.B2(n_1201),
.Y(n_3739)
);

AOI21xp33_ASAP7_75t_L g3740 ( 
.A1(n_3699),
.A2(n_801),
.B(n_802),
.Y(n_3740)
);

AOI22xp5_ASAP7_75t_L g3741 ( 
.A1(n_3697),
.A2(n_1208),
.B1(n_1210),
.B2(n_1207),
.Y(n_3741)
);

NOR2x1_ASAP7_75t_L g3742 ( 
.A(n_3715),
.B(n_803),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3696),
.B(n_806),
.Y(n_3743)
);

O2A1O1Ixp5_ASAP7_75t_SL g3744 ( 
.A1(n_3720),
.A2(n_809),
.B(n_807),
.C(n_808),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3722),
.B(n_813),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3725),
.B(n_816),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3726),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3727),
.B(n_818),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3728),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3729),
.B(n_820),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3730),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3731),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3732),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3733),
.B(n_821),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3734),
.B(n_822),
.Y(n_3755)
);

INVx1_ASAP7_75t_SL g3756 ( 
.A(n_3702),
.Y(n_3756)
);

AOI221xp5_ASAP7_75t_L g3757 ( 
.A1(n_3704),
.A2(n_1202),
.B1(n_1204),
.B2(n_1200),
.C(n_1199),
.Y(n_3757)
);

NOR2x1_ASAP7_75t_L g3758 ( 
.A(n_3724),
.B(n_823),
.Y(n_3758)
);

INVx1_ASAP7_75t_SL g3759 ( 
.A(n_3706),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3723),
.B(n_825),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3721),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3735),
.B(n_826),
.Y(n_3762)
);

AOI22xp33_ASAP7_75t_L g3763 ( 
.A1(n_3717),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3698),
.B(n_833),
.Y(n_3764)
);

OAI221xp5_ASAP7_75t_L g3765 ( 
.A1(n_3740),
.A2(n_3701),
.B1(n_3705),
.B2(n_3708),
.C(n_3700),
.Y(n_3765)
);

AOI221xp5_ASAP7_75t_L g3766 ( 
.A1(n_3757),
.A2(n_3716),
.B1(n_3703),
.B2(n_3714),
.C(n_3713),
.Y(n_3766)
);

OAI221xp5_ASAP7_75t_L g3767 ( 
.A1(n_3741),
.A2(n_3711),
.B1(n_3710),
.B2(n_3718),
.C(n_3719),
.Y(n_3767)
);

NAND3xp33_ASAP7_75t_L g3768 ( 
.A(n_3736),
.B(n_3758),
.C(n_3742),
.Y(n_3768)
);

AOI221xp5_ASAP7_75t_L g3769 ( 
.A1(n_3747),
.A2(n_3752),
.B1(n_3753),
.B2(n_3751),
.C(n_3749),
.Y(n_3769)
);

NOR4xp25_ASAP7_75t_L g3770 ( 
.A(n_3756),
.B(n_844),
.C(n_842),
.D(n_843),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3738),
.Y(n_3771)
);

NOR4xp25_ASAP7_75t_L g3772 ( 
.A(n_3759),
.B(n_849),
.C(n_846),
.D(n_848),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3743),
.A2(n_858),
.B(n_859),
.Y(n_3773)
);

OAI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3745),
.A2(n_860),
.B(n_861),
.Y(n_3774)
);

AOI222xp33_ASAP7_75t_L g3775 ( 
.A1(n_3761),
.A2(n_866),
.B1(n_868),
.B2(n_862),
.C1(n_863),
.C2(n_867),
.Y(n_3775)
);

AOI222xp33_ASAP7_75t_L g3776 ( 
.A1(n_3746),
.A2(n_3754),
.B1(n_3748),
.B2(n_3755),
.C1(n_3750),
.C2(n_3760),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3764),
.B(n_878),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3762),
.A2(n_879),
.B(n_880),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_SL g3779 ( 
.A(n_3739),
.B(n_881),
.Y(n_3779)
);

AOI322xp5_ASAP7_75t_L g3780 ( 
.A1(n_3763),
.A2(n_3744),
.A3(n_1192),
.B1(n_886),
.B2(n_884),
.C1(n_885),
.C2(n_883),
.Y(n_3780)
);

O2A1O1Ixp33_ASAP7_75t_SL g3781 ( 
.A1(n_3737),
.A2(n_889),
.B(n_887),
.C(n_888),
.Y(n_3781)
);

OAI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3737),
.A2(n_891),
.B(n_892),
.Y(n_3782)
);

OAI221xp5_ASAP7_75t_L g3783 ( 
.A1(n_3782),
.A2(n_907),
.B1(n_905),
.B2(n_906),
.C(n_908),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_3781),
.A2(n_910),
.B(n_911),
.Y(n_3784)
);

OAI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_3768),
.A2(n_918),
.B1(n_916),
.B2(n_917),
.Y(n_3785)
);

OAI221xp5_ASAP7_75t_L g3786 ( 
.A1(n_3766),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.C(n_923),
.Y(n_3786)
);

OAI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3765),
.A2(n_929),
.B1(n_926),
.B2(n_928),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_SL g3788 ( 
.A(n_3770),
.B(n_3772),
.Y(n_3788)
);

OAI211xp5_ASAP7_75t_SL g3789 ( 
.A1(n_3776),
.A2(n_935),
.B(n_932),
.C(n_934),
.Y(n_3789)
);

AOI211xp5_ASAP7_75t_SL g3790 ( 
.A1(n_3767),
.A2(n_943),
.B(n_936),
.C(n_939),
.Y(n_3790)
);

INVx3_ASAP7_75t_L g3791 ( 
.A(n_3771),
.Y(n_3791)
);

OAI221xp5_ASAP7_75t_L g3792 ( 
.A1(n_3769),
.A2(n_947),
.B1(n_945),
.B2(n_946),
.C(n_948),
.Y(n_3792)
);

OAI211xp5_ASAP7_75t_L g3793 ( 
.A1(n_3780),
.A2(n_956),
.B(n_953),
.C(n_954),
.Y(n_3793)
);

AOI21xp33_ASAP7_75t_L g3794 ( 
.A1(n_3779),
.A2(n_970),
.B(n_968),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3788),
.A2(n_3773),
.B(n_3778),
.Y(n_3795)
);

O2A1O1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3789),
.A2(n_3774),
.B(n_3775),
.C(n_3777),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3791),
.Y(n_3797)
);

AOI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3784),
.A2(n_972),
.B(n_973),
.Y(n_3798)
);

XOR2x2_ASAP7_75t_L g3799 ( 
.A(n_3790),
.B(n_974),
.Y(n_3799)
);

AOI22xp5_ASAP7_75t_L g3800 ( 
.A1(n_3793),
.A2(n_1187),
.B1(n_1189),
.B2(n_1186),
.Y(n_3800)
);

O2A1O1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_3785),
.A2(n_978),
.B(n_975),
.C(n_977),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_L g3802 ( 
.A1(n_3787),
.A2(n_1182),
.B(n_1181),
.Y(n_3802)
);

AOI211xp5_ASAP7_75t_SL g3803 ( 
.A1(n_3786),
.A2(n_3783),
.B(n_3794),
.C(n_3792),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3795),
.A2(n_3798),
.B(n_3796),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_SL g3805 ( 
.A1(n_3797),
.A2(n_992),
.B1(n_989),
.B2(n_991),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3799),
.Y(n_3806)
);

OAI22xp33_ASAP7_75t_SL g3807 ( 
.A1(n_3800),
.A2(n_1000),
.B1(n_998),
.B2(n_999),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3802),
.Y(n_3808)
);

NOR2x1_ASAP7_75t_L g3809 ( 
.A(n_3808),
.B(n_3801),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3806),
.B(n_3803),
.Y(n_3810)
);

AO22x2_ASAP7_75t_L g3811 ( 
.A1(n_3804),
.A2(n_1005),
.B1(n_1002),
.B2(n_1003),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3807),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3811),
.Y(n_3813)
);

INVxp67_ASAP7_75t_L g3814 ( 
.A(n_3809),
.Y(n_3814)
);

OR2x2_ASAP7_75t_L g3815 ( 
.A(n_3812),
.B(n_3805),
.Y(n_3815)
);

NAND4xp75_ASAP7_75t_L g3816 ( 
.A(n_3810),
.B(n_1008),
.C(n_1006),
.D(n_1007),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3813),
.Y(n_3817)
);

NOR4xp25_ASAP7_75t_L g3818 ( 
.A(n_3815),
.B(n_1013),
.C(n_1011),
.D(n_1012),
.Y(n_3818)
);

AND2x4_ASAP7_75t_L g3819 ( 
.A(n_3816),
.B(n_1015),
.Y(n_3819)
);

AOI222xp33_ASAP7_75t_L g3820 ( 
.A1(n_3814),
.A2(n_1018),
.B1(n_1020),
.B2(n_1016),
.C1(n_1017),
.C2(n_1019),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3817),
.A2(n_1021),
.B1(n_1018),
.B2(n_1019),
.Y(n_3821)
);

AND3x2_ASAP7_75t_L g3822 ( 
.A(n_3818),
.B(n_1022),
.C(n_1023),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3822),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3823),
.B(n_3819),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3824),
.Y(n_3825)
);

CKINVDCx20_ASAP7_75t_R g3826 ( 
.A(n_3825),
.Y(n_3826)
);

AOI22xp5_ASAP7_75t_L g3827 ( 
.A1(n_3826),
.A2(n_3820),
.B1(n_3821),
.B2(n_1026),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3827),
.A2(n_1190),
.B1(n_1028),
.B2(n_1025),
.Y(n_3828)
);

INVx2_ASAP7_75t_SL g3829 ( 
.A(n_3828),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_3829),
.A2(n_1030),
.B1(n_1027),
.B2(n_1029),
.Y(n_3830)
);

AO221x2_ASAP7_75t_L g3831 ( 
.A1(n_3830),
.A2(n_1033),
.B1(n_1031),
.B2(n_1032),
.C(n_1035),
.Y(n_3831)
);

AOI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_3831),
.A2(n_1036),
.B(n_1039),
.Y(n_3832)
);

AOI211xp5_ASAP7_75t_L g3833 ( 
.A1(n_3832),
.A2(n_1045),
.B(n_1041),
.C(n_1043),
.Y(n_3833)
);


endmodule