module fake_aes_1336_n_702 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_702);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_702;
wire n_117;
wire n_663;
wire n_513;
wire n_361;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_7), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_50), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_71), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_41), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_18), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_70), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_31), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_54), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_0), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_47), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_26), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_21), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_37), .Y(n_98) );
INVx4_ASAP7_75t_R g99 ( .A(n_67), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_9), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_69), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_22), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_33), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_30), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_56), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_75), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_32), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_53), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_5), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_24), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_40), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_5), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_11), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_44), .Y(n_124) );
NOR2xp67_ASAP7_75t_L g125 ( .A(n_23), .B(n_12), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_111), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_92), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_107), .B(n_38), .Y(n_136) );
NOR2xp33_ASAP7_75t_R g137 ( .A(n_86), .B(n_42), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_80), .B(n_1), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_110), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_107), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_124), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_120), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g144 ( .A1(n_100), .A2(n_4), .B1(n_6), .B2(n_8), .Y(n_144) );
OR2x2_ASAP7_75t_L g145 ( .A(n_123), .B(n_4), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_86), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_109), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_109), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_79), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_85), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_89), .A2(n_49), .B(n_76), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_87), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_110), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_103), .B(n_6), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_90), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_93), .Y(n_166) );
INVx6_ASAP7_75t_L g167 ( .A(n_99), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_123), .Y(n_168) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_93), .A2(n_48), .B(n_74), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_167), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_159), .B(n_81), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_159), .B(n_97), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_127), .B(n_126), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_159), .B(n_118), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_142), .Y(n_177) );
AND3x2_ASAP7_75t_L g178 ( .A(n_139), .B(n_91), .C(n_112), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_159), .B(n_88), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_139), .A2(n_121), .B1(n_117), .B2(n_105), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_145), .A2(n_108), .B1(n_115), .B2(n_113), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
NAND2xp33_ASAP7_75t_L g184 ( .A(n_136), .B(n_104), .Y(n_184) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_136), .B(n_104), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_146), .B(n_98), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_158), .B(n_98), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_158), .B(n_102), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_129), .B(n_125), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_130), .B(n_102), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_167), .B(n_106), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_127), .B(n_122), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_143), .B(n_122), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_130), .B(n_119), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_132), .B(n_119), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_167), .B(n_116), .Y(n_199) );
BUFx10_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
INVxp67_ASAP7_75t_SL g203 ( .A(n_168), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_133), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_136), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_150), .B(n_114), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_134), .B(n_101), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_134), .B(n_95), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_135), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_135), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_128), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_128), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_138), .A2(n_94), .B1(n_95), .B2(n_11), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_141), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_164), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_138), .B(n_94), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_151), .B(n_51), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_151), .B(n_36), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_128), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_141), .Y(n_221) );
BUFx10_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_165), .B(n_9), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_164), .B(n_52), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_164), .B(n_55), .Y(n_225) );
BUFx8_ASAP7_75t_SL g226 ( .A(n_162), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_145), .B(n_10), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_141), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_141), .B(n_35), .Y(n_229) );
NAND2xp33_ASAP7_75t_SL g230 ( .A(n_137), .B(n_10), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_147), .B(n_13), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_200), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_227), .B(n_169), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_184), .A2(n_156), .B(n_169), .Y(n_235) );
AOI21xp33_ASAP7_75t_L g236 ( .A1(n_203), .A2(n_156), .B(n_144), .Y(n_236) );
INVx5_ASAP7_75t_L g237 ( .A(n_222), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_222), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_194), .B(n_149), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_195), .B(n_149), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_179), .B(n_147), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_191), .B(n_136), .Y(n_244) );
INVxp67_ASAP7_75t_SL g245 ( .A(n_227), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_175), .A2(n_164), .B1(n_163), .B2(n_131), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_210), .B(n_136), .Y(n_248) );
NOR3xp33_ASAP7_75t_SL g249 ( .A(n_177), .B(n_15), .C(n_16), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_226), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_194), .A2(n_136), .B1(n_164), .B2(n_156), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_181), .A2(n_163), .B1(n_131), .B2(n_154), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_188), .B(n_163), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_182), .B(n_15), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_231), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_187), .B(n_156), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_231), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_182), .A2(n_163), .B1(n_131), .B2(n_154), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_171), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_174), .B(n_131), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_174), .B(n_140), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_218), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_180), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_205), .B(n_152), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_183), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_181), .A2(n_140), .B1(n_154), .B2(n_160), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_205), .B(n_152), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_193), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_196), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_176), .B(n_140), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_197), .A2(n_140), .B1(n_154), .B2(n_160), .Y(n_275) );
BUFx12f_ASAP7_75t_L g276 ( .A(n_190), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_214), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_221), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_176), .B(n_160), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_201), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_202), .B(n_160), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_204), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_228), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_190), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_209), .B(n_157), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_206), .B(n_160), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_178), .Y(n_288) );
NOR2xp67_ASAP7_75t_SL g289 ( .A(n_185), .B(n_160), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_186), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_190), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_172), .B(n_157), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_207), .B(n_16), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_230), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_197), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_217), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_207), .Y(n_297) );
HAxp5_ASAP7_75t_L g298 ( .A(n_285), .B(n_213), .CON(n_298), .SN(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_297), .B(n_238), .Y(n_299) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_235), .A2(n_217), .B(n_219), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_280), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_245), .A2(n_197), .B1(n_198), .B2(n_208), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_241), .A2(n_216), .B1(n_219), .B2(n_192), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_256), .A2(n_199), .B(n_229), .C(n_189), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_236), .A2(n_253), .B(n_247), .C(n_242), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_258), .A2(n_229), .B(n_170), .C(n_225), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_237), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_240), .A2(n_157), .B1(n_148), .B2(n_152), .C(n_153), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_238), .B(n_198), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_260), .A2(n_198), .B(n_224), .C(n_20), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_293), .B(n_198), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_237), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_280), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_283), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_290), .B(n_224), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_237), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_288), .B(n_224), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_237), .B(n_224), .Y(n_318) );
NOR2x1p5_ASAP7_75t_L g319 ( .A(n_250), .B(n_157), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_244), .A2(n_220), .B(n_212), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_264), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
OAI22xp5_ASAP7_75t_SL g325 ( .A1(n_285), .A2(n_157), .B1(n_153), .B2(n_152), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_248), .A2(n_220), .B(n_212), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_267), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_293), .B(n_157), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_291), .A2(n_153), .B1(n_152), .B2(n_148), .C(n_128), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_232), .B(n_153), .Y(n_331) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_233), .B(n_153), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_296), .A2(n_220), .B(n_212), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_291), .A2(n_153), .B1(n_152), .B2(n_148), .C(n_128), .Y(n_334) );
BUFx4_ASAP7_75t_SL g335 ( .A(n_250), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_257), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_257), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
OAI21xp33_ASAP7_75t_SL g339 ( .A1(n_270), .A2(n_17), .B(n_19), .Y(n_339) );
BUFx12f_ASAP7_75t_L g340 ( .A(n_276), .Y(n_340) );
BUFx12f_ASAP7_75t_L g341 ( .A(n_276), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_262), .B(n_148), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_272), .A2(n_25), .B(n_27), .C(n_28), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_294), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_294), .B(n_29), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_273), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_243), .A2(n_148), .B(n_128), .C(n_211), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_262), .Y(n_348) );
NOR2x1p5_ASAP7_75t_L g349 ( .A(n_234), .B(n_148), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_338), .B(n_296), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_299), .B(n_243), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_320), .A2(n_252), .B(n_259), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_311), .B(n_234), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_282), .B(n_292), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_322), .B(n_281), .Y(n_357) );
CKINVDCx10_ASAP7_75t_R g358 ( .A(n_335), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_333), .A2(n_279), .B(n_268), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_307), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_306), .A2(n_268), .B(n_271), .Y(n_361) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_300), .A2(n_234), .B(n_287), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_329), .A2(n_271), .B(n_286), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_329), .A2(n_286), .B(n_295), .C(n_254), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_347), .A2(n_261), .B(n_275), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_302), .A2(n_265), .B1(n_263), .B2(n_274), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_343), .A2(n_275), .B(n_284), .Y(n_369) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_312), .B(n_284), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_300), .A2(n_249), .B(n_278), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_304), .A2(n_278), .B(n_277), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_346), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_310), .A2(n_277), .B(n_266), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_303), .A2(n_315), .B(n_305), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_307), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_301), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_303), .A2(n_266), .B(n_251), .Y(n_379) );
AO32x2_ASAP7_75t_L g380 ( .A1(n_325), .A2(n_289), .A3(n_60), .B1(n_61), .B2(n_62), .Y(n_380) );
OAI21x1_ASAP7_75t_SL g381 ( .A1(n_302), .A2(n_251), .B(n_246), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_349), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_375), .A2(n_332), .B(n_319), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_371), .A2(n_344), .B1(n_345), .B2(n_325), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_358), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_339), .B1(n_298), .B2(n_317), .C(n_308), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_316), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_377), .Y(n_388) );
OA21x2_ASAP7_75t_L g389 ( .A1(n_376), .A2(n_330), .B(n_334), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_352), .Y(n_390) );
BUFx10_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_353), .B(n_309), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_352), .B(n_339), .Y(n_394) );
OR2x6_ASAP7_75t_L g395 ( .A(n_355), .B(n_301), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_358), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_374), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_375), .A2(n_342), .B(n_331), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_355), .B(n_321), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_351), .A2(n_336), .B1(n_318), .B2(n_313), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_373), .B(n_318), .C(n_348), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_378), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_350), .A2(n_337), .B(n_348), .C(n_321), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_362), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_341), .B1(n_337), .B2(n_348), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_350), .Y(n_409) );
CKINVDCx11_ASAP7_75t_R g410 ( .A(n_362), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_395), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_409), .B(n_372), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_397), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_397), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_390), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_402), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_402), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_403), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_403), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_394), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_409), .B(n_372), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_387), .B(n_364), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_388), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_398), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_399), .B(n_364), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_391), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_407), .B(n_371), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_399), .B(n_378), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_391), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_410), .B(n_382), .C(n_357), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_392), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_399), .B(n_355), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_395), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_383), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_427), .B(n_382), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_412), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_417), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_428), .A2(n_391), .B1(n_400), .B2(n_404), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_437), .A2(n_386), .B1(n_355), .B2(n_384), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_420), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_429), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_429), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_415), .A2(n_386), .B1(n_408), .B2(n_393), .C(n_368), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_424), .B(n_425), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_424), .B(n_363), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_428), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_363), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_444), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_425), .B(n_363), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_434), .B(n_385), .C(n_396), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_427), .B(n_404), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_434), .B(n_404), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_430), .B(n_395), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_422), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_433), .B(n_400), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_430), .B(n_395), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_416), .B(n_395), .Y(n_478) );
OR2x6_ASAP7_75t_L g479 ( .A(n_444), .B(n_381), .Y(n_479) );
OAI21xp33_ASAP7_75t_L g480 ( .A1(n_445), .A2(n_405), .B(n_406), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_411), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_416), .B(n_391), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_423), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_418), .B(n_380), .Y(n_486) );
NOR2xp33_ASAP7_75t_R g487 ( .A(n_433), .B(n_313), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_418), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_418), .B(n_380), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_426), .B(n_380), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_429), .A2(n_401), .B(n_383), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_436), .A2(n_401), .B1(n_389), .B2(n_367), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g495 ( .A1(n_439), .A2(n_366), .A3(n_246), .B1(n_239), .B2(n_380), .B3(n_381), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_464), .B(n_443), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_494), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_456), .A2(n_421), .B1(n_411), .B2(n_442), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_463), .B(n_426), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_472), .B(n_413), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_481), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_470), .B(n_431), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_472), .B(n_413), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_464), .B(n_443), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_466), .B(n_421), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_463), .B(n_439), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_487), .Y(n_509) );
OAI321xp33_ASAP7_75t_L g510 ( .A1(n_480), .A2(n_436), .A3(n_441), .B1(n_431), .B2(n_442), .C(n_443), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_471), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_449), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_481), .B(n_421), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_494), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_448), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_467), .B(n_432), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_471), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_467), .B(n_432), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_462), .A2(n_441), .B1(n_411), .B2(n_435), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_468), .B(n_438), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_469), .B(n_438), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_468), .B(n_411), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_447), .B(n_435), .Y(n_523) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_488), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_469), .B(n_435), .Y(n_525) );
AO21x1_ASAP7_75t_SL g526 ( .A1(n_448), .A2(n_435), .B(n_380), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_488), .Y(n_527) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_482), .B(n_389), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_488), .Y(n_529) );
NAND2x1_ASAP7_75t_L g530 ( .A(n_482), .B(n_370), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_451), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_451), .B(n_383), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_490), .B(n_380), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_490), .B(n_354), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_450), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_452), .B(n_354), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_482), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_452), .B(n_453), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_453), .B(n_367), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_455), .B(n_367), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_455), .B(n_367), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_475), .B(n_370), .C(n_379), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_474), .B(n_389), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
NOR3xp33_ASAP7_75t_SL g547 ( .A(n_493), .B(n_57), .C(n_63), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_478), .B(n_378), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_450), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_457), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_478), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_454), .B(n_389), .C(n_211), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_457), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_497), .B(n_491), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_539), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_539), .B(n_476), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_512), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_501), .B(n_504), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_497), .B(n_491), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_506), .B(n_476), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
OAI21xp33_ASAP7_75t_L g563 ( .A1(n_519), .A2(n_495), .B(n_483), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_506), .B(n_483), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_508), .B(n_459), .Y(n_565) );
NAND2xp33_ASAP7_75t_SL g566 ( .A(n_538), .B(n_459), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_525), .B(n_492), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_525), .B(n_492), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_505), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_515), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_516), .B(n_492), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_510), .B(n_461), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_511), .B(n_485), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_498), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_517), .B(n_477), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_465), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_500), .B(n_477), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_531), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_550), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_516), .B(n_492), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_509), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_553), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_514), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_501), .B(n_465), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_514), .Y(n_585) );
OR2x6_ASAP7_75t_L g586 ( .A(n_538), .B(n_479), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_504), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_502), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_540), .B(n_461), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_534), .B(n_473), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_549), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_507), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_503), .Y(n_593) );
AOI221x1_ASAP7_75t_L g594 ( .A1(n_544), .A2(n_460), .B1(n_458), .B2(n_473), .C(n_489), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_523), .B(n_489), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_507), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_532), .Y(n_597) );
INVx4_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_502), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_535), .B(n_486), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_513), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_536), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_535), .B(n_486), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_593), .A2(n_499), .B1(n_552), .B2(n_533), .C(n_545), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_566), .A2(n_530), .B(n_524), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_581), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_589), .Y(n_609) );
AOI321xp33_ASAP7_75t_L g610 ( .A1(n_572), .A2(n_563), .A3(n_557), .B1(n_587), .B2(n_568), .C(n_567), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_566), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_589), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_572), .A2(n_528), .B1(n_548), .B2(n_533), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_599), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_559), .B(n_513), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_592), .B(n_518), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_555), .B(n_537), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_588), .A2(n_547), .B(n_527), .C(n_522), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_567), .A2(n_528), .B1(n_526), .B2(n_548), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_561), .B(n_537), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_586), .A2(n_522), .B1(n_527), .B2(n_479), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_520), .B1(n_479), .B2(n_529), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_586), .A2(n_479), .B(n_520), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_576), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_565), .A2(n_541), .B1(n_543), .B2(n_542), .C(n_518), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_601), .B(n_521), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_599), .A2(n_543), .B(n_542), .Y(n_629) );
OA21x2_ASAP7_75t_SL g630 ( .A1(n_556), .A2(n_548), .B(n_521), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_586), .A2(n_529), .B(n_541), .Y(n_631) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_591), .B(n_546), .C(n_356), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_596), .A2(n_546), .B1(n_460), .B2(n_458), .C(n_324), .Y(n_634) );
AO21x1_ASAP7_75t_L g635 ( .A1(n_598), .A2(n_324), .B(n_458), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_573), .A2(n_460), .B(n_458), .C(n_68), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_564), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_584), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_598), .B(n_460), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_598), .B(n_356), .C(n_361), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_584), .Y(n_641) );
O2A1O1Ixp5_ASAP7_75t_L g642 ( .A1(n_597), .A2(n_460), .B(n_65), .C(n_72), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_608), .B(n_570), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_613), .A2(n_568), .B1(n_571), .B2(n_580), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_627), .B(n_554), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_615), .B(n_578), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_616), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_610), .B(n_571), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_632), .B(n_594), .C(n_602), .Y(n_649) );
AOI221x1_ASAP7_75t_L g650 ( .A1(n_607), .A2(n_562), .B1(n_579), .B2(n_569), .C(n_582), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_618), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_633), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_614), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_617), .B(n_554), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_641), .B(n_560), .Y(n_656) );
AOI31xp33_ASAP7_75t_L g657 ( .A1(n_625), .A2(n_590), .A3(n_580), .B(n_575), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_628), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_614), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_611), .B(n_585), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_609), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_611), .A2(n_577), .B1(n_595), .B2(n_604), .C(n_605), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_638), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_606), .A2(n_560), .B1(n_585), .B2(n_583), .Y(n_664) );
XOR2xp5_ASAP7_75t_L g665 ( .A(n_621), .B(n_600), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_661), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_657), .A2(n_630), .B1(n_624), .B2(n_631), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_664), .A2(n_631), .B1(n_620), .B2(n_629), .C(n_623), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_648), .A2(n_624), .B1(n_622), .B2(n_626), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_660), .A2(n_639), .B(n_635), .Y(n_670) );
O2A1O1Ixp5_ASAP7_75t_L g671 ( .A1(n_660), .A2(n_612), .B(n_642), .C(n_619), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_664), .B(n_583), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_658), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_650), .A2(n_639), .B(n_636), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_662), .A2(n_634), .B(n_640), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g676 ( .A1(n_649), .A2(n_574), .B(n_558), .C(n_603), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_659), .B(n_574), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_654), .B(n_558), .C(n_603), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_658), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_666), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_667), .A2(n_645), .B(n_643), .C(n_663), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g682 ( .A1(n_670), .A2(n_644), .B(n_665), .C(n_643), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_669), .B(n_646), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_667), .A2(n_646), .B1(n_647), .B2(n_653), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g685 ( .A1(n_671), .A2(n_652), .B(n_651), .C(n_656), .Y(n_685) );
NOR2xp33_ASAP7_75t_SL g686 ( .A(n_674), .B(n_655), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_677), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_681), .A2(n_668), .B1(n_676), .B2(n_675), .C(n_672), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_680), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_686), .B(n_678), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_682), .B(n_673), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_682), .A2(n_679), .B1(n_369), .B2(n_361), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_689), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_691), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_688), .B(n_684), .C(n_683), .Y(n_695) );
AND3x1_ASAP7_75t_L g696 ( .A(n_694), .B(n_692), .C(n_685), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_693), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_695), .B1(n_690), .B2(n_687), .Y(n_698) );
AO22x2_ASAP7_75t_L g699 ( .A1(n_698), .A2(n_696), .B1(n_73), .B2(n_77), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_699), .A2(n_313), .B1(n_321), .B2(n_301), .Y(n_700) );
AOI22x1_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_64), .B1(n_211), .B2(n_239), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_359), .B1(n_365), .B2(n_369), .C1(n_694), .C2(n_697), .Y(n_702) );
endmodule