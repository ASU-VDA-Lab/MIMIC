module fake_jpeg_27645_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_33),
.B1(n_21),
.B2(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_43),
.Y(n_68)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_69),
.B1(n_33),
.B2(n_31),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_34),
.B1(n_26),
.B2(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_72),
.B1(n_64),
.B2(n_42),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_35),
.B(n_31),
.Y(n_56)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_47),
.B1(n_18),
.B2(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_73),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_110),
.B(n_29),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_107),
.B1(n_30),
.B2(n_16),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_86),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_34),
.B1(n_26),
.B2(n_21),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_109),
.Y(n_118)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_94),
.B(n_97),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_16),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_23),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_21),
.B1(n_30),
.B2(n_35),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_30),
.B1(n_19),
.B2(n_29),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_23),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx5_ASAP7_75t_SL g144 ( 
.A(n_106),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_58),
.A2(n_56),
.B1(n_19),
.B2(n_29),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_23),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_38),
.A3(n_36),
.B1(n_25),
.B2(n_48),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

AO22x2_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_57),
.B1(n_36),
.B2(n_38),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_18),
.B(n_2),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_88),
.B1(n_108),
.B2(n_89),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_48),
.C(n_44),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_77),
.C(n_114),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_36),
.B1(n_48),
.B2(n_44),
.Y(n_129)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_44),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_105),
.B(n_109),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_18),
.B1(n_27),
.B2(n_15),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_19),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_18),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_112),
.B1(n_92),
.B2(n_86),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_153),
.B1(n_161),
.B2(n_143),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_91),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_158),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_178),
.B(n_119),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_152),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_93),
.B1(n_90),
.B2(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_84),
.B1(n_96),
.B2(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_159),
.B1(n_164),
.B2(n_168),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_16),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_81),
.B1(n_82),
.B2(n_110),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_81),
.B1(n_82),
.B2(n_79),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_33),
.A3(n_25),
.B1(n_27),
.B2(n_32),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_173),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_128),
.A2(n_106),
.B1(n_77),
.B2(n_113),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_166),
.Y(n_203)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_100),
.C(n_32),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_121),
.C(n_124),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_120),
.A2(n_27),
.B1(n_32),
.B2(n_25),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_27),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_170),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_159),
.B1(n_151),
.B2(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_14),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_176),
.B(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_121),
.B(n_145),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_137),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_181),
.B(n_7),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_196),
.B(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_136),
.B1(n_126),
.B2(n_144),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_200),
.B1(n_201),
.B2(n_205),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_190),
.B1(n_209),
.B2(n_183),
.Y(n_222)
);

OAI22x1_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_140),
.B1(n_121),
.B2(n_129),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_187),
.A2(n_9),
.B(n_10),
.C(n_185),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_126),
.B1(n_143),
.B2(n_133),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_202),
.B(n_204),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_133),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_148),
.B(n_169),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_166),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_143),
.B1(n_145),
.B2(n_144),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_18),
.B(n_124),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_146),
.A2(n_122),
.B(n_129),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_1),
.B(n_2),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_13),
.C(n_3),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_4),
.C(n_5),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_153),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_174),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_162),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

AOI22x1_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_161),
.B1(n_168),
.B2(n_177),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_227),
.B1(n_238),
.B2(n_186),
.Y(n_251)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_165),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_199),
.C(n_181),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_158),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_237),
.Y(n_243)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_218),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_189),
.B(n_149),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_207),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

NAND2x1_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_150),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_187),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_208),
.B1(n_209),
.B2(n_193),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_189),
.B(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_192),
.Y(n_234)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_8),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_8),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_182),
.B(n_9),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_260),
.Y(n_262)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_251),
.B1(n_259),
.B2(n_235),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_197),
.C(n_193),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_254),
.C(n_243),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_231),
.B(n_225),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_233),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_180),
.B1(n_200),
.B2(n_202),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_220),
.B1(n_228),
.B2(n_227),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_243),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_184),
.C(n_180),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_206),
.B1(n_201),
.B2(n_194),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_191),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_264),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_265),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_231),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_270),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_277),
.C(n_238),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_250),
.B1(n_258),
.B2(n_241),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_237),
.C(n_212),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.C(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_215),
.C(n_226),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_274),
.A2(n_278),
.B1(n_251),
.B2(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_195),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_236),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_269),
.C(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_287),
.C(n_291),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_252),
.B1(n_244),
.B2(n_247),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_241),
.B1(n_218),
.B2(n_234),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_253),
.C(n_238),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_224),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_238),
.C(n_258),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_204),
.C(n_211),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_263),
.C(n_268),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_268),
.B1(n_275),
.B2(n_264),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_299),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_270),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_300),
.C(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_274),
.B(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_281),
.C(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_234),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_286),
.C(n_293),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_294),
.C(n_296),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_298),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_296),
.C(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_295),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_314),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_320),
.B(n_315),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_323),
.B(n_306),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_192),
.C(n_9),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_9),
.C(n_10),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_10),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_10),
.Y(n_330)
);


endmodule