module real_jpeg_33652_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_690, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_690;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_620;
wire n_328;
wire n_366;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_0),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_0),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_0),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_1),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_76),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_1),
.A2(n_76),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_1),
.A2(n_76),
.B1(n_343),
.B2(n_347),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_2),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_2),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_2),
.A2(n_48),
.B1(n_361),
.B2(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_2),
.A2(n_361),
.B1(n_563),
.B2(n_564),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_2),
.A2(n_361),
.B1(n_643),
.B2(n_647),
.Y(n_642)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_4),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_4),
.A2(n_52),
.B1(n_194),
.B2(n_200),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_4),
.A2(n_52),
.B1(n_150),
.B2(n_240),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_4),
.A2(n_52),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_5),
.A2(n_122),
.B1(n_123),
.B2(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_5),
.A2(n_122),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_5),
.A2(n_122),
.B1(n_350),
.B2(n_353),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_5),
.A2(n_122),
.B1(n_480),
.B2(n_482),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_6),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_6),
.A2(n_159),
.B1(n_171),
.B2(n_176),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_159),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_7),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_8),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_8),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_8),
.A2(n_254),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_8),
.A2(n_254),
.B1(n_448),
.B2(n_452),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_8),
.A2(n_254),
.B1(n_542),
.B2(n_545),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_9),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_9),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_9),
.A2(n_313),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_9),
.A2(n_313),
.B1(n_509),
.B2(n_513),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_9),
.A2(n_313),
.B1(n_606),
.B2(n_620),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_10),
.A2(n_90),
.B1(n_264),
.B2(n_269),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_10),
.A2(n_90),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_10),
.A2(n_90),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_14),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_20),
.B(n_687),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_15),
.B(n_688),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_16),
.B(n_93),
.Y(n_408)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_16),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_16),
.B(n_98),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_16),
.B(n_534),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_16),
.A2(n_459),
.B1(n_571),
.B2(n_576),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_L g660 ( 
.A1(n_16),
.A2(n_221),
.B(n_623),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_17),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_205),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_204),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_186),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_24),
.B(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_164),
.C(n_165),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_26),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_26),
.B(n_210),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_82),
.C(n_128),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_28),
.A2(n_128),
.B1(n_168),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_28),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_46),
.B1(n_61),
.B2(n_73),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_29),
.A2(n_46),
.B1(n_61),
.B2(n_170),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_29),
.A2(n_61),
.B(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_29),
.A2(n_73),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_29),
.A2(n_61),
.B1(n_263),
.B2(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_29),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_29),
.B(n_370),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_29),
.A2(n_61),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_62),
.Y(n_61)
);

AOI22x1_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_35),
.B1(n_38),
.B2(n_42),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_31),
.A2(n_147),
.B1(n_150),
.B2(n_153),
.Y(n_146)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_33),
.Y(n_352)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_34),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_34),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_34),
.Y(n_589)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_40),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_41),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_41),
.Y(n_356)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_45),
.Y(n_531)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_49),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_50),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_50),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_51),
.Y(n_175)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_51),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_51),
.Y(n_579)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_60),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_61),
.Y(n_262)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_61),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_61),
.B(n_370),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_64),
.Y(n_527)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_81),
.Y(n_371)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_82),
.B(n_166),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_83),
.B(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_97),
.B1(n_109),
.B2(n_121),
.Y(n_83)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_88),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_96),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_96),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_96),
.Y(n_365)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_97),
.A2(n_109),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_98),
.B(n_121),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_98),
.B(n_252),
.Y(n_318)
);

AO22x1_ASAP7_75t_SL g359 ( 
.A1(n_98),
.A2(n_110),
.B1(n_312),
.B2(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_98),
.B(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_104),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_106),
.Y(n_393)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_110),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_110),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_110),
.B(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_114),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_114),
.Y(n_415)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_168),
.B1(n_169),
.B2(n_177),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_144),
.B(n_156),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_129),
.A2(n_144),
.B1(n_156),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_129),
.A2(n_144),
.B1(n_447),
.B2(n_455),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_129),
.B(n_447),
.Y(n_516)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_130),
.Y(n_630)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_131),
.B(n_146),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_249)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_134),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_137),
.Y(n_297)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_137),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_138),
.Y(n_423)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_138),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_138),
.Y(n_549)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_140),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_142),
.Y(n_613)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_144),
.B(n_616),
.Y(n_615)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_144),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_152),
.Y(n_567)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_158),
.Y(n_454)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_158),
.Y(n_515)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_163),
.Y(n_451)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_163),
.Y(n_604)
);

INVxp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_178),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_177),
.C(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_171),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_175),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_185),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_202),
.B2(n_203),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_194),
.A2(n_459),
.B(n_460),
.Y(n_458)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_199),
.Y(n_403)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_323),
.B(n_681),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_270),
.Y(n_207)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_208),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B(n_212),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_258),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_214),
.A2(n_258),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_218),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_250),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_219),
.A2(n_220),
.B(n_236),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_236),
.Y(n_219)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

AOI21x1_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_227),
.B(n_230),
.Y(n_220)
);

OAI22x1_ASAP7_75t_SL g293 ( 
.A1(n_221),
.A2(n_230),
.B1(n_294),
.B2(n_301),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_221),
.A2(n_421),
.B1(n_479),
.B2(n_485),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_221),
.A2(n_619),
.B(n_623),
.Y(n_618)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_222),
.B(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_222),
.A2(n_342),
.B1(n_417),
.B2(n_420),
.Y(n_416)
);

AO22x1_ASAP7_75t_SL g540 ( 
.A1(n_222),
.A2(n_541),
.B1(n_550),
.B2(n_551),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_222),
.A2(n_638),
.B1(n_640),
.B2(n_641),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_R g658 ( 
.A(n_222),
.B(n_541),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_224),
.Y(n_340)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_233),
.Y(n_622)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_235),
.Y(n_346)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_235),
.Y(n_481)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_235),
.Y(n_599)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_235),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_247),
.B2(n_248),
.Y(n_237)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_238),
.A2(n_239),
.B1(n_248),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_238),
.A2(n_248),
.B1(n_288),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_238),
.A2(n_248),
.B1(n_508),
.B2(n_562),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_239),
.Y(n_276)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_260),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_251),
.B(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_253),
.Y(n_362)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_261),
.Y(n_282)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_319),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_271),
.B(n_319),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.C(n_283),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_273),
.B(n_282),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_278),
.B(n_279),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_277),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_284),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_304),
.C(n_309),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_287),
.B(n_293),
.Y(n_426)
);

BUFx4f_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_294),
.A2(n_339),
.B(n_341),
.Y(n_338)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_300),
.Y(n_544)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_300),
.Y(n_611)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_301),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_303),
.Y(n_657)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_310),
.Y(n_332)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_318),
.Y(n_310)
);

INVx11_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_318),
.B(n_457),
.Y(n_456)
);

NAND2x1_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_496),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_435),
.B(n_492),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_326),
.B(n_678),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_378),
.B(n_381),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_327),
.B(n_378),
.Y(n_495)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_328),
.B(n_379),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.C(n_335),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_330),
.A2(n_331),
.B1(n_334),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_334),
.Y(n_434)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_336),
.B(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_357),
.B(n_377),
.Y(n_336)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_348),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_338),
.B(n_348),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_340),
.Y(n_624)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_356),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_366),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_366),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_358),
.A2(n_359),
.B1(n_367),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

OAI22x1_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_375),
.B2(n_376),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_368),
.A2(n_387),
.B(n_394),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_368),
.A2(n_394),
.B(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_376),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

NOR2x1_ASAP7_75t_R g626 ( 
.A(n_376),
.B(n_459),
.Y(n_626)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_432),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_382),
.B(n_432),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_426),
.C(n_427),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_383),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_395),
.C(n_398),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_385),
.A2(n_386),
.B1(n_395),
.B2(n_396),
.Y(n_444)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_416),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_400),
.B(n_416),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_404),
.B1(n_408),
.B2(n_409),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_408),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_419),
.Y(n_666)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_426),
.A2(n_428),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_426),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_441),
.C(n_468),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_437),
.A2(n_679),
.B(n_680),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_441),
.Y(n_679)
);

MAJx2_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.C(n_466),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_442),
.A2(n_443),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_467),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_456),
.C(n_461),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_461),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_447),
.Y(n_629)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_471),
.Y(n_470)
);

OAI211xp5_ASAP7_75t_L g519 ( 
.A1(n_459),
.A2(n_520),
.B(n_524),
.C(n_528),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_459),
.B(n_602),
.Y(n_601)
);

OAI21xp33_ASAP7_75t_SL g616 ( 
.A1(n_459),
.A2(n_510),
.B(n_601),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_459),
.B(n_630),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_459),
.B(n_663),
.Y(n_662)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_489),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_469),
.B(n_489),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.C(n_473),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_470),
.B(n_553),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_472),
.A2(n_473),
.B1(n_474),
.B2(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_472),
.Y(n_554)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.C(n_487),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_503),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_478),
.A2(n_487),
.B1(n_488),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_478),
.Y(n_504)
);

INVxp33_ASAP7_75t_SL g550 ( 
.A(n_479),
.Y(n_550)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_484),
.Y(n_649)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B(n_495),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_677),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_555),
.B(n_675),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_552),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_500),
.B(n_676),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_505),
.C(n_517),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_502),
.B(n_558),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_505),
.A2(n_506),
.B1(n_517),
.B2(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_507),
.A2(n_508),
.B(n_516),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_516),
.B(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_540),
.Y(n_517)
);

XOR2x1_ASAP7_75t_L g580 ( 
.A(n_518),
.B(n_540),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_532),
.Y(n_518)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_535),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_SL g623 ( 
.A(n_541),
.B(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_552),
.Y(n_676)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_556),
.A2(n_581),
.B(n_674),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_557),
.B(n_560),
.Y(n_556)
);

NOR2x1_ASAP7_75t_L g674 ( 
.A(n_557),
.B(n_560),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_SL g560 ( 
.A(n_561),
.B(n_568),
.C(n_580),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_569),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_562),
.A2(n_628),
.B1(n_629),
.B2(n_630),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

BUFx2_ASAP7_75t_SL g572 ( 
.A(n_573),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_580),
.B(n_634),
.Y(n_633)
);

OAI321xp33_ASAP7_75t_L g581 ( 
.A1(n_582),
.A2(n_631),
.A3(n_635),
.B1(n_672),
.B2(n_673),
.C(n_690),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_617),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_583),
.B(n_617),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_614),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_584),
.B(n_614),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_585),
.A2(n_595),
.B1(n_600),
.B2(n_605),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_590),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_606),
.B(n_612),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_613),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_625),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_626),
.C(n_627),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_619),
.Y(n_640)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

BUFx2_ASAP7_75t_SL g621 ( 
.A(n_622),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_626),
.B(n_627),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_633),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_632),
.B(n_633),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_636),
.A2(n_651),
.B(n_671),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_637),
.B(n_650),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_650),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_642),
.A2(n_655),
.B(n_658),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

BUFx2_ASAP7_75t_SL g645 ( 
.A(n_646),
.Y(n_645)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_652),
.A2(n_659),
.B(n_670),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_653),
.B(n_654),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_653),
.B(n_654),
.Y(n_670)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_660),
.B(n_661),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_662),
.B(n_667),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_665),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_668),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_669),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_682),
.A2(n_684),
.B(n_685),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_683),
.Y(n_682)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_686),
.Y(n_685)
);


endmodule