module real_aes_17986_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_917;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_397;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_0), .Y(n_190) );
AND2x4_ASAP7_75t_L g114 ( .A(n_1), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g918 ( .A(n_2), .Y(n_918) );
BUFx3_ASAP7_75t_L g274 ( .A(n_3), .Y(n_274) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_5), .B(n_237), .Y(n_236) );
BUFx2_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
OR2x2_ASAP7_75t_L g127 ( .A(n_6), .B(n_20), .Y(n_127) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_7), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_8), .B(n_163), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_9), .B(n_163), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_10), .B(n_175), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_11), .A2(n_84), .B1(n_159), .B2(n_163), .Y(n_162) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_12), .A2(n_37), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_13), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_14), .B(n_182), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_15), .Y(n_588) );
AO32x1_ASAP7_75t_L g150 ( .A1(n_16), .A2(n_151), .A3(n_154), .B1(n_165), .B2(n_169), .Y(n_150) );
AO32x2_ASAP7_75t_L g282 ( .A1(n_16), .A2(n_151), .A3(n_154), .B1(n_165), .B2(n_169), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_17), .B(n_574), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_18), .B(n_169), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_19), .Y(n_612) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_21), .A2(n_44), .B1(n_182), .B2(n_183), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_22), .A2(n_92), .B1(n_159), .B2(n_161), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_23), .B(n_207), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_24), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_25), .B(n_205), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_26), .A2(n_64), .B1(n_161), .B2(n_297), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_27), .A2(n_32), .B1(n_894), .B2(n_895), .Y(n_893) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_27), .Y(n_894) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_28), .B(n_163), .Y(n_603) );
INVx2_ASAP7_75t_L g123 ( .A(n_29), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_30), .B(n_164), .Y(n_622) );
BUFx3_ASAP7_75t_L g118 ( .A(n_31), .Y(n_118) );
INVx1_ASAP7_75t_L g889 ( .A(n_31), .Y(n_889) );
INVx1_ASAP7_75t_L g895 ( .A(n_32), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_33), .B(n_212), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g904 ( .A(n_34), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_35), .B(n_566), .Y(n_628) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_35), .Y(n_899) );
AOI22x1_ASAP7_75t_SL g133 ( .A1(n_36), .A2(n_71), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_36), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_38), .Y(n_137) );
AND2x2_ASAP7_75t_L g594 ( .A(n_39), .B(n_566), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_40), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_41), .B(n_191), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_42), .B(n_574), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_43), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_45), .B(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_46), .A2(n_79), .B1(n_191), .B2(n_205), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_47), .B(n_297), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_48), .A2(n_155), .B(n_188), .C(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_49), .A2(n_81), .B1(n_159), .B2(n_163), .Y(n_270) );
INVx1_ASAP7_75t_L g153 ( .A(n_50), .Y(n_153) );
AND2x4_ASAP7_75t_L g167 ( .A(n_51), .B(n_168), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_52), .A2(n_53), .B1(n_161), .B2(n_183), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_54), .B(n_169), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_55), .B(n_566), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_56), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g129 ( .A(n_57), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_58), .B(n_161), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_59), .B(n_159), .Y(n_235) );
INVx1_ASAP7_75t_L g168 ( .A(n_60), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_61), .B(n_169), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_62), .A2(n_188), .B(n_189), .C(n_192), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_63), .B(n_159), .C(n_240), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_65), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_66), .B(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_67), .B(n_169), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_68), .B(n_548), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_69), .Y(n_300) );
AND2x2_ASAP7_75t_L g195 ( .A(n_70), .B(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g135 ( .A(n_71), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_72), .B(n_164), .C(n_182), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_73), .A2(n_96), .B1(n_163), .B2(n_191), .Y(n_223) );
INVx2_ASAP7_75t_L g157 ( .A(n_74), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_75), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_76), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_77), .B(n_186), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_78), .B(n_163), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_80), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_82), .B(n_258), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_83), .A2(n_91), .B1(n_574), .B2(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_85), .B(n_163), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_86), .B(n_240), .Y(n_239) );
NAND2xp33_ASAP7_75t_SL g564 ( .A(n_87), .B(n_237), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_88), .B(n_254), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_89), .A2(n_103), .B1(n_161), .B2(n_183), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_90), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_93), .B(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_94), .A2(n_898), .B1(n_899), .B2(n_900), .Y(n_897) );
INVx1_ASAP7_75t_L g900 ( .A(n_94), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_95), .B(n_175), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_97), .B(n_237), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_98), .B(n_566), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_99), .B(n_186), .C(n_237), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_100), .B(n_548), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_101), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_102), .B(n_574), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_119), .B(n_917), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx12f_ASAP7_75t_L g921 ( .A(n_107), .Y(n_921) );
AND2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_112), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
NOR3x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .C(n_118), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g533 ( .A(n_117), .Y(n_533) );
INVx1_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
NOR2x1_ASAP7_75t_L g916 ( .A(n_118), .B(n_127), .Y(n_916) );
AO21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_128), .B(n_882), .Y(n_119) );
BUFx12f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_SL g121 ( .A(n_122), .B(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g884 ( .A(n_123), .B(n_885), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_123), .B(n_914), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x6_ASAP7_75t_SL g886 ( .A(n_126), .B(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
XNOR2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_140), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_136), .B1(n_137), .B2(n_138), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_137), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_139), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_531), .B1(n_532), .B2(n_534), .Y(n_140) );
XNOR2xp5_ASAP7_75t_L g892 ( .A(n_141), .B(n_893), .Y(n_892) );
NOR2x1p5_ASAP7_75t_L g141 ( .A(n_142), .B(n_451), .Y(n_141) );
NAND4xp75_ASAP7_75t_L g142 ( .A(n_143), .B(n_330), .C(n_383), .D(n_428), .Y(n_142) );
NOR2x1_ASAP7_75t_L g143 ( .A(n_144), .B(n_287), .Y(n_143) );
OAI21xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_215), .B(n_244), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_170), .Y(n_146) );
AND2x4_ASAP7_75t_L g419 ( .A(n_147), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_147), .B(n_293), .Y(n_447) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_148), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g412 ( .A(n_149), .Y(n_412) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_149), .Y(n_434) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_L g318 ( .A(n_150), .B(n_294), .Y(n_318) );
INVx1_ASAP7_75t_L g340 ( .A(n_150), .Y(n_340) );
AND2x2_ASAP7_75t_L g374 ( .A(n_150), .B(n_294), .Y(n_374) );
INVx4_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
INVx2_ASAP7_75t_SL g201 ( .A(n_151), .Y(n_201) );
BUFx3_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
INVx2_ASAP7_75t_L g249 ( .A(n_151), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_151), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_151), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_SL g554 ( .A(n_151), .B(n_242), .Y(n_554) );
INVx1_ASAP7_75t_SL g557 ( .A(n_151), .Y(n_557) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B1(n_162), .B2(n_164), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g251 ( .A1(n_155), .A2(n_252), .B(n_253), .C(n_255), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_155), .A2(n_547), .B(n_549), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_155), .A2(n_563), .B(n_564), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_155), .A2(n_572), .B(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_155), .A2(n_602), .B(n_603), .Y(n_601) );
BUFx4f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g240 ( .A(n_156), .Y(n_240) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx8_ASAP7_75t_L g164 ( .A(n_157), .Y(n_164) );
INVx1_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
INVx2_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx2_ASAP7_75t_SL g205 ( .A(n_159), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_159), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_160), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_160), .Y(n_163) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
INVx1_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
INVx1_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_160), .Y(n_237) );
INVx1_ASAP7_75t_L g254 ( .A(n_160), .Y(n_254) );
INVx3_ASAP7_75t_L g548 ( .A(n_160), .Y(n_548) );
INVx1_ASAP7_75t_L g575 ( .A(n_160), .Y(n_575) );
INVx2_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_161), .A2(n_548), .B1(n_592), .B2(n_593), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_161), .A2(n_622), .B(n_623), .Y(n_621) );
INVx2_ASAP7_75t_L g649 ( .A(n_161), .Y(n_649) );
INVx3_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_163), .A2(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g627 ( .A(n_163), .Y(n_627) );
INVx6_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_164), .A2(n_235), .B(n_236), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_164), .A2(n_213), .B1(n_270), .B2(n_271), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_164), .A2(n_605), .B(n_606), .Y(n_604) );
O2A1O1Ixp5_ASAP7_75t_L g611 ( .A1(n_164), .A2(n_253), .B(n_612), .C(n_613), .Y(n_611) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_165), .A2(n_203), .B(n_209), .Y(n_202) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_SL g224 ( .A(n_166), .Y(n_224) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
BUFx10_ASAP7_75t_L g242 ( .A(n_167), .Y(n_242) );
AO31x2_ASAP7_75t_L g294 ( .A1(n_167), .A2(n_219), .A3(n_295), .B(n_299), .Y(n_294) );
BUFx10_ASAP7_75t_L g584 ( .A(n_167), .Y(n_584) );
INVx2_ASAP7_75t_L g268 ( .A(n_169), .Y(n_268) );
INVxp33_ASAP7_75t_L g369 ( .A(n_170), .Y(n_369) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OR2x2_ASAP7_75t_L g481 ( .A(n_171), .B(n_318), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_198), .Y(n_171) );
OR2x2_ASAP7_75t_L g361 ( .A(n_172), .B(n_199), .Y(n_361) );
INVx1_ASAP7_75t_L g394 ( .A(n_172), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_172), .Y(n_398) );
AND2x2_ASAP7_75t_L g514 ( .A(n_172), .B(n_329), .Y(n_514) );
OR2x2_ASAP7_75t_L g520 ( .A(n_172), .B(n_340), .Y(n_520) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g279 ( .A(n_173), .Y(n_279) );
AOI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_178), .B(n_195), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp67_ASAP7_75t_SL g582 ( .A(n_175), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AO31x2_ASAP7_75t_L g646 ( .A1(n_176), .A2(n_584), .A3(n_647), .B(n_651), .Y(n_646) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g197 ( .A(n_177), .Y(n_197) );
INVx2_ASAP7_75t_L g232 ( .A(n_177), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_187), .B(n_194), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_180), .B(n_185), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_180) );
INVx2_ASAP7_75t_L g297 ( .A(n_182), .Y(n_297) );
INVx1_ASAP7_75t_L g260 ( .A(n_183), .Y(n_260) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_185), .A2(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_SL g222 ( .A(n_186), .Y(n_222) );
INVx1_ASAP7_75t_L g552 ( .A(n_188), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx2_ASAP7_75t_L g208 ( .A(n_192), .Y(n_208) );
INVx2_ASAP7_75t_L g590 ( .A(n_192), .Y(n_590) );
BUFx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g259 ( .A(n_193), .Y(n_259) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_197), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_197), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g414 ( .A(n_198), .B(n_364), .Y(n_414) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g280 ( .A(n_199), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g284 ( .A(n_199), .B(n_281), .Y(n_284) );
AND2x2_ASAP7_75t_L g291 ( .A(n_199), .B(n_282), .Y(n_291) );
INVx2_ASAP7_75t_L g315 ( .A(n_199), .Y(n_315) );
INVx1_ASAP7_75t_L g338 ( .A(n_199), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_199), .B(n_294), .Y(n_411) );
AND2x2_ASAP7_75t_L g420 ( .A(n_199), .B(n_278), .Y(n_420) );
INVxp67_ASAP7_75t_L g490 ( .A(n_199), .Y(n_490) );
BUFx2_ASAP7_75t_L g498 ( .A(n_199), .Y(n_498) );
INVx1_ASAP7_75t_L g528 ( .A(n_199), .Y(n_528) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OAI21x1_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_214), .Y(n_200) );
AOI21x1_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B(n_208), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_207), .A2(n_239), .B(n_241), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_208), .A2(n_213), .B1(n_296), .B2(n_298), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_208), .A2(n_577), .B(n_578), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_213), .A2(n_221), .B1(n_222), .B2(n_223), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_213), .A2(n_590), .B1(n_648), .B2(n_650), .Y(n_647) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
OR2x2_ASAP7_75t_L g286 ( .A(n_217), .B(n_247), .Y(n_286) );
AND2x2_ASAP7_75t_L g436 ( .A(n_217), .B(n_320), .Y(n_436) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g264 ( .A(n_218), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g312 ( .A(n_218), .Y(n_312) );
AND2x2_ASAP7_75t_L g335 ( .A(n_218), .B(n_306), .Y(n_335) );
INVx1_ASAP7_75t_L g368 ( .A(n_218), .Y(n_368) );
AND2x2_ASAP7_75t_L g404 ( .A(n_218), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g409 ( .A(n_218), .B(n_265), .Y(n_409) );
AND2x2_ASAP7_75t_L g467 ( .A(n_218), .B(n_309), .Y(n_467) );
OR2x2_ASAP7_75t_L g476 ( .A(n_218), .B(n_248), .Y(n_476) );
AO31x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .A3(n_224), .B(n_225), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_227), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g352 ( .A(n_228), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_228), .B(n_305), .Y(n_393) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g322 ( .A(n_229), .Y(n_322) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g346 ( .A(n_230), .B(n_266), .Y(n_346) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_233), .B(n_243), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_231), .A2(n_233), .B(n_243), .Y(n_263) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_231), .A2(n_570), .B(n_579), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_231), .A2(n_610), .B(n_618), .Y(n_609) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_231), .A2(n_610), .B(n_618), .Y(n_633) );
OAI21xp33_ASAP7_75t_SL g642 ( .A1(n_231), .A2(n_570), .B(n_579), .Y(n_642) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g566 ( .A(n_232), .Y(n_566) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_238), .B(n_242), .Y(n_233) );
INVx2_ASAP7_75t_L g617 ( .A(n_237), .Y(n_617) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_242), .A2(n_251), .B(n_256), .Y(n_250) );
AOI31xp67_ASAP7_75t_L g267 ( .A1(n_242), .A2(n_268), .A3(n_269), .B(n_272), .Y(n_267) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_242), .A2(n_559), .B(n_562), .Y(n_558) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_242), .A2(n_571), .B(n_576), .Y(n_570) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_242), .A2(n_601), .B(n_604), .Y(n_600) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_242), .A2(n_611), .B(n_614), .Y(n_610) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_242), .A2(n_621), .B(n_624), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_275), .B1(n_283), .B2(n_285), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_246), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_264), .Y(n_246) );
INVx1_ASAP7_75t_L g417 ( .A(n_247), .Y(n_417) );
OR2x2_ASAP7_75t_L g530 ( .A(n_247), .B(n_426), .Y(n_530) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_263), .Y(n_247) );
INVx2_ASAP7_75t_SL g302 ( .A(n_248), .Y(n_302) );
BUFx2_ASAP7_75t_L g343 ( .A(n_248), .Y(n_343) );
AND2x2_ASAP7_75t_L g367 ( .A(n_248), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g405 ( .A(n_248), .Y(n_405) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_262), .Y(n_248) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_249), .A2(n_250), .B(n_262), .Y(n_309) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_249), .A2(n_600), .B(n_607), .Y(n_599) );
OA21x2_ASAP7_75t_L g619 ( .A1(n_249), .A2(n_620), .B(n_628), .Y(n_619) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_249), .A2(n_620), .B(n_628), .Y(n_645) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_249), .A2(n_600), .B(n_607), .Y(n_679) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_259), .B1(n_260), .B2(n_261), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_258), .A2(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_259), .A2(n_551), .B1(n_552), .B2(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g308 ( .A(n_263), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g468 ( .A(n_263), .B(n_306), .Y(n_468) );
INVx1_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g306 ( .A(n_267), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
AND2x2_ASAP7_75t_L g524 ( .A(n_277), .B(n_291), .Y(n_524) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g293 ( .A(n_279), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g328 ( .A(n_279), .Y(n_328) );
INVx1_ASAP7_75t_L g341 ( .A(n_279), .Y(n_341) );
INVx1_ASAP7_75t_L g433 ( .A(n_279), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_280), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g332 ( .A(n_280), .B(n_293), .Y(n_332) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g364 ( .A(n_282), .B(n_329), .Y(n_364) );
INVx1_ASAP7_75t_L g382 ( .A(n_282), .Y(n_382) );
INVx2_ASAP7_75t_L g477 ( .A(n_283), .Y(n_477) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI321xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_301), .A3(n_303), .B1(n_307), .B2(n_313), .C(n_316), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g313 ( .A(n_293), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g354 ( .A(n_293), .B(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g329 ( .A(n_294), .Y(n_329) );
AND2x2_ASAP7_75t_L g432 ( .A(n_294), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_302), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_304), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g377 ( .A(n_305), .Y(n_377) );
AND2x2_ASAP7_75t_L g439 ( .A(n_305), .B(n_368), .Y(n_439) );
AND2x2_ASAP7_75t_L g459 ( .A(n_305), .B(n_322), .Y(n_459) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g353 ( .A(n_306), .B(n_309), .Y(n_353) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
AND2x2_ASAP7_75t_L g438 ( .A(n_308), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g478 ( .A(n_308), .Y(n_478) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g316 ( .A1(n_310), .A2(n_317), .A3(n_319), .B1(n_324), .B2(n_326), .Y(n_316) );
OR2x2_ASAP7_75t_L g350 ( .A(n_310), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g344 ( .A(n_311), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_311), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g511 ( .A(n_311), .B(n_346), .Y(n_511) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g358 ( .A(n_312), .B(n_322), .Y(n_358) );
OR2x2_ASAP7_75t_L g527 ( .A(n_312), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_314), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g317 ( .A(n_315), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
OR2x2_ASAP7_75t_L g372 ( .A(n_315), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g505 ( .A(n_315), .B(n_432), .Y(n_505) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_315), .Y(n_519) );
INVx2_ASAP7_75t_L g456 ( .A(n_318), .Y(n_456) );
OR2x2_ASAP7_75t_L g497 ( .A(n_318), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g501 ( .A(n_319), .Y(n_501) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g515 ( .A(n_320), .B(n_335), .Y(n_515) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g376 ( .A(n_321), .B(n_377), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g472 ( .A(n_327), .Y(n_472) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
INVx1_ASAP7_75t_L g424 ( .A(n_329), .Y(n_424) );
NOR2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_347), .Y(n_330) );
AO22x1_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_336), .B2(n_342), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g426 ( .A(n_335), .Y(n_426) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_337), .A2(n_430), .B1(n_435), .B2(n_437), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g380 ( .A(n_341), .Y(n_380) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g408 ( .A(n_343), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g445 ( .A(n_343), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_344), .A2(n_450), .B1(n_483), .B2(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g366 ( .A(n_346), .Y(n_366) );
OR2x2_ASAP7_75t_L g491 ( .A(n_346), .B(n_476), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_370), .Y(n_347) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_354), .B(n_356), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_349), .A2(n_371), .B1(n_375), .B2(n_378), .Y(n_370) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_L g427 ( .A(n_352), .Y(n_427) );
AND2x2_ASAP7_75t_L g484 ( .A(n_352), .B(n_367), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_353), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g386 ( .A(n_355), .B(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_365), .B2(n_369), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_361), .B(n_373), .Y(n_483) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp33_ASAP7_75t_R g378 ( .A(n_363), .B(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g396 ( .A(n_364), .B(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g450 ( .A(n_364), .B(n_394), .Y(n_450) );
BUFx2_ASAP7_75t_L g513 ( .A(n_364), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g444 ( .A(n_366), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g488 ( .A(n_366), .B(n_404), .Y(n_488) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_373), .Y(n_443) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g461 ( .A(n_374), .B(n_398), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g509 ( .A(n_380), .Y(n_509) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g504 ( .A(n_382), .Y(n_504) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_406), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B(n_395), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_385), .A2(n_486), .B(n_494), .Y(n_485) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g455 ( .A(n_394), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g458 ( .A(n_404), .B(n_459), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_410), .B(n_413), .C(n_418), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g494 ( .A1(n_410), .A2(n_491), .B(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI211xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_425), .C(n_427), .Y(n_418) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_420), .Y(n_493) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g522 ( .A(n_427), .Y(n_522) );
NOR3x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_440), .C(n_448), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_438), .A2(n_442), .B1(n_444), .B2(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g523 ( .A(n_439), .Y(n_523) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_444), .B(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_444), .A2(n_518), .B1(n_521), .B2(n_524), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_444), .A2(n_461), .B1(n_526), .B2(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND4xp75_ASAP7_75t_L g451 ( .A(n_452), .B(n_485), .C(n_499), .D(n_516), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g452 ( .A(n_453), .B(n_469), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B1(n_460), .B2(n_462), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g464 ( .A(n_458), .Y(n_464) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g474 ( .A(n_468), .B(n_475), .Y(n_474) );
OAI321xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .A3(n_477), .B1(n_478), .B2(n_479), .C(n_482), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_472), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_474), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .B1(n_491), .B2(n_492), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_497), .Y(n_510) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_510), .B(n_511), .C(n_512), .Y(n_506) );
INVxp33_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
NOR2x1p5_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
BUFx8_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g915 ( .A(n_533), .B(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND4xp75_ASAP7_75t_L g535 ( .A(n_536), .B(n_728), .C(n_801), .D(n_860), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_684), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_654), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_595), .B1(n_629), .B2(n_634), .C(n_638), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI21xp33_ASAP7_75t_SL g638 ( .A1(n_540), .A2(n_639), .B(n_643), .Y(n_638) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_567), .Y(n_540) );
AND2x2_ASAP7_75t_L g681 ( .A(n_541), .B(n_641), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_541), .B(n_692), .Y(n_754) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_555), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g640 ( .A(n_543), .Y(n_640) );
INVx4_ASAP7_75t_L g660 ( .A(n_543), .Y(n_660) );
AND2x2_ASAP7_75t_L g688 ( .A(n_543), .B(n_568), .Y(n_688) );
OR2x2_ASAP7_75t_L g850 ( .A(n_543), .B(n_637), .Y(n_850) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_550), .B(n_554), .Y(n_545) );
INVx2_ASAP7_75t_L g663 ( .A(n_555), .Y(n_663) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_555), .Y(n_689) );
INVx1_ASAP7_75t_L g699 ( .A(n_555), .Y(n_699) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g637 ( .A(n_556), .Y(n_637) );
AND2x2_ASAP7_75t_L g790 ( .A(n_556), .B(n_581), .Y(n_790) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_565), .Y(n_556) );
INVx2_ASAP7_75t_L g747 ( .A(n_567), .Y(n_747) );
AND2x2_ASAP7_75t_L g751 ( .A(n_567), .B(n_663), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_567), .B(n_782), .Y(n_880) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_580), .Y(n_567) );
INVx2_ASAP7_75t_L g714 ( .A(n_568), .Y(n_714) );
AND2x2_ASAP7_75t_L g808 ( .A(n_568), .B(n_674), .Y(n_808) );
AND2x2_ASAP7_75t_L g859 ( .A(n_568), .B(n_660), .Y(n_859) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g641 ( .A(n_580), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g662 ( .A(n_581), .Y(n_662) );
AOI21x1_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_594), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_608), .Y(n_596) );
INVx2_ASAP7_75t_L g630 ( .A(n_597), .Y(n_630) );
AND2x2_ASAP7_75t_L g791 ( .A(n_597), .B(n_644), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_597), .B(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_597), .B(n_812), .Y(n_821) );
OR2x2_ASAP7_75t_L g844 ( .A(n_597), .B(n_703), .Y(n_844) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp67_ASAP7_75t_L g727 ( .A(n_598), .B(n_670), .Y(n_727) );
AND2x2_ASAP7_75t_L g833 ( .A(n_598), .B(n_645), .Y(n_833) );
BUFx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g667 ( .A(n_599), .Y(n_667) );
AND2x2_ASAP7_75t_L g720 ( .A(n_608), .B(n_665), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_608), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_608), .B(n_776), .Y(n_784) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_619), .Y(n_608) );
AND2x2_ASAP7_75t_L g696 ( .A(n_609), .B(n_645), .Y(n_696) );
INVx1_ASAP7_75t_L g840 ( .A(n_609), .Y(n_840) );
AND2x2_ASAP7_75t_L g631 ( .A(n_619), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g703 ( .A(n_619), .B(n_646), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_619), .B(n_646), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_630), .B(n_744), .Y(n_743) );
AND2x4_ASAP7_75t_L g866 ( .A(n_630), .B(n_669), .Y(n_866) );
AND2x2_ASAP7_75t_L g796 ( .A(n_631), .B(n_797), .Y(n_796) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_632), .Y(n_653) );
AND2x2_ASAP7_75t_L g677 ( .A(n_632), .B(n_678), .Y(n_677) );
BUFx3_ASAP7_75t_L g683 ( .A(n_632), .Y(n_683) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_632), .Y(n_719) );
INVx1_ASAP7_75t_L g744 ( .A(n_632), .Y(n_744) );
AND2x2_ASAP7_75t_L g750 ( .A(n_632), .B(n_645), .Y(n_750) );
INVx1_ASAP7_75t_L g831 ( .A(n_632), .Y(n_831) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g673 ( .A(n_635), .B(n_674), .Y(n_673) );
AOI32xp33_ASAP7_75t_SL g805 ( .A1(n_635), .A2(n_697), .A3(n_806), .B1(n_808), .B2(n_809), .Y(n_805) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx2_ASAP7_75t_L g658 ( .A(n_636), .Y(n_658) );
OR2x2_ASAP7_75t_L g707 ( .A(n_636), .B(n_663), .Y(n_707) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_637), .Y(n_711) );
INVxp67_ASAP7_75t_L g737 ( .A(n_637), .Y(n_737) );
OR2x2_ASAP7_75t_L g839 ( .A(n_637), .B(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OR3x2_ASAP7_75t_L g704 ( .A(n_640), .B(n_705), .C(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g810 ( .A(n_640), .Y(n_810) );
AND2x2_ASAP7_75t_L g738 ( .A(n_641), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g794 ( .A(n_641), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_641), .B(n_689), .Y(n_800) );
BUFx2_ASAP7_75t_L g693 ( .A(n_642), .Y(n_693) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_653), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_644), .B(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_644), .Y(n_873) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g670 ( .A(n_645), .Y(n_670) );
INVx1_ASAP7_75t_L g812 ( .A(n_645), .Y(n_812) );
INVx1_ASAP7_75t_L g671 ( .A(n_646), .Y(n_671) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_646), .Y(n_717) );
OR2x2_ASAP7_75t_L g758 ( .A(n_646), .B(n_679), .Y(n_758) );
AND2x2_ASAP7_75t_L g776 ( .A(n_646), .B(n_679), .Y(n_776) );
AND2x2_ASAP7_75t_L g797 ( .A(n_646), .B(n_667), .Y(n_797) );
BUFx2_ASAP7_75t_L g865 ( .A(n_653), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_672), .C(n_680), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_664), .Y(n_655) );
INVx3_ASAP7_75t_L g787 ( .A(n_656), .Y(n_787) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_661), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x2_ASAP7_75t_L g817 ( .A(n_658), .B(n_773), .Y(n_817) );
INVx1_ASAP7_75t_L g739 ( .A(n_659), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_659), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g824 ( .A(n_659), .B(n_663), .Y(n_824) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g698 ( .A(n_660), .B(n_699), .Y(n_698) );
NAND2x1_ASAP7_75t_L g713 ( .A(n_660), .B(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g782 ( .A(n_660), .Y(n_782) );
NAND2xp33_ASAP7_75t_R g765 ( .A(n_661), .B(n_688), .Y(n_765) );
AND2x2_ASAP7_75t_L g781 ( .A(n_661), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g847 ( .A(n_661), .Y(n_847) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx2_ASAP7_75t_L g674 ( .A(n_662), .Y(n_674) );
INVx1_ASAP7_75t_L g706 ( .A(n_662), .Y(n_706) );
INVx2_ASAP7_75t_L g773 ( .A(n_662), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_663), .B(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g695 ( .A(n_666), .B(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g682 ( .A(n_669), .B(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g853 ( .A(n_669), .B(n_744), .Y(n_853) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AND2x2_ASAP7_75t_L g734 ( .A(n_671), .B(n_679), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g701 ( .A(n_677), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g804 ( .A(n_678), .Y(n_804) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx2_ASAP7_75t_L g862 ( .A(n_681), .Y(n_862) );
INVx1_ASAP7_75t_L g690 ( .A(n_682), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_683), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g760 ( .A(n_683), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g807 ( .A(n_683), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g856 ( .A(n_683), .B(n_757), .Y(n_856) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_691), .C(n_708), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g722 ( .A(n_688), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g815 ( .A(n_688), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B1(n_700), .B2(n_704), .Y(n_691) );
NAND3x2_ASAP7_75t_L g834 ( .A(n_692), .B(n_835), .C(n_836), .Y(n_834) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
NAND2x1_ASAP7_75t_L g774 ( .A(n_696), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g746 ( .A(n_698), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g818 ( .A(n_698), .Y(n_818) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g870 ( .A(n_702), .B(n_803), .Y(n_870) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g732 ( .A(n_703), .Y(n_732) );
NOR2x1p5_ASAP7_75t_SL g779 ( .A(n_705), .B(n_707), .Y(n_779) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g723 ( .A(n_706), .Y(n_723) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_706), .Y(n_825) );
OAI22xp33_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_715), .B1(n_721), .B2(n_724), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g868 ( .A(n_711), .B(n_815), .Y(n_868) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g788 ( .A(n_713), .B(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_SL g715 ( .A(n_716), .B(n_720), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g770 ( .A(n_717), .Y(n_770) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_722), .A2(n_838), .B1(n_843), .B2(n_845), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_722), .A2(n_816), .B1(n_873), .B2(n_874), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_722), .B(n_870), .Y(n_877) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_762), .Y(n_728) );
NAND3xp33_ASAP7_75t_SL g729 ( .A(n_730), .B(n_740), .C(n_752), .Y(n_729) );
AO21x1_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g832 ( .A(n_731), .Y(n_832) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2x1p5_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
AOI32xp33_ASAP7_75t_L g852 ( .A1(n_736), .A2(n_853), .A3(n_854), .B1(n_855), .B2(n_857), .Y(n_852) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g835 ( .A(n_739), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_745), .B1(n_748), .B2(n_751), .Y(n_740) );
INVxp67_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g768 ( .A(n_744), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_744), .B(n_776), .Y(n_777) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_745), .A2(n_753), .B1(n_755), .B2(n_759), .Y(n_752) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g849 ( .A(n_747), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI322xp33_ASAP7_75t_L g861 ( .A1(n_749), .A2(n_842), .A3(n_862), .B1(n_863), .B2(n_867), .C1(n_868), .C2(n_869), .Y(n_861) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g881 ( .A(n_750), .B(n_770), .Y(n_881) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g842 ( .A(n_758), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_759), .B(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g799 ( .A(n_761), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_785), .Y(n_762) );
AOI211xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B(n_771), .C(n_780), .Y(n_763) );
INVxp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B1(n_777), .B2(n_778), .Y(n_771) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_776), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_776), .B(n_812), .Y(n_875) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_791), .B(n_792), .Y(n_785) );
NAND2x1_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
NOR2x1_ASAP7_75t_SL g814 ( .A(n_789), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g836 ( .A(n_789), .Y(n_836) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g851 ( .A(n_791), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B1(n_798), .B2(n_800), .Y(n_792) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g854 ( .A(n_794), .Y(n_854) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR3x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_826), .C(n_848), .Y(n_801) );
OAI211xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B(n_813), .C(n_822), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVxp67_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g820 ( .A(n_807), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_808), .B(n_810), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI21xp5_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_816), .B(n_819), .Y(n_813) );
AND2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVxp67_ASAP7_75t_L g867 ( .A(n_817), .Y(n_867) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_834), .B(n_837), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_832), .C(n_833), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_SL g845 ( .A(n_846), .B(n_847), .Y(n_845) );
OAI21xp5_ASAP7_75t_SL g848 ( .A1(n_849), .A2(n_851), .B(n_852), .Y(n_848) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
NOR3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_871), .C(n_876), .Y(n_860) );
NAND2x1p5_ASAP7_75t_L g863 ( .A(n_864), .B(n_866), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND2xp33_ASAP7_75t_SL g876 ( .A(n_877), .B(n_878), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_881), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
OAI21xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_890), .B(n_902), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_884), .Y(n_883) );
INVx5_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
CKINVDCx8_ASAP7_75t_R g907 ( .A(n_886), .Y(n_907) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_896), .B1(n_897), .B2(n_901), .Y(n_891) );
INVx2_ASAP7_75t_SL g901 ( .A(n_892), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_908), .Y(n_902) );
NOR2xp67_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
INVx4_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx3_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
BUFx10_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_920), .Y(n_919) );
CKINVDCx6p67_ASAP7_75t_R g920 ( .A(n_921), .Y(n_920) );
endmodule