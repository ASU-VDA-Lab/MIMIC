module fake_jpeg_12844_n_555 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_555);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_555;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_62),
.B(n_96),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_69),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_70),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_55),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_72),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_79),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_84),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_23),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_92),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_95),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_16),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx2_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_98),
.B(n_1),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_99),
.B(n_100),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_37),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_103),
.Y(n_183)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_118),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_42),
.B(n_16),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_36),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_54),
.Y(n_146)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_42),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_125),
.Y(n_199)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_123),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_21),
.B(n_15),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_0),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_34),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_48),
.B1(n_38),
.B2(n_43),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_131),
.A2(n_135),
.B1(n_159),
.B2(n_114),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_133),
.B(n_172),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_77),
.A2(n_48),
.B1(n_38),
.B2(n_43),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_25),
.B1(n_43),
.B2(n_49),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_69),
.A2(n_25),
.B1(n_49),
.B2(n_48),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_87),
.A2(n_38),
.B1(n_46),
.B2(n_45),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_69),
.A2(n_49),
.B1(n_46),
.B2(n_51),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_146),
.B(n_63),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_148),
.B(n_160),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_70),
.A2(n_46),
.B1(n_53),
.B2(n_51),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_149),
.A2(n_163),
.B1(n_171),
.B2(n_178),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_82),
.B(n_28),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_162),
.B(n_190),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_70),
.A2(n_57),
.B1(n_35),
.B2(n_53),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_88),
.A2(n_57),
.B1(n_35),
.B2(n_47),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_164),
.A2(n_140),
.B(n_187),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_80),
.A2(n_47),
.B1(n_39),
.B2(n_33),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_98),
.B(n_93),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_67),
.A2(n_39),
.B1(n_33),
.B2(n_30),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_211),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_74),
.A2(n_54),
.B1(n_3),
.B2(n_4),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_181),
.A2(n_208),
.B1(n_94),
.B2(n_109),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_2),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_80),
.A2(n_106),
.B1(n_113),
.B2(n_71),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_197),
.A2(n_202),
.B1(n_213),
.B2(n_11),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_89),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_200),
.B(n_201),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_60),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_106),
.A2(n_76),
.B1(n_75),
.B2(n_65),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_85),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_120),
.B(n_4),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_73),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_220),
.B(n_238),
.Y(n_334)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_221),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_115),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_222),
.B(n_227),
.Y(n_320)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_155),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_224),
.B(n_225),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_127),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_226),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_115),
.Y(n_227)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_229),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_133),
.A2(n_107),
.B1(n_116),
.B2(n_112),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_231),
.B1(n_245),
.B2(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_232),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_233),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_110),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_234),
.B(n_244),
.Y(n_311)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_235),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_239),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_240),
.B(n_286),
.C(n_210),
.Y(n_340)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_241),
.Y(n_339)
);

AO22x1_ASAP7_75t_SL g242 ( 
.A1(n_147),
.A2(n_104),
.B1(n_72),
.B2(n_121),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_252),
.Y(n_289)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_184),
.B(n_95),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_142),
.A2(n_108),
.B1(n_101),
.B2(n_90),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_111),
.B1(n_8),
.B2(n_9),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_246),
.A2(n_212),
.B1(n_137),
.B2(n_196),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_172),
.A2(n_111),
.B(n_8),
.C(n_9),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_247),
.A2(n_248),
.B(n_213),
.C(n_204),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_194),
.A2(n_5),
.B(n_8),
.C(n_9),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_251),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_9),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx11_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_157),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_128),
.B(n_183),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_161),
.Y(n_257)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx6_ASAP7_75t_SL g258 ( 
.A(n_134),
.Y(n_258)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_150),
.B(n_10),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_171),
.B(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_266),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_177),
.Y(n_264)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_174),
.Y(n_265)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_166),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_268),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_143),
.B(n_175),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_269),
.B(n_271),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_208),
.A2(n_12),
.B1(n_181),
.B2(n_141),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_153),
.B(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_273),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_167),
.B(n_12),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_167),
.B(n_176),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_276),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_179),
.B(n_138),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_134),
.A2(n_187),
.B1(n_132),
.B2(n_138),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_161),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_282),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_285),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_284),
.A2(n_204),
.B(n_169),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_163),
.B(n_130),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_186),
.B(n_130),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_216),
.B(n_240),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_313),
.C(n_238),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_SL g362 ( 
.A1(n_298),
.A2(n_325),
.B(n_255),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_220),
.A2(n_149),
.B1(n_144),
.B2(n_202),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_309),
.A2(n_326),
.B1(n_132),
.B2(n_286),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_217),
.A2(n_285),
.A3(n_218),
.B1(n_247),
.B2(n_237),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_226),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_216),
.B(n_169),
.C(n_166),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_231),
.A2(n_168),
.B1(n_212),
.B2(n_137),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_327),
.A2(n_328),
.B1(n_182),
.B2(n_185),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_270),
.A2(n_236),
.B1(n_228),
.B2(n_245),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_252),
.B(n_216),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_336),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_240),
.B(n_168),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_242),
.B(n_205),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_337),
.B(n_196),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_286),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_295),
.B(n_250),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_341),
.B(n_345),
.Y(n_415)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_343),
.B(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_292),
.B(n_284),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_348),
.C(n_375),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_248),
.B(n_258),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_242),
.C(n_273),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_254),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_349),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_302),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_350),
.Y(n_391)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_351),
.Y(n_411)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_354),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_321),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_372),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_321),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_357),
.Y(n_392)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_358),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g359 ( 
.A(n_331),
.B(n_272),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_359),
.A2(n_360),
.B(n_364),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_282),
.B(n_233),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_253),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_361),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_362),
.A2(n_363),
.B(n_365),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_303),
.A2(n_266),
.B(n_215),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_277),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_337),
.A2(n_205),
.B1(n_235),
.B2(n_223),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_366),
.A2(n_371),
.B1(n_287),
.B2(n_297),
.Y(n_400)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_374),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_328),
.A2(n_246),
.B1(n_185),
.B2(n_182),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_368),
.A2(n_381),
.B1(n_326),
.B2(n_312),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_289),
.A2(n_241),
.B1(n_265),
.B2(n_229),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_334),
.A2(n_313),
.B(n_322),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_269),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_373),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_295),
.B(n_243),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_261),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_377),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_333),
.A2(n_265),
.B1(n_221),
.B2(n_283),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_378),
.A2(n_294),
.B1(n_264),
.B2(n_323),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_288),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_293),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_289),
.B(n_281),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_324),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_382),
.A2(n_384),
.B1(n_389),
.B2(n_393),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_368),
.A2(n_333),
.B1(n_305),
.B2(n_322),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_381),
.A2(n_305),
.B1(n_319),
.B2(n_336),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_310),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_409),
.C(n_414),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_342),
.A2(n_319),
.B1(n_298),
.B2(n_327),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_344),
.A2(n_348),
.B1(n_359),
.B2(n_360),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_398),
.A2(n_404),
.B1(n_371),
.B2(n_369),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_402),
.B1(n_357),
.B2(n_339),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_364),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_370),
.A2(n_380),
.B1(n_376),
.B2(n_363),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_359),
.A2(n_312),
.B1(n_296),
.B2(n_330),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_405),
.A2(n_354),
.B(n_356),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_338),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_351),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_300),
.C(n_332),
.Y(n_414)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_390),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_419),
.C(n_420),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_355),
.C(n_375),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_412),
.C(n_386),
.Y(n_420)
);

AOI22x1_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_365),
.B1(n_372),
.B2(n_369),
.Y(n_422)
);

AO22x1_ASAP7_75t_SL g466 ( 
.A1(n_422),
.A2(n_444),
.B1(n_405),
.B2(n_324),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_359),
.Y(n_423)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_341),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_427),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_425),
.A2(n_440),
.B1(n_408),
.B2(n_394),
.Y(n_456)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_411),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_345),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_374),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_431),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_365),
.C(n_352),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_439),
.C(n_419),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_433),
.A2(n_438),
.B(n_441),
.Y(n_464)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_415),
.B(n_353),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_442),
.B1(n_443),
.B2(n_388),
.Y(n_447)
);

MAJx2_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_401),
.C(n_339),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_387),
.A2(n_304),
.B(n_317),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_398),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_389),
.A2(n_366),
.B1(n_330),
.B2(n_367),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_403),
.A2(n_393),
.B(n_387),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

OA22x2_ASAP7_75t_L g444 ( 
.A1(n_384),
.A2(n_317),
.B1(n_307),
.B2(n_291),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_414),
.B(n_318),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_404),
.Y(n_461)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_443),
.A2(n_408),
.B1(n_395),
.B2(n_382),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_456),
.Y(n_477)
);

FAx1_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_407),
.CI(n_400),
.CON(n_450),
.SN(n_450)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_450),
.A2(n_459),
.B(n_462),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_441),
.A2(n_407),
.B(n_403),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_468),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_460),
.C(n_467),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_421),
.A2(n_394),
.B1(n_383),
.B2(n_410),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_420),
.C(n_417),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_461),
.B(n_444),
.Y(n_491)
);

A2O1A1O1Ixp25_ASAP7_75t_L g462 ( 
.A1(n_422),
.A2(n_406),
.B(n_385),
.C(n_392),
.D(n_388),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_385),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_421),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_392),
.C(n_307),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_416),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_423),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_425),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_472),
.B(n_481),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_432),
.C(n_445),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_486),
.C(n_489),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_479),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_377),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_460),
.B(n_442),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_482),
.B(n_485),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_471),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_491),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_435),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_487),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_448),
.B(n_434),
.C(n_444),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_438),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_488),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_433),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_440),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_490),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_444),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_494),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_473),
.A2(n_462),
.B(n_459),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_497),
.A2(n_506),
.B(n_464),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_478),
.A2(n_456),
.B1(n_452),
.B2(n_446),
.Y(n_498)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_480),
.A2(n_446),
.B1(n_452),
.B2(n_453),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_505),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_484),
.A2(n_454),
.B(n_464),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_477),
.A2(n_453),
.B1(n_457),
.B2(n_463),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_449),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_484),
.B(n_457),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_508),
.B(n_492),
.Y(n_509)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_514),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_513),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_486),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_479),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g515 ( 
.A(n_496),
.B(n_450),
.CI(n_476),
.CON(n_515),
.SN(n_515)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_487),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_508),
.A2(n_450),
.B1(n_466),
.B2(n_491),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_516),
.A2(n_498),
.B1(n_466),
.B2(n_499),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_474),
.C(n_475),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_518),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_474),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_504),
.C(n_506),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_489),
.C(n_497),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_522),
.A2(n_515),
.B(n_510),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_513),
.C(n_520),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_524),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_502),
.C(n_504),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_528),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_500),
.C(n_499),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_529),
.A2(n_522),
.B1(n_521),
.B2(n_511),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_470),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_495),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_510),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_533),
.B(n_534),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_536),
.A2(n_533),
.B(n_539),
.Y(n_546)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_538),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_532),
.A2(n_516),
.B1(n_495),
.B2(n_515),
.Y(n_539)
);

AO21x1_ASAP7_75t_L g545 ( 
.A1(n_539),
.A2(n_540),
.B(n_294),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_535),
.A2(n_526),
.B(n_525),
.Y(n_542)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_542),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_537),
.A2(n_530),
.B(n_290),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_543),
.B(n_545),
.C(n_546),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_534),
.C(n_536),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_547),
.B(n_544),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_550),
.A2(n_551),
.B(n_214),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_548),
.A2(n_538),
.B(n_290),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_552),
.A2(n_239),
.B(n_257),
.Y(n_553)
);

AOI31xp33_ASAP7_75t_L g554 ( 
.A1(n_553),
.A2(n_280),
.A3(n_210),
.B(n_186),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_329),
.B(n_258),
.Y(n_555)
);


endmodule