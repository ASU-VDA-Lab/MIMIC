module fake_jpeg_11588_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_20),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_57),
.B(n_58),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_62),
.Y(n_132)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_69),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_30),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_65),
.B(n_76),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_66),
.B(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_1),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_15),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_73),
.Y(n_131)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_23),
.B(n_15),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_78),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_79),
.B(n_85),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_1),
.Y(n_86)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_1),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_98),
.C(n_99),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_2),
.Y(n_93)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_19),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_96),
.A2(n_48),
.B1(n_47),
.B2(n_44),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_27),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_29),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_29),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_102),
.B1(n_43),
.B2(n_38),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

BUFx16f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_33),
.B1(n_50),
.B2(n_19),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_105),
.A2(n_115),
.B1(n_127),
.B2(n_152),
.Y(n_199)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_33),
.B1(n_50),
.B2(n_19),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_25),
.B1(n_41),
.B2(n_50),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_96),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_64),
.A2(n_41),
.B1(n_25),
.B2(n_31),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_122),
.A2(n_160),
.B1(n_44),
.B2(n_39),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_56),
.A2(n_41),
.B1(n_25),
.B2(n_33),
.Y(n_123)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_41),
.B1(n_25),
.B2(n_34),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_55),
.A2(n_60),
.B1(n_82),
.B2(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_58),
.A2(n_52),
.B1(n_31),
.B2(n_35),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_128),
.B(n_3),
.Y(n_213)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_74),
.Y(n_179)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_31),
.B1(n_52),
.B2(n_34),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_103),
.A2(n_52),
.B1(n_34),
.B2(n_51),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_155),
.A2(n_89),
.B1(n_6),
.B2(n_7),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_163),
.B(n_166),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_164),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_75),
.B1(n_77),
.B2(n_80),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_168),
.A2(n_197),
.B1(n_135),
.B2(n_156),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_73),
.B(n_91),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_169),
.A2(n_8),
.B(n_9),
.Y(n_249)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_173),
.B(n_185),
.Y(n_260)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_178),
.B1(n_188),
.B2(n_158),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_95),
.B1(n_90),
.B2(n_68),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_67),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_209),
.C(n_62),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_78),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_71),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_123),
.A2(n_72),
.B1(n_87),
.B2(n_63),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_79),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_189),
.B(n_212),
.Y(n_254)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_193),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_121),
.A2(n_65),
.B1(n_100),
.B2(n_99),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_139),
.B(n_89),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_130),
.B(n_97),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_198),
.Y(n_251)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_196),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_85),
.B1(n_43),
.B2(n_48),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_132),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_203),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g201 ( 
.A(n_132),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_51),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_157),
.B(n_47),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_125),
.B(n_129),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_210),
.Y(n_227)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_136),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_211),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_109),
.B(n_89),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_39),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_155),
.A2(n_62),
.B(n_4),
.C(n_5),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_216),
.B1(n_134),
.B2(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_215),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_3),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_218),
.A2(n_236),
.B1(n_237),
.B2(n_263),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_222),
.B(n_223),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_105),
.B1(n_115),
.B2(n_152),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_228),
.B1(n_233),
.B2(n_234),
.Y(n_269)
);

OAI22x1_ASAP7_75t_SL g228 ( 
.A1(n_179),
.A2(n_127),
.B1(n_134),
.B2(n_138),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_248),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_156),
.B1(n_119),
.B2(n_150),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_176),
.A2(n_162),
.B1(n_135),
.B2(n_150),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_162),
.B1(n_139),
.B2(n_116),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_240),
.B1(n_241),
.B2(n_244),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_179),
.A2(n_120),
.B1(n_101),
.B2(n_151),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_192),
.A2(n_151),
.B1(n_6),
.B2(n_7),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_180),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_192),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_189),
.B(n_181),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_245),
.B(n_184),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_249),
.B(n_201),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_177),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_181),
.B(n_8),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_267),
.C(n_182),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_178),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_13),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_169),
.B(n_12),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_192),
.B1(n_191),
.B2(n_175),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_268),
.A2(n_236),
.B1(n_218),
.B2(n_237),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_172),
.B(n_163),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_271),
.B(n_282),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_239),
.B(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_215),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_287),
.C(n_305),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_274),
.B(n_275),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_225),
.A2(n_211),
.B1(n_183),
.B2(n_212),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_280),
.A2(n_281),
.B1(n_222),
.B2(n_223),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_248),
.A2(n_214),
.B1(n_195),
.B2(n_170),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_239),
.A2(n_198),
.B(n_201),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_166),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_288),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_296),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_239),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_286),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_171),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_231),
.A2(n_171),
.B(n_167),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_289),
.A2(n_290),
.B(n_295),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_SL g292 ( 
.A(n_243),
.B(n_167),
.Y(n_292)
);

HAxp5_ASAP7_75t_SL g317 ( 
.A(n_292),
.B(n_250),
.CON(n_317),
.SN(n_317)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_247),
.B(n_165),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_293),
.B(n_298),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_227),
.Y(n_295)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_177),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_190),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_304),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_247),
.B(n_165),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_300),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_228),
.A2(n_217),
.B(n_184),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_301),
.Y(n_354)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_204),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_217),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_311),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_196),
.C(n_164),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_256),
.C(n_230),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_206),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_249),
.B(n_186),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_317),
.B(n_305),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_261),
.B1(n_238),
.B2(n_234),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_324),
.B1(n_327),
.B2(n_341),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_297),
.A2(n_261),
.B1(n_238),
.B2(n_233),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_326),
.A2(n_329),
.B1(n_353),
.B2(n_290),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_270),
.A2(n_244),
.B1(n_255),
.B2(n_246),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_269),
.A2(n_263),
.B1(n_229),
.B2(n_255),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_285),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_339),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_346),
.C(n_282),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_285),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_246),
.B1(n_221),
.B2(n_252),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_271),
.A2(n_221),
.B1(n_252),
.B2(n_230),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_342),
.A2(n_348),
.B1(n_349),
.B2(n_303),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_267),
.C(n_235),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_269),
.A2(n_230),
.B1(n_196),
.B2(n_224),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_283),
.A2(n_224),
.B1(n_266),
.B2(n_258),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_279),
.A2(n_265),
.B1(n_262),
.B2(n_266),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_288),
.Y(n_355)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_355),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_292),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_367),
.C(n_378),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_334),
.B(n_306),
.Y(n_361)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_335),
.B(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_337),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_364),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_349),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_368),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_273),
.Y(n_367)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_294),
.C(n_300),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_336),
.B(n_294),
.Y(n_369)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_301),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_370),
.A2(n_390),
.B(n_352),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_330),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_376),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_315),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_341),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_379),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_330),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_307),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NOR2x1p5_ASAP7_75t_SL g384 ( 
.A(n_327),
.B(n_279),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_384),
.A2(n_324),
.B1(n_354),
.B2(n_348),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_289),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_385),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_322),
.A2(n_268),
.B1(n_277),
.B2(n_313),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_354),
.B1(n_314),
.B2(n_329),
.Y(n_393)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_316),
.B(n_304),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_351),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_330),
.A2(n_313),
.B(n_284),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_391),
.A2(n_399),
.B(n_296),
.Y(n_433)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_386),
.B1(n_358),
.B2(n_370),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_400),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_371),
.A2(n_318),
.B(n_314),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_315),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_346),
.C(n_323),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_404),
.C(n_405),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_323),
.C(n_316),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_286),
.C(n_331),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_331),
.C(n_352),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_410),
.C(n_411),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_409),
.A2(n_417),
.B1(n_370),
.B2(n_374),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_345),
.C(n_274),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_298),
.C(n_333),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_356),
.B(n_333),
.C(n_350),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_418),
.C(n_420),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_360),
.A2(n_351),
.B1(n_325),
.B2(n_353),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_343),
.C(n_347),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_343),
.C(n_310),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_412),
.B(n_363),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_426),
.B(n_427),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

XOR2x1_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_393),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_380),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_431),
.B(n_435),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_384),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_449),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_433),
.A2(n_439),
.B(n_441),
.Y(n_469)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_397),
.Y(n_434)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_434),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_258),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_402),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_438),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_421),
.Y(n_437)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_407),
.A2(n_377),
.B1(n_366),
.B2(n_384),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_399),
.A2(n_296),
.B(n_383),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_326),
.B1(n_387),
.B2(n_373),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_442),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_381),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_445),
.Y(n_450)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_447),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_362),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_420),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_448),
.A2(n_404),
.B1(n_406),
.B2(n_410),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_362),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_392),
.C(n_403),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_452),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_443),
.A2(n_409),
.B1(n_406),
.B2(n_408),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_467),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_430),
.C(n_444),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_455),
.B(n_460),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_425),
.B(n_398),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_456),
.B(n_425),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_392),
.C(n_405),
.Y(n_460)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_391),
.C(n_394),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_465),
.C(n_466),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_401),
.C(n_415),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_357),
.C(n_344),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_424),
.A2(n_357),
.B1(n_311),
.B2(n_344),
.Y(n_467)
);

BUFx12_ASAP7_75t_L g468 ( 
.A(n_427),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_468),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_466),
.Y(n_472)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_472),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_448),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_474),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_449),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_447),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_477),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_432),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_482),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_452),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_437),
.Y(n_480)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_424),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_456),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_469),
.A2(n_433),
.B(n_441),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_485),
.A2(n_469),
.B(n_439),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_470),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_487),
.B(n_458),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_496),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_451),
.C(n_460),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_493),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_463),
.C(n_454),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_441),
.B(n_468),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_450),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_459),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_504),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_480),
.B(n_485),
.Y(n_499)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_499),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_500),
.B(n_442),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_486),
.A2(n_423),
.B1(n_436),
.B2(n_471),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_321),
.B1(n_312),
.B2(n_278),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_481),
.A2(n_423),
.B(n_468),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_479),
.B(n_486),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_438),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_472),
.C(n_484),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_509),
.Y(n_521)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_507),
.A2(n_508),
.B(n_514),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_489),
.A2(n_429),
.B(n_467),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_511),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_440),
.C(n_434),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_504),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_490),
.A2(n_321),
.B(n_278),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_497),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_494),
.C(n_496),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_519),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_498),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_520),
.B(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_517),
.B(n_503),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_516),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_498),
.Y(n_526)
);

XOR2x2_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_511),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_518),
.A2(n_506),
.B(n_507),
.Y(n_528)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_528),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_531),
.C(n_525),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_530),
.B(n_523),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_532),
.B(n_527),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_521),
.C(n_524),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_535),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_534),
.B1(n_536),
.B2(n_512),
.Y(n_538)
);

A2O1A1O1Ixp25_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_491),
.B(n_276),
.C(n_312),
.D(n_13),
.Y(n_539)
);


endmodule