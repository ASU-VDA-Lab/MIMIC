module fake_jpeg_12126_n_577 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_577);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_577;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_1),
.B(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_102),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_9),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_62),
.B(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_10),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_74),
.B(n_81),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g162 ( 
.A(n_80),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_10),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_86),
.Y(n_172)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_30),
.A2(n_10),
.B1(n_17),
.B2(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_36),
.B1(n_46),
.B2(n_35),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_16),
.Y(n_157)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_50),
.B(n_8),
.Y(n_101)
);

NAND2xp67_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_17),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_8),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_104),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_30),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_30),
.Y(n_120)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_120),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_29),
.C(n_42),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_52),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_123),
.B(n_135),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_52),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_79),
.B1(n_70),
.B2(n_108),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_60),
.A2(n_53),
.B1(n_29),
.B2(n_41),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_72),
.A2(n_53),
.B1(n_29),
.B2(n_41),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_73),
.A2(n_53),
.B1(n_51),
.B2(n_41),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_55),
.A2(n_45),
.B1(n_51),
.B2(n_33),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_49),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_46),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_43),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_167),
.B(n_107),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_80),
.A2(n_33),
.B1(n_48),
.B2(n_51),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_168),
.A2(n_89),
.B1(n_75),
.B2(n_69),
.Y(n_221)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_183),
.Y(n_241)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_184),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_35),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_185),
.B(n_195),
.Y(n_273)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_189),
.B(n_196),
.Y(n_253)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_109),
.A2(n_104),
.B(n_94),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_166),
.B(n_48),
.Y(n_239)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_114),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_197),
.A2(n_124),
.B1(n_151),
.B2(n_110),
.Y(n_257)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_83),
.B1(n_63),
.B2(n_64),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_201),
.A2(n_45),
.B1(n_20),
.B2(n_40),
.Y(n_284)
);

BUFx4f_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_138),
.Y(n_204)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_205),
.B(n_212),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_211),
.Y(n_285)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_131),
.B(n_43),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_214),
.B(n_222),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_142),
.A2(n_105),
.B1(n_48),
.B2(n_98),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_215),
.A2(n_228),
.B1(n_230),
.B2(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_155),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_220),
.Y(n_270)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_111),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_166),
.B1(n_130),
.B2(n_124),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_152),
.B(n_36),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_32),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

BUFx4f_ASAP7_75t_SL g255 ( 
.A(n_226),
.Y(n_255)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_168),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_231),
.B(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_234),
.A2(n_235),
.B1(n_139),
.B2(n_116),
.Y(n_268)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_112),
.Y(n_235)
);

OAI32xp33_ASAP7_75t_L g236 ( 
.A1(n_164),
.A2(n_130),
.A3(n_142),
.B1(n_112),
.B2(n_143),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_186),
.A2(n_148),
.B1(n_118),
.B2(n_143),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_238),
.A2(n_257),
.B1(n_261),
.B2(n_279),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_239),
.A2(n_291),
.B(n_1),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_175),
.B(n_65),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_242),
.B(n_248),
.C(n_258),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_246),
.A2(n_269),
.B1(n_196),
.B2(n_194),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_59),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_176),
.B(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_259),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_106),
.C(n_58),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_32),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_197),
.A2(n_148),
.B1(n_139),
.B2(n_118),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_174),
.A2(n_85),
.B1(n_95),
.B2(n_92),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_218),
.A2(n_86),
.B1(n_116),
.B2(n_173),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_219),
.B(n_49),
.CI(n_12),
.CON(n_278),
.SN(n_278)
);

MAJIxp5_ASAP7_75t_SL g337 ( 
.A(n_278),
.B(n_11),
.C(n_12),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_197),
.A2(n_71),
.B1(n_173),
.B2(n_45),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_289),
.B1(n_226),
.B2(n_187),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_191),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_219),
.A2(n_0),
.B(n_1),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_197),
.A2(n_210),
.B1(n_230),
.B2(n_207),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_292),
.A2(n_194),
.B1(n_193),
.B2(n_198),
.Y(n_308)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_294),
.B(n_295),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_188),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_252),
.A2(n_228),
.B1(n_227),
.B2(n_178),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_306),
.B1(n_307),
.B2(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_263),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_263),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_242),
.B(n_181),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_301),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_179),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_209),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_302),
.B(n_316),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_R g304 ( 
.A(n_248),
.B(n_239),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g375 ( 
.A1(n_304),
.A2(n_324),
.B(n_332),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_241),
.B(n_235),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_274),
.A2(n_217),
.B1(n_204),
.B2(n_233),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_308),
.A2(n_339),
.B1(n_313),
.B2(n_326),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_309),
.A2(n_310),
.B1(n_315),
.B2(n_323),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_279),
.A2(n_200),
.B1(n_199),
.B2(n_190),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_312),
.Y(n_355)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_274),
.A2(n_206),
.B(n_202),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_314),
.A2(n_342),
.B(n_254),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_216),
.B1(n_203),
.B2(n_202),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_282),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_253),
.A2(n_7),
.B(n_15),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_317),
.A2(n_330),
.B(n_337),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_0),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_338),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_8),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_276),
.C(n_286),
.Y(n_349)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_257),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_7),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_325),
.B(n_328),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_269),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_258),
.B(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_246),
.A2(n_7),
.B(n_13),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_260),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_331),
.A2(n_339),
.B1(n_286),
.B2(n_276),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_R g332 ( 
.A(n_278),
.B(n_11),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_11),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_333),
.B(n_334),
.Y(n_386)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_335),
.A2(n_340),
.B1(n_244),
.B2(n_254),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_341),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_238),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_245),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_277),
.B(n_13),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_251),
.B(n_18),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_299),
.A2(n_251),
.B1(n_283),
.B2(n_250),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_344),
.A2(n_345),
.B1(n_347),
.B2(n_348),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_299),
.A2(n_283),
.B1(n_250),
.B2(n_271),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_303),
.A2(n_290),
.B1(n_287),
.B2(n_264),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_303),
.A2(n_290),
.B1(n_287),
.B2(n_264),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_301),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx3_ASAP7_75t_SL g357 ( 
.A(n_305),
.Y(n_357)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_367),
.B1(n_372),
.B2(n_383),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_285),
.C(n_237),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_366),
.C(n_349),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_305),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_362),
.Y(n_392)
);

AO22x1_ASAP7_75t_SL g362 ( 
.A1(n_304),
.A2(n_243),
.B1(n_240),
.B2(n_262),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_297),
.A2(n_278),
.B(n_262),
.C(n_255),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_374),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_240),
.C(n_243),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_336),
.A2(n_267),
.B1(n_272),
.B2(n_244),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_314),
.A2(n_265),
.B1(n_288),
.B2(n_272),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_368),
.A2(n_382),
.B1(n_364),
.B2(n_347),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_296),
.A2(n_265),
.B1(n_288),
.B2(n_255),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_314),
.A2(n_255),
.B(n_4),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_376),
.A2(n_325),
.B(n_317),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_294),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_380),
.Y(n_402)
);

OAI32xp33_ASAP7_75t_L g380 ( 
.A1(n_328),
.A2(n_5),
.A3(n_298),
.B1(n_300),
.B2(n_295),
.Y(n_380)
);

AOI22x1_ASAP7_75t_L g381 ( 
.A1(n_306),
.A2(n_5),
.B1(n_307),
.B2(n_318),
.Y(n_381)
);

AO21x2_ASAP7_75t_L g400 ( 
.A1(n_381),
.A2(n_376),
.B(n_352),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_309),
.A2(n_328),
.B1(n_310),
.B2(n_308),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_384),
.A2(n_332),
.B(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_354),
.A2(n_328),
.B1(n_323),
.B2(n_330),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_388),
.A2(n_399),
.B1(n_408),
.B2(n_416),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_324),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_389),
.A2(n_394),
.B(n_411),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_396),
.C(n_406),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_398),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_354),
.A2(n_315),
.B1(n_316),
.B2(n_342),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_400),
.A2(n_412),
.B1(n_420),
.B2(n_422),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_363),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_403),
.B(n_414),
.Y(n_430)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_319),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_293),
.C(n_311),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_344),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_374),
.A2(n_329),
.B1(n_327),
.B2(n_312),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_370),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_409),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_379),
.A2(n_333),
.B1(n_341),
.B2(n_322),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_321),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_377),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_363),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_378),
.A2(n_331),
.B1(n_335),
.B2(n_334),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_353),
.A2(n_340),
.B(n_335),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_417),
.A2(n_418),
.B(n_419),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_378),
.A2(n_375),
.B(n_370),
.Y(n_418)
);

AO22x1_ASAP7_75t_L g419 ( 
.A1(n_380),
.A2(n_362),
.B1(n_346),
.B2(n_382),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_359),
.A2(n_377),
.B1(n_372),
.B2(n_384),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_386),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_355),
.Y(n_444)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_424),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_345),
.Y(n_426)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_392),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_446),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_432),
.B(n_440),
.C(n_449),
.Y(n_486)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_422),
.A2(n_357),
.B1(n_361),
.B2(n_350),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_425),
.B1(n_390),
.B2(n_416),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_437),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_373),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_373),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_388),
.A2(n_364),
.B1(n_348),
.B2(n_368),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_441),
.A2(n_447),
.B1(n_450),
.B2(n_415),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_386),
.Y(n_443)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_444),
.A2(n_424),
.B1(n_356),
.B2(n_400),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_404),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_391),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_365),
.B(n_362),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_381),
.B1(n_362),
.B2(n_371),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_385),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_390),
.A2(n_381),
.B1(n_385),
.B2(n_355),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_452),
.Y(n_462)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_421),
.Y(n_453)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_453),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_407),
.B(n_356),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_417),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_430),
.B(n_418),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_458),
.B(n_459),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_429),
.B(n_413),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_474),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_456),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_477),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_464),
.A2(n_482),
.B1(n_441),
.B2(n_447),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_402),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_468),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_467),
.A2(n_426),
.B1(n_439),
.B2(n_450),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_402),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_437),
.B(n_397),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_469),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_435),
.B(n_394),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_443),
.Y(n_471)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_431),
.A2(n_400),
.B1(n_392),
.B2(n_415),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_472),
.A2(n_479),
.B1(n_445),
.B2(n_433),
.Y(n_495)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_473),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_389),
.Y(n_474)
);

XNOR2x1_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_389),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_440),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_452),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_431),
.A2(n_400),
.B1(n_419),
.B2(n_410),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_434),
.A2(n_393),
.B1(n_410),
.B2(n_419),
.Y(n_482)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_483),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_456),
.B(n_411),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_454),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_467),
.B1(n_480),
.B2(n_474),
.Y(n_525)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_490),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_491),
.A2(n_495),
.B1(n_461),
.B2(n_478),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_502),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_499),
.A2(n_478),
.B(n_477),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_454),
.C(n_436),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_509),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_428),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_483),
.Y(n_503)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_503),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_438),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_476),
.Y(n_526)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_506),
.Y(n_527)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_510),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_453),
.C(n_448),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_451),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_464),
.B1(n_482),
.B2(n_485),
.Y(n_511)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_511),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_499),
.A2(n_463),
.B(n_479),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_514),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_472),
.B(n_461),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_526),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_468),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_516),
.B(n_520),
.Y(n_536)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_517),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_465),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_491),
.A2(n_504),
.B1(n_494),
.B2(n_498),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_522),
.B(n_496),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_489),
.A2(n_460),
.B(n_480),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_523),
.A2(n_493),
.B(n_500),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_525),
.A2(n_528),
.B1(n_490),
.B2(n_488),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_487),
.A2(n_462),
.B1(n_442),
.B2(n_455),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_498),
.A2(n_455),
.B(n_452),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_528),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_505),
.C(n_509),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_531),
.Y(n_547)
);

OAI321xp33_ASAP7_75t_L g531 ( 
.A1(n_524),
.A2(n_510),
.A3(n_493),
.B1(n_503),
.B2(n_506),
.C(n_507),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_532),
.A2(n_534),
.B(n_517),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_502),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_545),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_511),
.B1(n_515),
.B2(n_529),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_497),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_543),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_496),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_492),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_544),
.B(n_522),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_519),
.B(n_492),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_535),
.A2(n_523),
.B(n_524),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_546),
.A2(n_555),
.B(n_556),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_538),
.A2(n_514),
.B1(n_512),
.B2(n_518),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_550),
.B(n_557),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_518),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_552),
.B(n_553),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_530),
.B(n_519),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_527),
.C(n_452),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_547),
.B(n_536),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_559),
.B(n_548),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_532),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_563),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_556),
.A2(n_541),
.B(n_527),
.Y(n_563)
);

AOI221xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_549),
.B1(n_551),
.B2(n_554),
.C(n_546),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_565),
.B(n_564),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_557),
.C(n_553),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_566),
.B(n_567),
.Y(n_570)
);

MAJx2_ASAP7_75t_L g572 ( 
.A(n_569),
.B(n_561),
.C(n_539),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_568),
.B(n_562),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_571),
.B(n_544),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_573),
.C(n_570),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_571),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_537),
.C(n_543),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_537),
.B(n_542),
.Y(n_577)
);


endmodule