module real_aes_8224_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_602;
wire n_552;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g458 ( .A1(n_0), .A2(n_159), .B(n_459), .C(n_462), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_1), .B(n_453), .Y(n_463) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g157 ( .A(n_3), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_4), .B(n_160), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_5), .A2(n_448), .B(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_6), .A2(n_182), .B(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_7), .A2(n_39), .B1(n_147), .B2(n_205), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_8), .A2(n_9), .B1(n_710), .B2(n_711), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_8), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_9), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_10), .B(n_182), .Y(n_190) );
AND2x6_ASAP7_75t_L g162 ( .A(n_11), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_12), .A2(n_162), .B(n_439), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_13), .B(n_40), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_13), .B(n_40), .Y(n_122) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
INVx1_ASAP7_75t_L g138 ( .A(n_15), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_16), .B(n_143), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_17), .B(n_160), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_18), .B(n_134), .Y(n_192) );
AO32x2_ASAP7_75t_L g243 ( .A1(n_19), .A2(n_133), .A3(n_176), .B1(n_182), .B2(n_244), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_20), .A2(n_30), .B1(n_124), .B2(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_20), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_21), .B(n_147), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_22), .B(n_134), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_23), .A2(n_56), .B1(n_147), .B2(n_205), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_24), .A2(n_81), .B1(n_143), .B2(n_147), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_25), .B(n_147), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_26), .A2(n_176), .B(n_439), .C(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_27), .A2(n_176), .B(n_439), .C(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_29), .B(n_178), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_30), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_30), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_31), .A2(n_448), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_32), .B(n_178), .Y(n_220) );
INVx2_ASAP7_75t_L g145 ( .A(n_33), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_34), .A2(n_445), .B(n_488), .C(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_35), .B(n_147), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_36), .B(n_178), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_37), .A2(n_103), .B1(n_116), .B2(n_739), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_38), .B(n_227), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_41), .B(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_42), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_43), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_44), .B(n_160), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_45), .B(n_448), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_46), .A2(n_445), .B(n_488), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_47), .B(n_147), .Y(n_185) );
INVx1_ASAP7_75t_L g460 ( .A(n_48), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_49), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_50), .A2(n_90), .B1(n_205), .B2(n_206), .Y(n_204) );
INVx1_ASAP7_75t_L g513 ( .A(n_51), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_52), .B(n_147), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_53), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_54), .B(n_448), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_55), .B(n_155), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_57), .A2(n_61), .B1(n_143), .B2(n_147), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_58), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_59), .B(n_147), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_60), .B(n_147), .Y(n_224) );
INVx1_ASAP7_75t_L g163 ( .A(n_62), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_63), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_64), .B(n_453), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_65), .A2(n_149), .B(n_155), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_66), .B(n_147), .Y(n_158) );
INVx1_ASAP7_75t_L g137 ( .A(n_67), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_68), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_69), .B(n_160), .Y(n_491) );
AO32x2_ASAP7_75t_L g202 ( .A1(n_70), .A2(n_176), .A3(n_182), .B1(n_203), .B2(n_208), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_71), .B(n_161), .Y(n_504) );
INVx1_ASAP7_75t_L g172 ( .A(n_72), .Y(n_172) );
INVx1_ASAP7_75t_L g215 ( .A(n_73), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_74), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_75), .B(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_76), .A2(n_439), .B(n_441), .C(n_445), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_77), .B(n_143), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_78), .Y(n_522) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_80), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_82), .B(n_205), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_83), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_84), .B(n_143), .Y(n_219) );
INVx2_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_86), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_87), .B(n_175), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_88), .B(n_143), .Y(n_186) );
INVx2_ASAP7_75t_L g112 ( .A(n_89), .Y(n_112) );
OR2x2_ASAP7_75t_L g120 ( .A(n_89), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g727 ( .A(n_89), .B(n_719), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_91), .A2(n_101), .B1(n_143), .B2(n_144), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_92), .B(n_448), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_93), .Y(n_490) );
INVxp67_ASAP7_75t_L g525 ( .A(n_94), .Y(n_525) );
XNOR2xp5_ASAP7_75t_L g728 ( .A(n_95), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_96), .B(n_143), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g442 ( .A(n_98), .Y(n_442) );
INVx1_ASAP7_75t_L g500 ( .A(n_99), .Y(n_500) );
AND2x2_ASAP7_75t_L g515 ( .A(n_100), .B(n_178), .Y(n_515) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g740 ( .A(n_106), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g121 ( .A(n_111), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g430 ( .A(n_112), .B(n_121), .Y(n_430) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_112), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO221x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_721), .B1(n_724), .B2(n_733), .C(n_735), .Y(n_116) );
OAI222xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_709), .B1(n_712), .B2(n_716), .C1(n_717), .C2(n_720), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B1(n_429), .B2(n_431), .Y(n_118) );
INVx2_ASAP7_75t_L g714 ( .A(n_119), .Y(n_714) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g719 ( .A(n_121), .Y(n_719) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_123), .A2(n_431), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_125), .A2(n_126), .B1(n_730), .B2(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR5x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_320), .C(n_378), .D(n_414), .E(n_421), .Y(n_126) );
NAND3xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_266), .C(n_290), .Y(n_127) );
AOI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_198), .B1(n_232), .B2(n_237), .C(n_247), .Y(n_128) );
OAI21xp5_ASAP7_75t_SL g400 ( .A1(n_129), .A2(n_401), .B(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_179), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_130), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
INVx2_ASAP7_75t_L g236 ( .A(n_131), .Y(n_236) );
AND2x2_ASAP7_75t_L g249 ( .A(n_131), .B(n_181), .Y(n_249) );
AND2x2_ASAP7_75t_L g303 ( .A(n_131), .B(n_180), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_131), .B(n_166), .Y(n_318) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_164), .Y(n_131) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_132), .A2(n_167), .B(n_177), .Y(n_166) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_133), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_135), .B(n_136), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_153), .B(n_162), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_146), .C(n_149), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_142), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_142), .A2(n_533), .B(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx3_ASAP7_75t_L g214 ( .A(n_147), .Y(n_214) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_147), .Y(n_444) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g205 ( .A(n_148), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
AND2x6_ASAP7_75t_L g439 ( .A(n_148), .B(n_440), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_L g441 ( .A1(n_149), .A2(n_442), .B(n_443), .C(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_150), .A2(n_218), .B(n_219), .Y(n_217) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g472 ( .A(n_151), .Y(n_472) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
INVx1_ASAP7_75t_L g227 ( .A(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g440 ( .A(n_152), .Y(n_440) );
AND2x2_ASAP7_75t_L g449 ( .A(n_152), .B(n_156), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_157), .B(n_158), .C(n_159), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g171 ( .A1(n_154), .A2(n_172), .B(n_173), .C(n_174), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_154), .A2(n_471), .B(n_473), .Y(n_470) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_159), .A2(n_188), .B(n_189), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_159), .A2(n_175), .B1(n_195), .B2(n_196), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_159), .A2(n_175), .B1(n_245), .B2(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_160), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_160), .A2(n_185), .B(n_186), .Y(n_184) );
O2A1O1Ixp5_ASAP7_75t_SL g213 ( .A1(n_160), .A2(n_214), .B(n_215), .C(n_216), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_160), .B(n_525), .Y(n_524) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_161), .A2(n_175), .B1(n_204), .B2(n_207), .Y(n_203) );
BUFx3_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_162), .A2(n_184), .B(n_187), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_162), .A2(n_213), .B(n_217), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_162), .A2(n_223), .B(n_228), .Y(n_222) );
INVx4_ASAP7_75t_SL g446 ( .A(n_162), .Y(n_446) );
AND2x4_ASAP7_75t_L g448 ( .A(n_162), .B(n_449), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_162), .B(n_449), .Y(n_501) );
AND2x2_ASAP7_75t_L g336 ( .A(n_165), .B(n_277), .Y(n_336) );
AND2x2_ASAP7_75t_L g369 ( .A(n_165), .B(n_181), .Y(n_369) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OR2x2_ASAP7_75t_L g276 ( .A(n_166), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g289 ( .A(n_166), .B(n_181), .Y(n_289) );
AND2x2_ASAP7_75t_L g296 ( .A(n_166), .B(n_277), .Y(n_296) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_166), .Y(n_305) );
AND2x2_ASAP7_75t_L g312 ( .A(n_166), .B(n_180), .Y(n_312) );
INVx1_ASAP7_75t_L g343 ( .A(n_166), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_176), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_174), .A2(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g461 ( .A(n_175), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g193 ( .A(n_176), .B(n_194), .C(n_197), .Y(n_193) );
INVx2_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_178), .A2(n_212), .B(n_220), .Y(n_211) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_178), .A2(n_222), .B(n_231), .Y(n_221) );
INVx1_ASAP7_75t_L g478 ( .A(n_178), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_178), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_178), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g319 ( .A(n_179), .Y(n_319) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_191), .Y(n_179) );
INVx2_ASAP7_75t_L g275 ( .A(n_180), .Y(n_275) );
AND2x2_ASAP7_75t_L g297 ( .A(n_180), .B(n_236), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_180), .B(n_343), .Y(n_348) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_181), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g420 ( .A(n_181), .B(n_384), .Y(n_420) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_190), .Y(n_181) );
INVx4_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_182), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_182), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g234 ( .A(n_191), .Y(n_234) );
INVx3_ASAP7_75t_L g335 ( .A(n_191), .Y(n_335) );
OR2x2_ASAP7_75t_L g365 ( .A(n_191), .B(n_366), .Y(n_365) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_191), .B(n_275), .Y(n_391) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_L g278 ( .A(n_192), .Y(n_278) );
AO21x1_ASAP7_75t_L g277 ( .A1(n_194), .A2(n_197), .B(n_278), .Y(n_277) );
AO21x2_ASAP7_75t_L g436 ( .A1(n_197), .A2(n_437), .B(n_450), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_197), .B(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g453 ( .A(n_197), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_197), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_197), .A2(n_499), .B(n_506), .Y(n_498) );
AOI33xp33_ASAP7_75t_L g411 ( .A1(n_198), .A2(n_249), .A3(n_263), .B1(n_335), .B2(n_412), .B3(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
OR2x2_ASAP7_75t_L g264 ( .A(n_200), .B(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_200), .B(n_261), .Y(n_323) );
OR2x2_ASAP7_75t_L g376 ( .A(n_200), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g302 ( .A(n_201), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g327 ( .A(n_201), .B(n_209), .Y(n_327) );
AND2x2_ASAP7_75t_L g394 ( .A(n_201), .B(n_239), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_201), .A2(n_294), .B(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
INVx1_ASAP7_75t_L g254 ( .A(n_202), .Y(n_254) );
AND2x2_ASAP7_75t_L g273 ( .A(n_202), .B(n_243), .Y(n_273) );
AND2x2_ASAP7_75t_L g322 ( .A(n_202), .B(n_242), .Y(n_322) );
INVx2_ASAP7_75t_L g462 ( .A(n_206), .Y(n_462) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_206), .Y(n_492) );
INVx1_ASAP7_75t_L g475 ( .A(n_208), .Y(n_475) );
INVx2_ASAP7_75t_SL g364 ( .A(n_209), .Y(n_364) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
INVx2_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
INVx1_ASAP7_75t_L g415 ( .A(n_210), .Y(n_415) );
AND2x2_ASAP7_75t_L g428 ( .A(n_210), .B(n_309), .Y(n_428) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g255 ( .A(n_211), .Y(n_255) );
OR2x2_ASAP7_75t_L g261 ( .A(n_211), .B(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
AND2x2_ASAP7_75t_L g256 ( .A(n_221), .B(n_242), .Y(n_256) );
INVx1_ASAP7_75t_L g262 ( .A(n_221), .Y(n_262) );
INVx1_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
AND2x2_ASAP7_75t_L g294 ( .A(n_221), .B(n_243), .Y(n_294) );
INVx2_ASAP7_75t_L g310 ( .A(n_221), .Y(n_310) );
AND2x2_ASAP7_75t_L g403 ( .A(n_221), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_221), .B(n_284), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx1_ASAP7_75t_L g287 ( .A(n_234), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_234), .B(n_318), .Y(n_384) );
INVx1_ASAP7_75t_SL g344 ( .A(n_235), .Y(n_344) );
INVx2_ASAP7_75t_L g265 ( .A(n_236), .Y(n_265) );
AND2x2_ASAP7_75t_L g334 ( .A(n_236), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g350 ( .A(n_236), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx1_ASAP7_75t_L g412 ( .A(n_238), .Y(n_412) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g267 ( .A(n_240), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g370 ( .A(n_240), .B(n_360), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_240), .A2(n_381), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x2_ASAP7_75t_L g283 ( .A(n_241), .B(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g308 ( .A(n_241), .Y(n_308) );
INVx1_ASAP7_75t_L g332 ( .A(n_241), .Y(n_332) );
OR2x2_ASAP7_75t_L g396 ( .A(n_242), .B(n_255), .Y(n_396) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_242), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g309 ( .A(n_243), .B(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g316 ( .A(n_243), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B1(n_257), .B2(n_259), .Y(n_247) );
OR2x2_ASAP7_75t_L g326 ( .A(n_248), .B(n_276), .Y(n_326) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_249), .A2(n_368), .B1(n_370), .B2(n_371), .C1(n_372), .C2(n_375), .Y(n_367) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_256), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g314 ( .A(n_253), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_255), .B(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_255), .Y(n_339) );
AND2x2_ASAP7_75t_L g387 ( .A(n_255), .B(n_256), .Y(n_387) );
INVx1_ASAP7_75t_L g405 ( .A(n_255), .Y(n_405) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g371 ( .A(n_258), .B(n_297), .Y(n_371) );
AND2x2_ASAP7_75t_L g413 ( .A(n_258), .B(n_289), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_260), .B(n_308), .Y(n_395) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_261), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g288 ( .A(n_265), .B(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g356 ( .A(n_265), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_274), .C(n_279), .Y(n_266) );
INVxp67_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_268), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_268), .B(n_315), .Y(n_410) );
BUFx3_ASAP7_75t_L g374 ( .A(n_269), .Y(n_374) );
INVx1_ASAP7_75t_L g281 ( .A(n_270), .Y(n_281) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g300 ( .A(n_272), .B(n_294), .Y(n_300) );
INVx1_ASAP7_75t_SL g340 ( .A(n_273), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g330 ( .A(n_275), .Y(n_330) );
AND2x2_ASAP7_75t_L g353 ( .A(n_275), .B(n_336), .Y(n_353) );
INVx1_ASAP7_75t_SL g324 ( .A(n_276), .Y(n_324) );
INVx1_ASAP7_75t_L g351 ( .A(n_277), .Y(n_351) );
AOI31xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .A3(n_282), .B(n_285), .Y(n_279) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g372 ( .A(n_283), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g346 ( .A(n_284), .Y(n_346) );
BUFx2_ASAP7_75t_L g360 ( .A(n_284), .Y(n_360) );
AND2x2_ASAP7_75t_L g388 ( .A(n_284), .B(n_309), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g361 ( .A(n_288), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_289), .B(n_356), .Y(n_402) );
AND2x2_ASAP7_75t_L g409 ( .A(n_289), .B(n_335), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B(n_298), .C(n_313), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_295), .A2(n_322), .B1(n_323), .B2(n_324), .C(n_325), .Y(n_321) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g329 ( .A(n_296), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g366 ( .A(n_297), .Y(n_366) );
OAI32xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .A3(n_304), .B1(n_306), .B2(n_311), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_300), .A2(n_353), .B(n_354), .C(n_357), .Y(n_352) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
OAI21xp5_ASAP7_75t_SL g416 ( .A1(n_308), .A2(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g377 ( .A(n_309), .Y(n_377) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_315), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g363 ( .A(n_315), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g380 ( .A(n_317), .Y(n_380) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND4xp25_ASAP7_75t_SL g320 ( .A(n_321), .B(n_333), .C(n_352), .D(n_367), .Y(n_320) );
AND2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g381 ( .A(n_322), .B(n_374), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_324), .B(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_328), .B2(n_331), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_326), .A2(n_377), .B1(n_408), .B2(n_410), .Y(n_407) );
O2A1O1Ixp33_ASAP7_75t_L g414 ( .A1(n_326), .A2(n_415), .B(n_416), .C(n_419), .Y(n_414) );
INVx2_ASAP7_75t_L g385 ( .A(n_327), .Y(n_385) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g379 ( .A1(n_329), .A2(n_363), .B1(n_380), .B2(n_381), .C1(n_382), .C2(n_385), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_337), .C(n_341), .Y(n_333) );
INVx1_ASAP7_75t_L g399 ( .A(n_334), .Y(n_399) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_338), .A2(n_342), .B1(n_345), .B2(n_347), .Y(n_341) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g368 ( .A(n_350), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g426 ( .A(n_353), .Y(n_426) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B1(n_362), .B2(n_365), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_360), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
INVx1_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_371), .Y(n_425) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND5xp2_ASAP7_75t_L g378 ( .A(n_379), .B(n_386), .C(n_400), .D(n_406), .E(n_411), .Y(n_378) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_389), .C(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI31xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .A3(n_396), .B(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI222xp33_ASAP7_75t_L g421 ( .A1(n_408), .A2(n_410), .B1(n_422), .B2(n_425), .C1(n_426), .C2(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g715 ( .A(n_429), .Y(n_715) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR3x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_617), .C(n_666), .Y(n_431) );
NAND5xp2_ASAP7_75t_L g432 ( .A(n_433), .B(n_551), .C(n_580), .D(n_588), .E(n_603), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_479), .B(n_495), .C(n_535), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_464), .Y(n_434) );
AND2x2_ASAP7_75t_L g546 ( .A(n_435), .B(n_543), .Y(n_546) );
AND2x2_ASAP7_75t_L g579 ( .A(n_435), .B(n_465), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_435), .B(n_483), .Y(n_672) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_452), .Y(n_435) );
INVx2_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
BUFx2_ASAP7_75t_L g646 ( .A(n_436), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_447), .Y(n_437) );
INVx5_ASAP7_75t_L g457 ( .A(n_439), .Y(n_457) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_SL g455 ( .A1(n_446), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_446), .A2(n_457), .B(n_522), .C(n_523), .Y(n_521) );
BUFx2_ASAP7_75t_L g468 ( .A(n_448), .Y(n_468) );
AND2x2_ASAP7_75t_L g464 ( .A(n_452), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g544 ( .A(n_452), .Y(n_544) );
AND2x2_ASAP7_75t_L g630 ( .A(n_452), .B(n_543), .Y(n_630) );
AND2x2_ASAP7_75t_L g685 ( .A(n_452), .B(n_482), .Y(n_685) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_463), .Y(n_452) );
INVx2_ASAP7_75t_L g488 ( .A(n_457), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g602 ( .A(n_464), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_464), .B(n_483), .Y(n_649) );
INVx5_ASAP7_75t_L g543 ( .A(n_465), .Y(n_543) );
AND2x4_ASAP7_75t_L g564 ( .A(n_465), .B(n_544), .Y(n_564) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_465), .Y(n_586) );
AND2x2_ASAP7_75t_L g661 ( .A(n_465), .B(n_646), .Y(n_661) );
AND2x2_ASAP7_75t_L g664 ( .A(n_465), .B(n_484), .Y(n_664) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
AOI21xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_469), .B(n_475), .Y(n_466) );
INVx2_ASAP7_75t_L g474 ( .A(n_472), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_474), .A2(n_490), .B(n_491), .C(n_492), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_474), .A2(n_492), .B(n_513), .C(n_514), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_479), .B(n_544), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_479), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
AND2x2_ASAP7_75t_L g569 ( .A(n_481), .B(n_544), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_481), .B(n_484), .Y(n_587) );
INVx1_ASAP7_75t_L g607 ( .A(n_481), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_481), .B(n_543), .Y(n_652) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_481), .Y(n_694) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_482), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_483), .B(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_483), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_483), .A2(n_539), .B(n_600), .C(n_602), .Y(n_599) );
AND2x2_ASAP7_75t_L g606 ( .A(n_483), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g615 ( .A(n_483), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g619 ( .A(n_483), .B(n_543), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_483), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g634 ( .A(n_483), .B(n_544), .Y(n_634) );
AND2x2_ASAP7_75t_L g684 ( .A(n_483), .B(n_685), .Y(n_684) );
INVx5_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g548 ( .A(n_484), .Y(n_548) );
AND2x2_ASAP7_75t_L g589 ( .A(n_484), .B(n_542), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_484), .B(n_576), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_484), .B(n_630), .Y(n_648) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_516), .Y(n_495) );
INVx1_ASAP7_75t_L g537 ( .A(n_496), .Y(n_537) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
OR2x2_ASAP7_75t_L g539 ( .A(n_497), .B(n_508), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_497), .B(n_546), .C(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_497), .B(n_518), .Y(n_556) );
OR2x2_ASAP7_75t_L g571 ( .A(n_497), .B(n_559), .Y(n_571) );
AND2x2_ASAP7_75t_L g577 ( .A(n_497), .B(n_527), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_497), .B(n_708), .Y(n_707) );
INVx5_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_498), .B(n_518), .Y(n_574) );
AND2x2_ASAP7_75t_L g613 ( .A(n_498), .B(n_528), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_498), .B(n_527), .Y(n_641) );
OR2x2_ASAP7_75t_L g644 ( .A(n_498), .B(n_527), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_502), .Y(n_499) );
INVx5_ASAP7_75t_SL g559 ( .A(n_508), .Y(n_559) );
OR2x2_ASAP7_75t_L g565 ( .A(n_508), .B(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g581 ( .A(n_508), .B(n_582), .Y(n_581) );
AOI321xp33_ASAP7_75t_L g588 ( .A1(n_508), .A2(n_589), .A3(n_590), .B1(n_591), .B2(n_597), .C(n_599), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_508), .B(n_516), .Y(n_598) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_508), .Y(n_611) );
OR2x2_ASAP7_75t_L g658 ( .A(n_508), .B(n_556), .Y(n_658) );
AND2x2_ASAP7_75t_L g680 ( .A(n_508), .B(n_577), .Y(n_680) );
AND2x2_ASAP7_75t_L g699 ( .A(n_508), .B(n_518), .Y(n_699) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_518), .B(n_527), .Y(n_540) );
AND2x2_ASAP7_75t_L g549 ( .A(n_518), .B(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g576 ( .A(n_518), .Y(n_576) );
AND2x2_ASAP7_75t_L g582 ( .A(n_518), .B(n_577), .Y(n_582) );
INVxp67_ASAP7_75t_L g612 ( .A(n_518), .Y(n_612) );
OR2x2_ASAP7_75t_L g654 ( .A(n_518), .B(n_559), .Y(n_654) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_526), .Y(n_518) );
OR2x2_ASAP7_75t_L g536 ( .A(n_527), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_SL g550 ( .A(n_527), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_527), .B(n_539), .Y(n_583) );
AND2x2_ASAP7_75t_L g632 ( .A(n_527), .B(n_576), .Y(n_632) );
AND2x2_ASAP7_75t_L g670 ( .A(n_527), .B(n_559), .Y(n_670) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_528), .B(n_559), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_538), .B(n_541), .C(n_545), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_536), .A2(n_538), .B1(n_663), .B2(n_665), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_538), .A2(n_561), .B1(n_616), .B2(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_SL g690 ( .A(n_539), .Y(n_690) );
INVx1_ASAP7_75t_SL g590 ( .A(n_540), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_542), .B(n_562), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g603 ( .A1(n_542), .A2(n_583), .B1(n_590), .B2(n_604), .C1(n_608), .C2(n_614), .Y(n_603) );
AND2x2_ASAP7_75t_L g693 ( .A(n_542), .B(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g568 ( .A(n_543), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_543), .B(n_563), .Y(n_638) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_543), .Y(n_675) );
AND2x2_ASAP7_75t_L g678 ( .A(n_543), .B(n_587), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_543), .B(n_694), .Y(n_704) );
INVx1_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_544), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g686 ( .A1(n_546), .A2(n_687), .B(n_688), .C(n_691), .Y(n_686) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_548), .B(n_610), .C(n_613), .Y(n_609) );
OR2x2_ASAP7_75t_L g637 ( .A(n_548), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_548), .B(n_564), .Y(n_665) );
OR2x2_ASAP7_75t_L g570 ( .A(n_550), .B(n_571), .Y(n_570) );
AOI211xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_554), .B(n_560), .C(n_572), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_553), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g659 ( .A(n_554), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_555), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g573 ( .A(n_558), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_559), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g627 ( .A(n_559), .B(n_577), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_559), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_559), .B(n_576), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_565), .B1(n_566), .B2(n_570), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_562), .B(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_564), .B(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_SL g628 ( .A1(n_565), .A2(n_629), .B1(n_631), .B2(n_633), .C(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g683 ( .A(n_568), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g696 ( .A(n_568), .B(n_685), .Y(n_696) );
INVx1_ASAP7_75t_L g616 ( .A(n_569), .Y(n_616) );
INVx1_ASAP7_75t_L g687 ( .A(n_570), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_571), .A2(n_654), .B(n_677), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_578), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_583), .B(n_584), .Y(n_580) );
INVx1_ASAP7_75t_L g620 ( .A(n_581), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_582), .A2(n_668), .B1(n_671), .B2(n_673), .C(n_676), .Y(n_667) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_590), .A2(n_680), .B1(n_681), .B2(n_683), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g656 ( .A(n_592), .Y(n_656) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp67_ASAP7_75t_SL g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g660 ( .A(n_596), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g625 ( .A(n_601), .Y(n_625) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_606), .B(n_630), .Y(n_682) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_612), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g698 ( .A(n_613), .B(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_L g705 ( .A(n_613), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI211xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_620), .B(n_621), .C(n_655), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI211xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B(n_628), .C(n_647), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g708 ( .A(n_632), .Y(n_708) );
AND2x2_ASAP7_75t_L g645 ( .A(n_634), .B(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .B1(n_643), .B2(n_645), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
OR2x2_ASAP7_75t_L g653 ( .A(n_641), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g706 ( .A(n_642), .Y(n_706) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI31xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .A3(n_650), .B(n_653), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B(n_659), .C(n_662), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
CKINVDCx16_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
NAND5xp2_ASAP7_75t_L g666 ( .A(n_667), .B(n_679), .C(n_686), .D(n_700), .E(n_703), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_678), .A2(n_704), .B1(n_705), .B2(n_707), .Y(n_703) );
INVx1_ASAP7_75t_SL g702 ( .A(n_680), .Y(n_702) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B(n_697), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g716 ( .A(n_709), .Y(n_716) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_SL g734 ( .A(n_722), .Y(n_734) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g738 ( .A(n_727), .Y(n_738) );
INVx1_ASAP7_75t_L g732 ( .A(n_730), .Y(n_732) );
BUFx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
endmodule