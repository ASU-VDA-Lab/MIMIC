module fake_jpeg_11509_n_293 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_293);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_9),
.B(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_56),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_61),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_2),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_2),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_36),
.B1(n_22),
.B2(n_34),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_98),
.C(n_52),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_4),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_34),
.B1(n_41),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_85),
.B1(n_93),
.B2(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_37),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_91),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_22),
.B1(n_25),
.B2(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_25),
.B1(n_40),
.B2(n_39),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_25),
.B1(n_40),
.B2(n_39),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_34),
.B1(n_41),
.B2(n_28),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_41),
.B1(n_37),
.B2(n_31),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_48),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_26),
.B1(n_30),
.B2(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_23),
.B1(n_33),
.B2(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_33),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_4),
.Y(n_116)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_52),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_130),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_68),
.B1(n_49),
.B2(n_67),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_95),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_56),
.B1(n_65),
.B2(n_7),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_136),
.Y(n_163)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_137),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_73),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_138),
.Y(n_153)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_7),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_13),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_71),
.B(n_8),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_75),
.B(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_9),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_11),
.Y(n_172)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

CKINVDCx10_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_147),
.B1(n_174),
.B2(n_99),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_71),
.B1(n_96),
.B2(n_99),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_172),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_100),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_170),
.Y(n_178)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_83),
.B1(n_77),
.B2(n_104),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_134),
.B1(n_123),
.B2(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_83),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_127),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_120),
.A2(n_97),
.B(n_96),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_82),
.B(n_112),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_111),
.B(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_136),
.B1(n_117),
.B2(n_128),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_180),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_118),
.C(n_115),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_181),
.C(n_90),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_167),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_184),
.B(n_186),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_139),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_137),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_190),
.Y(n_218)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_115),
.B1(n_116),
.B2(n_94),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_194),
.B1(n_171),
.B2(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_198),
.B(n_90),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_152),
.B(n_82),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_132),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_145),
.A2(n_110),
.B1(n_140),
.B2(n_123),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_199),
.B1(n_171),
.B2(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_144),
.B1(n_141),
.B2(n_125),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_126),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_135),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_160),
.B1(n_170),
.B2(n_163),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_207),
.B1(n_208),
.B2(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_185),
.C(n_183),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_165),
.B1(n_149),
.B2(n_162),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_162),
.B1(n_165),
.B2(n_149),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_148),
.A3(n_154),
.B1(n_156),
.B2(n_158),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_175),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_175),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_228),
.C(n_219),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_176),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_179),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_235),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_218),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_238),
.B(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_175),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_207),
.B1(n_215),
.B2(n_188),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_182),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_185),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_252),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_248),
.C(n_251),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_212),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_211),
.B1(n_213),
.B2(n_203),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_253),
.B1(n_226),
.B2(n_243),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_226),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_211),
.C(n_209),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_215),
.B1(n_216),
.B2(n_221),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_182),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_238),
.C(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_240),
.B(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_259),
.Y(n_270)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_240),
.B(n_237),
.C(n_233),
.D(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_265),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_251),
.C(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_271),
.C(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_254),
.C(n_250),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_256),
.B(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_246),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_230),
.CI(n_259),
.CON(n_277),
.SN(n_277)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_229),
.B(n_262),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_275),
.B1(n_272),
.B2(n_268),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_283),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_269),
.B(n_227),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_272),
.B1(n_221),
.B2(n_216),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_200),
.B1(n_177),
.B2(n_235),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.C(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_286),
.B(n_177),
.Y(n_288)
);

AOI221xp5_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_180),
.B1(n_191),
.B2(n_193),
.C(n_198),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_289),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_290),
.B(n_286),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_11),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_292),
.B(n_12),
.CI(n_286),
.CON(n_293),
.SN(n_293)
);


endmodule