module fake_jpeg_27079_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_32),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_57),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_16),
.B1(n_18),
.B2(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_53),
.B(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_24),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_40),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_26),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_30),
.B1(n_23),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_75),
.B1(n_47),
.B2(n_36),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_18),
.B1(n_26),
.B2(n_17),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_16),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_37),
.B(n_36),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_46),
.B1(n_21),
.B2(n_30),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_86),
.B1(n_56),
.B2(n_37),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_79),
.B1(n_38),
.B2(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_38),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_104),
.B(n_101),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_38),
.B(n_35),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_76),
.B(n_67),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_79),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_69),
.B(n_88),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_84),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_22),
.B(n_19),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_37),
.B1(n_36),
.B2(n_56),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_36),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_77),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_63),
.B1(n_58),
.B2(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_68),
.Y(n_124)
);

OAI221xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_108),
.B1(n_22),
.B2(n_0),
.C(n_3),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_74),
.B1(n_86),
.B2(n_78),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_137),
.B1(n_90),
.B2(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_122),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

XOR2x1_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_87),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_127),
.B(n_102),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_130),
.B1(n_103),
.B2(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_126),
.B1(n_133),
.B2(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_60),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_66),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_129),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_69),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_93),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_97),
.B1(n_102),
.B2(n_90),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_96),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_134),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_92),
.B(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_19),
.B1(n_22),
.B2(n_0),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_89),
.B(n_19),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_0),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_115),
.B1(n_137),
.B2(n_135),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_133),
.B1(n_121),
.B2(n_124),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_156),
.B(n_135),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_90),
.B(n_112),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_154),
.B(n_2),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_106),
.C(n_89),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_152),
.C(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_106),
.C(n_105),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_92),
.B(n_96),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_5),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_8),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_7),
.C(n_1),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_7),
.C(n_1),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_10),
.C(n_2),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_169),
.B(n_175),
.Y(n_189)
);

OAI322xp33_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_128),
.A3(n_136),
.B1(n_123),
.B2(n_138),
.C1(n_122),
.C2(n_117),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_151),
.B1(n_157),
.B2(n_140),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_11),
.C(n_1),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_173),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_172),
.B1(n_160),
.B2(n_149),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_171),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_117),
.B(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_174),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_177),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_5),
.C(n_6),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_173),
.C(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_184),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_141),
.A3(n_146),
.B1(n_151),
.B2(n_153),
.C1(n_148),
.C2(n_157),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_145),
.C(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_188),
.Y(n_199)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_148),
.C(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_167),
.B1(n_139),
.B2(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_191),
.A2(n_175),
.B(n_176),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_191),
.B1(n_190),
.B2(n_184),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_198),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_197),
.B(n_182),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_189),
.A2(n_162),
.B(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_202),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_139),
.B(n_162),
.Y(n_197)
);

INVxp33_ASAP7_75t_SL g200 ( 
.A(n_181),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_200),
.A2(n_189),
.B1(n_181),
.B2(n_187),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_179),
.B1(n_190),
.B2(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_209),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_212),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_211),
.B(n_12),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_185),
.B1(n_183),
.B2(n_178),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_193),
.B1(n_195),
.B2(n_13),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_159),
.B1(n_177),
.B2(n_11),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_8),
.C(n_10),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_215),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_10),
.B(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_211),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_205),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_220),
.A2(n_221),
.B1(n_218),
.B2(n_212),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_222),
.B1(n_205),
.B2(n_210),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_217),
.B(n_213),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_207),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_227),
.B(n_223),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_15),
.Y(n_230)
);


endmodule