module fake_jpeg_28616_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_0),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_61),
.B1(n_52),
.B2(n_50),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_93),
.B1(n_58),
.B2(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_49),
.B1(n_55),
.B2(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_70),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_58),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_58),
.B1(n_54),
.B2(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_108),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_62),
.B(n_66),
.C(n_65),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_113),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_111),
.Y(n_118)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_96),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_64),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_2),
.B(n_3),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_3),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_132),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_55),
.C(n_49),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_29),
.C(n_47),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_131),
.B1(n_9),
.B2(n_11),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_8),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_7),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_142),
.B(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_138),
.C(n_146),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_28),
.C(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_141),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_118),
.B(n_127),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_148),
.B(n_124),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_32),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_33),
.C(n_12),
.Y(n_147)
);

BUFx10_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_126),
.A3(n_9),
.B1(n_16),
.B2(n_20),
.C1(n_21),
.C2(n_23),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_119),
.B(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_149),
.B(n_143),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_140),
.B(n_137),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_14),
.C(n_26),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_27),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_151),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_151),
.B1(n_162),
.B2(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_156),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_148),
.A3(n_37),
.B1(n_39),
.B2(n_40),
.C1(n_35),
.C2(n_41),
.Y(n_167)
);


endmodule