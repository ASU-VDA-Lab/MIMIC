module fake_jpeg_11722_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_3),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_26),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_0),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_91),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_98),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_77),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_76),
.B(n_61),
.C(n_69),
.Y(n_98)
);

CKINVDCx9p33_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_69),
.B1(n_75),
.B2(n_64),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_106),
.C(n_5),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_67),
.B1(n_71),
.B2(n_60),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_66),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_49),
.B1(n_73),
.B2(n_72),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_111),
.B1(n_115),
.B2(n_110),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OR2x4_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_58),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_71),
.B1(n_67),
.B2(n_68),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_28),
.B1(n_46),
.B2(n_45),
.Y(n_132)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_65),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_59),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_70),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_51),
.B1(n_57),
.B2(n_29),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_129),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_63),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_137),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_134),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_61),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_31),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_8),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_9),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_155),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_10),
.CI(n_17),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_41),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_159),
.Y(n_168)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_32),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_133),
.B1(n_126),
.B2(n_128),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_148),
.B1(n_160),
.B2(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_126),
.C(n_162),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_153),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_176),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_171),
.B1(n_163),
.B2(n_168),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_179),
.Y(n_180)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_177),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_154),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_166),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_175),
.Y(n_186)
);


endmodule