module real_jpeg_14598_n_16 (n_5, n_4, n_8, n_0, n_12, n_413, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_412, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_413;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_412;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_0),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_3),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_3),
.B(n_32),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_3),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_3),
.B(n_52),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_3),
.B(n_40),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_5),
.B(n_32),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_110),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_5),
.B(n_29),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_5),
.B(n_40),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_5),
.B(n_45),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_6),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_29),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_6),
.B(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_32),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_6),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_52),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_6),
.B(n_40),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_6),
.B(n_45),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_7),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_7),
.B(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_7),
.B(n_40),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_7),
.B(n_110),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_7),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_7),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_52),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_10),
.B(n_26),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_10),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_40),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_12),
.B(n_110),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_12),
.B(n_115),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_12),
.B(n_26),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_12),
.B(n_29),
.Y(n_327)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_13),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_13),
.B(n_115),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_13),
.B(n_32),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_13),
.B(n_26),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_52),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_40),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_110),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_14),
.B(n_115),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_14),
.B(n_26),
.Y(n_248)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_79),
.B(n_344),
.C(n_408),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_89),
.B(n_407),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_21),
.B(n_77),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.C(n_64),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_22),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.C(n_54),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_23),
.B(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_37),
.C(n_41),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_25),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_56),
.C(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_25),
.A2(n_62),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_25),
.B(n_233),
.C(n_234),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_25),
.A2(n_31),
.B1(n_62),
.B2(n_182),
.Y(n_385)
);

INVx5_ASAP7_75t_SL g124 ( 
.A(n_26),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_28),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_28),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_28),
.B(n_273),
.C(n_276),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_28),
.A2(n_277),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_30),
.B(n_38),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_31),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_31),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_31),
.B(n_178),
.C(n_180),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_31),
.A2(n_136),
.B1(n_137),
.B2(n_182),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_31),
.B(n_136),
.C(n_248),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_33),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_33),
.B(n_50),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_33),
.B(n_43),
.Y(n_252)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_38),
.B(n_109),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_43),
.B(n_227),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_44),
.B(n_157),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_44),
.B(n_111),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_44),
.B(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_47),
.A2(n_54),
.B1(n_55),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_47),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.C(n_51),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_48),
.B(n_51),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_49),
.A2(n_87),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

NOR3xp33_ASAP7_75t_L g408 ( 
.A(n_49),
.B(n_68),
.C(n_85),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_52),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_56),
.A2(n_57),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_57),
.B(n_117),
.C(n_233),
.Y(n_340)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_66),
.C(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_60),
.A2(n_61),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_61),
.B(n_246),
.C(n_248),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_63),
.B(n_64),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_72),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_74),
.C(n_75),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_66),
.A2(n_70),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_66),
.B(n_353),
.C(n_354),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_69),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_68),
.A2(n_69),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_69),
.B(n_287),
.C(n_289),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_88),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_85),
.A2(n_86),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_86),
.B(n_309),
.C(n_312),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_402),
.B(n_406),
.Y(n_89)
);

OAI321xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_370),
.A3(n_390),
.B1(n_400),
.B2(n_401),
.C(n_412),
.Y(n_90)
);

AOI321xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_298),
.A3(n_330),
.B1(n_364),
.B2(n_369),
.C(n_413),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_237),
.C(n_293),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_205),
.B(n_236),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_172),
.B(n_204),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_141),
.B(n_171),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_118),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_97),
.B(n_118),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_112),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_121),
.B1(n_122),
.B2(n_130),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_98),
.B(n_168),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.CI(n_101),
.CON(n_98),
.SN(n_98)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_102),
.A2(n_103),
.B1(n_112),
.B2(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_105),
.B(n_157),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_107),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_109),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_116),
.A2(n_117),
.B1(n_186),
.B2(n_187),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_116),
.A2(n_117),
.B1(n_232),
.B2(n_233),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_117),
.B(n_187),
.C(n_290),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_131),
.B2(n_140),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_130),
.C(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_126),
.C(n_129),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_134),
.C(n_135),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_136),
.A2(n_137),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_136),
.A2(n_137),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_136),
.B(n_344),
.C(n_346),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_138),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_137),
.B(n_325),
.C(n_327),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_138),
.A2(n_139),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_138),
.B(n_260),
.C(n_263),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_165),
.B(n_170),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_154),
.B(n_164),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_152),
.C(n_153),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_159),
.B(n_163),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_167),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_174),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_190),
.B2(n_191),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_192),
.C(n_203),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_184),
.C(n_185),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_188),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_202),
.B2(n_203),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_201),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_198),
.C(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_197),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_207),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_223),
.B2(n_235),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_222),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_210),
.B(n_222),
.C(n_235),
.Y(n_294)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_219),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_220),
.C(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_214),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.CI(n_217),
.CON(n_214),
.SN(n_214)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_216),
.C(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_223),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.CI(n_230),
.CON(n_223),
.SN(n_223)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_225),
.C(n_230),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_228),
.B(n_229),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_229),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g365 ( 
.A1(n_238),
.A2(n_366),
.B(n_367),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_269),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_239),
.B(n_269),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_257),
.C(n_268),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_256),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_249),
.C(n_256),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_245),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_247),
.A2(n_248),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_253),
.C(n_255),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_257),
.A2(n_258),
.B1(n_268),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_265),
.C(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_262),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_292),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_281),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_281),
.C(n_292),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_279),
.C(n_280),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_294),
.B(n_295),
.Y(n_366)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_299),
.A2(n_365),
.B(n_368),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_300),
.B(n_301),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_329),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_304),
.C(n_329),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_321),
.B2(n_322),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_323),
.C(n_324),
.Y(n_363)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_315),
.C(n_320),
.Y(n_336)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_327),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_332),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_363),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_348),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_348),
.C(n_363),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_339),
.C(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_346),
.Y(n_339)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_340),
.Y(n_346)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_355),
.B2(n_356),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_357),
.C(n_362),
.Y(n_373)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_352),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_361),
.B2(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_371),
.B(n_372),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_391),
.Y(n_401)
);

FAx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.CI(n_389),
.CON(n_372),
.SN(n_372)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_379),
.C(n_382),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_380),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_387),
.C(n_388),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_399),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_397),
.B2(n_398),
.Y(n_392)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_398),
.C(n_399),
.Y(n_403)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_404),
.Y(n_406)
);


endmodule