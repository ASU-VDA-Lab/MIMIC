module real_aes_5677_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_1077, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_1076, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_1077;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_1076;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_635;
wire n_792;
wire n_673;
wire n_386;
wire n_503;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_320;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_1053;
wire n_1049;
wire n_636;
wire n_466;
wire n_559;
wire n_976;
wire n_906;
wire n_477;
wire n_872;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_1031;
wire n_432;
wire n_880;
wire n_1037;
wire n_1008;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_1041;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_288;
wire n_1073;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_354;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1051;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_1071;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_0), .A2(n_19), .B1(n_389), .B2(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_1), .A2(n_52), .B1(n_795), .B2(n_799), .Y(n_802) );
AOI21xp33_ASAP7_75t_L g1064 ( .A1(n_2), .A2(n_402), .B(n_1065), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_3), .Y(n_292) );
AND2x4_ASAP7_75t_L g789 ( .A(n_3), .B(n_790), .Y(n_789) );
AND2x4_ASAP7_75t_L g798 ( .A(n_3), .B(n_274), .Y(n_798) );
INVx1_ASAP7_75t_L g544 ( .A(n_4), .Y(n_544) );
INVx1_ASAP7_75t_L g392 ( .A(n_5), .Y(n_392) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_6), .B(n_442), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_7), .A2(n_62), .B1(n_431), .B2(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_8), .B(n_471), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_9), .A2(n_120), .B1(n_499), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_10), .A2(n_94), .B1(n_471), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_11), .A2(n_217), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI21xp33_ASAP7_75t_SL g550 ( .A1(n_12), .A2(n_551), .B(n_552), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_13), .A2(n_84), .B1(n_788), .B2(n_792), .Y(n_801) );
INVx1_ASAP7_75t_L g453 ( .A(n_14), .Y(n_453) );
INVx1_ASAP7_75t_L g300 ( .A(n_15), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_16), .A2(n_232), .B1(n_354), .B2(n_358), .Y(n_1057) );
INVx1_ASAP7_75t_L g825 ( .A(n_17), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_18), .A2(n_192), .B1(n_371), .B2(n_372), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_20), .A2(n_139), .B1(n_389), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_21), .A2(n_56), .B1(n_389), .B2(n_406), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_22), .A2(n_178), .B1(n_415), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_23), .A2(n_121), .B1(n_415), .B2(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_24), .A2(n_243), .B1(n_406), .B2(n_459), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_25), .A2(n_81), .B1(n_830), .B2(n_842), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_26), .A2(n_111), .B1(n_420), .B2(n_422), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_27), .A2(n_69), .B1(n_341), .B2(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g487 ( .A(n_28), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_29), .A2(n_255), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_30), .A2(n_107), .B1(n_305), .B2(n_375), .Y(n_735) );
INVx1_ASAP7_75t_L g467 ( .A(n_31), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_32), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g895 ( .A(n_33), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_34), .B(n_644), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_35), .A2(n_72), .B1(n_366), .B2(n_369), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_36), .B(n_221), .Y(n_290) );
INVx1_ASAP7_75t_L g324 ( .A(n_36), .Y(n_324) );
INVxp67_ASAP7_75t_L g351 ( .A(n_36), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_37), .A2(n_95), .B1(n_821), .B2(n_835), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_38), .A2(n_131), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_39), .A2(n_75), .B1(n_496), .B2(n_611), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_40), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_41), .A2(n_102), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_42), .A2(n_640), .B1(n_657), .B2(n_658), .Y(n_639) );
INVxp67_ASAP7_75t_L g658 ( .A(n_42), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_43), .A2(n_88), .B1(n_447), .B2(n_564), .Y(n_1043) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_44), .B(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_45), .A2(n_92), .B1(n_664), .B2(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_46), .B(n_396), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_47), .A2(n_114), .B1(n_354), .B2(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_48), .B(n_309), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_49), .A2(n_182), .B1(n_564), .B2(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_50), .A2(n_244), .B1(n_328), .B2(n_344), .Y(n_1067) );
INVx1_ASAP7_75t_SL g626 ( .A(n_51), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_53), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_54), .A2(n_280), .B1(n_827), .B2(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_55), .A2(n_198), .B1(n_524), .B2(n_526), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_57), .A2(n_91), .B1(n_332), .B2(n_341), .Y(n_736) );
INVxp67_ASAP7_75t_R g828 ( .A(n_58), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_59), .A2(n_222), .B1(n_406), .B2(n_506), .Y(n_558) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_60), .B(n_304), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_61), .A2(n_202), .B1(n_433), .B2(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g628 ( .A(n_63), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_64), .A2(n_181), .B1(n_427), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_65), .A2(n_116), .B1(n_463), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_66), .A2(n_173), .B1(n_445), .B2(n_568), .Y(n_1040) );
INVx2_ASAP7_75t_L g287 ( .A(n_67), .Y(n_287) );
AOI21xp33_ASAP7_75t_L g532 ( .A1(n_68), .A2(n_402), .B(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_70), .A2(n_195), .B1(n_564), .B2(n_566), .Y(n_563) );
INVx1_ASAP7_75t_SL g791 ( .A(n_71), .Y(n_791) );
AND2x4_ASAP7_75t_L g793 ( .A(n_71), .B(n_287), .Y(n_793) );
INVx1_ASAP7_75t_L g797 ( .A(n_71), .Y(n_797) );
XOR2x2_ASAP7_75t_L g700 ( .A(n_73), .B(n_701), .Y(n_700) );
XOR2x2_ASAP7_75t_L g747 ( .A(n_73), .B(n_701), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_74), .A2(n_226), .B1(n_366), .B2(n_369), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_76), .A2(n_483), .B(n_486), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_77), .A2(n_166), .B1(n_494), .B2(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_78), .A2(n_212), .B1(n_788), .B2(n_792), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_79), .A2(n_148), .B1(n_431), .B2(n_433), .Y(n_430) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_80), .Y(n_309) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_81), .B(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_82), .A2(n_163), .B1(n_328), .B2(n_344), .Y(n_737) );
INVx1_ASAP7_75t_L g377 ( .A(n_83), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_85), .A2(n_213), .B1(n_328), .B2(n_330), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_86), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g409 ( .A(n_87), .Y(n_409) );
INVx1_ASAP7_75t_L g623 ( .A(n_89), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_90), .A2(n_241), .B1(n_445), .B2(n_561), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_93), .A2(n_146), .B1(n_425), .B2(n_427), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_96), .A2(n_105), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_97), .A2(n_1030), .B(n_1031), .Y(n_1029) );
CKINVDCx16_ASAP7_75t_R g823 ( .A(n_98), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_99), .A2(n_194), .B1(n_551), .B2(n_774), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_100), .A2(n_183), .B1(n_821), .B2(n_881), .Y(n_880) );
XNOR2x1_ASAP7_75t_L g384 ( .A(n_101), .B(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_103), .A2(n_234), .B1(n_561), .B2(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g310 ( .A(n_104), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_104), .B(n_220), .Y(n_348) );
INVx1_ASAP7_75t_L g534 ( .A(n_106), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_108), .A2(n_130), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_109), .A2(n_174), .B1(n_431), .B2(n_568), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_110), .A2(n_172), .B1(n_506), .B2(n_1035), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_112), .A2(n_211), .B1(n_420), .B2(n_422), .Y(n_448) );
INVx1_ASAP7_75t_L g809 ( .A(n_113), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_115), .A2(n_185), .B1(n_833), .B2(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_117), .B(n_396), .Y(n_1062) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_118), .A2(n_199), .B1(n_420), .B2(n_422), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_119), .A2(n_273), .B1(n_354), .B2(n_360), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_122), .A2(n_238), .B1(n_561), .B2(n_1039), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_123), .A2(n_154), .B1(n_633), .B2(n_672), .C(n_673), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_123), .A2(n_154), .B1(n_633), .B2(n_672), .C(n_673), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_124), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_125), .A2(n_214), .B1(n_436), .B2(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_126), .A2(n_229), .B1(n_406), .B2(n_411), .Y(n_530) );
INVx1_ASAP7_75t_L g553 ( .A(n_127), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_128), .A2(n_224), .B1(n_420), .B2(n_422), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_129), .A2(n_264), .B1(n_433), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_132), .A2(n_137), .B1(n_600), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_133), .A2(n_200), .B1(n_420), .B2(n_526), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_134), .A2(n_180), .B1(n_445), .B2(n_561), .Y(n_655) );
INVx1_ASAP7_75t_L g1032 ( .A(n_135), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_136), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_136), .A2(n_190), .B1(n_827), .B2(n_830), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_138), .A2(n_203), .B1(n_422), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g464 ( .A(n_140), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_141), .A2(n_228), .B1(n_358), .B2(n_372), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_142), .A2(n_219), .B1(n_360), .B2(n_363), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_143), .A2(n_249), .B1(n_363), .B2(n_371), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_144), .A2(n_162), .B1(n_687), .B2(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g605 ( .A(n_145), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_147), .A2(n_150), .B1(n_360), .B2(n_363), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_149), .A2(n_250), .B1(n_436), .B2(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g1066 ( .A(n_151), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_152), .A2(n_231), .B1(n_436), .B2(n_438), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_153), .A2(n_272), .B1(n_568), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_155), .A2(n_204), .B1(n_691), .B2(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g601 ( .A(n_156), .Y(n_601) );
INVx1_ASAP7_75t_L g593 ( .A(n_157), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_158), .A2(n_233), .B1(n_360), .B2(n_363), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_159), .A2(n_276), .B1(n_664), .B2(n_666), .Y(n_771) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_160), .A2(n_455), .B(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_161), .A2(n_179), .B1(n_562), .B2(n_566), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_164), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_165), .A2(n_225), .B1(n_722), .B2(n_723), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_167), .A2(n_188), .B1(n_354), .B2(n_358), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_168), .A2(n_254), .B1(n_427), .B2(n_566), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_169), .A2(n_256), .B1(n_795), .B2(n_799), .Y(n_794) );
INVx1_ASAP7_75t_L g813 ( .A(n_170), .Y(n_813) );
INVx1_ASAP7_75t_L g811 ( .A(n_171), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_175), .A2(n_189), .B1(n_502), .B2(n_611), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_176), .A2(n_245), .B1(n_420), .B2(n_422), .Y(n_1042) );
CKINVDCx14_ASAP7_75t_R g731 ( .A(n_177), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_184), .A2(n_1053), .B1(n_1054), .B2(n_1068), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1053 ( .A(n_184), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_186), .B(n_676), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_187), .B(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_191), .A2(n_389), .B(n_391), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_193), .A2(n_251), .B1(n_415), .B2(n_471), .Y(n_470) );
OA22x2_ASAP7_75t_L g314 ( .A1(n_196), .A2(n_221), .B1(n_309), .B2(n_313), .Y(n_314) );
INVx1_ASAP7_75t_L g337 ( .A(n_196), .Y(n_337) );
INVx1_ASAP7_75t_L g461 ( .A(n_197), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_201), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_205), .A2(n_270), .B1(n_455), .B2(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g614 ( .A(n_206), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_207), .A2(n_259), .B1(n_450), .B2(n_611), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_208), .A2(n_223), .B1(n_489), .B2(n_506), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_209), .A2(n_258), .B1(n_687), .B2(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g404 ( .A(n_210), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_215), .B(n_396), .Y(n_395) );
CKINVDCx6p67_ASAP7_75t_R g822 ( .A(n_216), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_218), .A2(n_237), .B1(n_366), .B2(n_369), .Y(n_365) );
INVx1_ASAP7_75t_L g326 ( .A(n_220), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_220), .B(n_335), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g338 ( .A1(n_221), .A2(n_242), .B(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_227), .A2(n_246), .B1(n_821), .B2(n_835), .Y(n_834) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_230), .A2(n_551), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g630 ( .A(n_235), .Y(n_630) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_236), .Y(n_677) );
INVx1_ASAP7_75t_L g400 ( .A(n_239), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_240), .A2(n_277), .B1(n_371), .B2(n_372), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_242), .B(n_268), .Y(n_291) );
INVx1_ASAP7_75t_L g312 ( .A(n_242), .Y(n_312) );
INVx1_ASAP7_75t_L g1025 ( .A(n_246), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_246), .B(n_1041), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_246), .A2(n_1052), .B1(n_1069), .B2(n_1071), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_247), .A2(n_279), .B1(n_427), .B2(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g896 ( .A(n_248), .Y(n_896) );
INVx1_ASAP7_75t_L g647 ( .A(n_252), .Y(n_647) );
INVx1_ASAP7_75t_SL g613 ( .A(n_253), .Y(n_613) );
INVx1_ASAP7_75t_L g514 ( .A(n_256), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_257), .A2(n_715), .B(n_716), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_260), .A2(n_269), .B1(n_436), .B2(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g718 ( .A(n_261), .Y(n_718) );
AOI21xp33_ASAP7_75t_SL g374 ( .A1(n_262), .A2(n_375), .B(n_376), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_263), .B(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_265), .Y(n_775) );
AOI22xp5_ASAP7_75t_SL g1063 ( .A1(n_266), .A2(n_275), .B1(n_332), .B2(n_341), .Y(n_1063) );
INVx1_ASAP7_75t_L g674 ( .A(n_267), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_268), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_271), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g790 ( .A(n_274), .Y(n_790) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_274), .Y(n_1073) );
INVx1_ASAP7_75t_L g457 ( .A(n_278), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_293), .B(n_780), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
BUFx4_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NAND3xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .C(n_292), .Y(n_284) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_285), .B(n_1049), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_285), .B(n_1050), .Y(n_1070) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_285), .A2(n_292), .B(n_791), .Y(n_1074) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AO21x1_ASAP7_75t_L g1072 ( .A1(n_286), .A2(n_1073), .B(n_1074), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND3x4_ASAP7_75t_L g788 ( .A(n_287), .B(n_789), .C(n_791), .Y(n_788) );
AND2x2_ASAP7_75t_L g796 ( .A(n_287), .B(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_288), .B(n_1050), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_289), .A2(n_381), .B(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g1050 ( .A(n_292), .Y(n_1050) );
XNOR2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_636), .Y(n_293) );
XOR2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_476), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_441), .B1(n_474), .B2(n_475), .Y(n_297) );
INVx1_ASAP7_75t_L g475 ( .A(n_298), .Y(n_475) );
XNOR2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_384), .Y(n_298) );
XNOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_302), .B(n_352), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_327), .C(n_340), .Y(n_302) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_315), .Y(n_305) );
AND2x4_ASAP7_75t_L g328 ( .A(n_306), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g354 ( .A(n_306), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g360 ( .A(n_306), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g398 ( .A(n_306), .B(n_315), .Y(n_398) );
AND2x2_ASAP7_75t_L g413 ( .A(n_306), .B(n_329), .Y(n_413) );
AND2x4_ASAP7_75t_L g426 ( .A(n_306), .B(n_373), .Y(n_426) );
AND2x2_ASAP7_75t_L g437 ( .A(n_306), .B(n_361), .Y(n_437) );
AND2x2_ASAP7_75t_L g565 ( .A(n_306), .B(n_361), .Y(n_565) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_314), .Y(n_306) );
INVx1_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
NAND2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g313 ( .A(n_309), .Y(n_313) );
INVx3_ASAP7_75t_L g319 ( .A(n_309), .Y(n_319) );
NAND2xp33_ASAP7_75t_L g325 ( .A(n_309), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_310), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_312), .A2(n_339), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g349 ( .A(n_314), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
AND2x4_ASAP7_75t_L g332 ( .A(n_315), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g369 ( .A(n_315), .B(n_367), .Y(n_369) );
AND2x2_ASAP7_75t_L g375 ( .A(n_315), .B(n_342), .Y(n_375) );
AND2x4_ASAP7_75t_L g403 ( .A(n_315), .B(n_342), .Y(n_403) );
AND2x4_ASAP7_75t_L g407 ( .A(n_315), .B(n_333), .Y(n_407) );
AND2x2_ASAP7_75t_L g423 ( .A(n_315), .B(n_367), .Y(n_423) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g329 ( .A(n_317), .B(n_321), .Y(n_329) );
AND2x2_ASAP7_75t_L g345 ( .A(n_317), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g356 ( .A(n_317), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g361 ( .A(n_317), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_319), .B(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g335 ( .A(n_319), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_320), .B(n_334), .C(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
AND2x4_ASAP7_75t_L g341 ( .A(n_329), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g366 ( .A(n_329), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g390 ( .A(n_329), .B(n_342), .Y(n_390) );
AND2x4_ASAP7_75t_L g421 ( .A(n_329), .B(n_367), .Y(n_421) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g358 ( .A(n_333), .B(n_355), .Y(n_358) );
AND2x4_ASAP7_75t_L g363 ( .A(n_333), .B(n_361), .Y(n_363) );
AND2x4_ASAP7_75t_L g428 ( .A(n_333), .B(n_355), .Y(n_428) );
AND2x4_ASAP7_75t_L g440 ( .A(n_333), .B(n_361), .Y(n_440) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_338), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x4_ASAP7_75t_L g367 ( .A(n_343), .B(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g717 ( .A(n_344), .Y(n_717) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
AND2x4_ASAP7_75t_L g416 ( .A(n_345), .B(n_349), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
NAND4xp25_ASAP7_75t_SL g352 ( .A(n_353), .B(n_359), .C(n_364), .D(n_374), .Y(n_352) );
AND2x4_ASAP7_75t_L g434 ( .A(n_355), .B(n_367), .Y(n_434) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g373 ( .A(n_356), .Y(n_373) );
INVx1_ASAP7_75t_L g362 ( .A(n_357), .Y(n_362) );
AND2x4_ASAP7_75t_L g371 ( .A(n_361), .B(n_367), .Y(n_371) );
AND2x4_ASAP7_75t_L g432 ( .A(n_361), .B(n_367), .Y(n_432) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_370), .Y(n_364) );
AND2x4_ASAP7_75t_L g372 ( .A(n_367), .B(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_378), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g720 ( .A(n_378), .Y(n_720) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g394 ( .A(n_379), .Y(n_394) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_379), .Y(n_648) );
INVx2_ASAP7_75t_SL g676 ( .A(n_379), .Y(n_676) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g473 ( .A(n_380), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_417), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_399), .C(n_408), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_395), .Y(n_387) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g456 ( .A(n_390), .Y(n_456) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_390), .Y(n_505) );
BUFx3_ASAP7_75t_L g529 ( .A(n_390), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g469 ( .A(n_397), .Y(n_469) );
INVx2_ASAP7_75t_L g485 ( .A(n_397), .Y(n_485) );
INVx2_ASAP7_75t_L g644 ( .A(n_397), .Y(n_644) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g557 ( .A(n_398), .Y(n_557) );
BUFx3_ASAP7_75t_L g592 ( .A(n_398), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_404), .B2(n_405), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx3_ASAP7_75t_L g463 ( .A(n_403), .Y(n_463) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_403), .Y(n_551) );
INVx2_ASAP7_75t_L g590 ( .A(n_403), .Y(n_590) );
BUFx8_ASAP7_75t_SL g722 ( .A(n_403), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_405), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g669 ( .A(n_406), .Y(n_669) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx3_ASAP7_75t_L g465 ( .A(n_407), .Y(n_465) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_407), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_414), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_412), .Y(n_727) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
BUFx4f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx5_ASAP7_75t_L g490 ( .A(n_416), .Y(n_490) );
BUFx2_ASAP7_75t_L g549 ( .A(n_416), .Y(n_549) );
BUFx2_ASAP7_75t_L g650 ( .A(n_416), .Y(n_650) );
NOR2xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_429), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_424), .Y(n_418) );
BUFx12f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_421), .Y(n_494) );
INVx3_ASAP7_75t_L g525 ( .A(n_421), .Y(n_525) );
INVx1_ASAP7_75t_L g615 ( .A(n_422), .Y(n_615) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g526 ( .A(n_423), .Y(n_526) );
BUFx5_ASAP7_75t_L g689 ( .A(n_423), .Y(n_689) );
INVx1_ASAP7_75t_L g707 ( .A(n_423), .Y(n_707) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_426), .Y(n_447) );
BUFx3_ASAP7_75t_L g502 ( .A(n_426), .Y(n_502) );
BUFx12f_ASAP7_75t_L g566 ( .A(n_426), .Y(n_566) );
BUFx3_ASAP7_75t_L g682 ( .A(n_427), .Y(n_682) );
BUFx12f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx6_ASAP7_75t_L g519 ( .A(n_428), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_435), .Y(n_429) );
BUFx12f_ASAP7_75t_L g608 ( .A(n_431), .Y(n_608) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_431), .Y(n_691) );
BUFx12f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_432), .Y(n_445) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_432), .Y(n_499) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_433), .Y(n_757) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_434), .Y(n_500) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_434), .Y(n_521) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_434), .Y(n_561) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx8_ASAP7_75t_L g611 ( .A(n_437), .Y(n_611) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx4_ASAP7_75t_L g450 ( .A(n_439), .Y(n_450) );
INVx4_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
INVx1_ASAP7_75t_L g568 ( .A(n_439), .Y(n_568) );
INVx4_ASAP7_75t_L g584 ( .A(n_439), .Y(n_584) );
INVx1_ASAP7_75t_L g712 ( .A(n_439), .Y(n_712) );
INVx8_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_451), .Y(n_442) );
AND4x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .C(n_448), .D(n_449), .Y(n_443) );
BUFx3_ASAP7_75t_L g600 ( .A(n_447), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_460), .C(n_466), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_457), .B2(n_458), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g1030 ( .A(n_456), .Y(n_1030) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_464), .B2(n_465), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g508 ( .A(n_465), .Y(n_508) );
INVx2_ASAP7_75t_L g774 ( .A(n_465), .Y(n_774) );
OAI21xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g624 ( .A(n_471), .Y(n_624) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g769 ( .A(n_472), .Y(n_769) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g535 ( .A(n_473), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_594), .B1(n_634), .B2(n_635), .Y(n_476) );
INVx1_ASAP7_75t_L g635 ( .A(n_477), .Y(n_635) );
XNOR2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_539), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_510), .B1(n_536), .B2(n_538), .Y(n_478) );
INVx1_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
XNOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_509), .Y(n_480) );
NAND4xp75_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .C(n_497), .D(n_503), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_491), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g633 ( .A(n_490), .Y(n_633) );
INVx2_ASAP7_75t_L g1035 ( .A(n_490), .Y(n_1035) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
BUFx3_ASAP7_75t_L g681 ( .A(n_500), .Y(n_681) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx3_ASAP7_75t_L g631 ( .A(n_506), .Y(n_631) );
BUFx3_ASAP7_75t_L g666 ( .A(n_506), .Y(n_666) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g537 ( .A(n_513), .Y(n_537) );
XNOR2x1_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_516), .B(n_527), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .C(n_522), .D(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g604 ( .A(n_518), .Y(n_604) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_518), .Y(n_763) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g562 ( .A(n_519), .Y(n_562) );
INVx1_ASAP7_75t_L g710 ( .A(n_519), .Y(n_710) );
INVx2_ASAP7_75t_L g1039 ( .A(n_519), .Y(n_1039) );
BUFx3_ASAP7_75t_L g609 ( .A(n_521), .Y(n_609) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_525), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g687 ( .A(n_525), .Y(n_687) );
BUFx2_ASAP7_75t_L g752 ( .A(n_526), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .C(n_531), .D(n_532), .Y(n_527) );
INVx2_ASAP7_75t_L g665 ( .A(n_529), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_535), .B(n_1066), .Y(n_1065) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
XNOR2x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_576), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .B(n_570), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_543), .B(n_558), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_546), .B(n_559), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_554), .C(n_558), .Y(n_546) );
INVx1_ASAP7_75t_L g574 ( .A(n_547), .Y(n_574) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
BUFx3_ASAP7_75t_L g668 ( .A(n_551), .Y(n_668) );
INVxp67_ASAP7_75t_L g572 ( .A(n_554), .Y(n_572) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g715 ( .A(n_556), .Y(n_715) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g620 ( .A(n_557), .Y(n_620) );
INVx1_ASAP7_75t_L g575 ( .A(n_559), .Y(n_575) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .C(n_567), .D(n_569), .Y(n_559) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_565), .Y(n_654) );
BUFx3_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .C(n_574), .Y(n_571) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
XOR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_593), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_585), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .C(n_582), .D(n_583), .Y(n_579) );
BUFx2_ASAP7_75t_L g692 ( .A(n_584), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_588), .D(n_591), .Y(n_585) );
INVx2_ASAP7_75t_L g627 ( .A(n_589), .Y(n_627) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g773 ( .A(n_590), .Y(n_773) );
BUFx3_ASAP7_75t_L g767 ( .A(n_592), .Y(n_767) );
INVx2_ASAP7_75t_L g634 ( .A(n_594), .Y(n_634) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_616), .Y(n_596) );
NOR3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_606), .C(n_612), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B1(n_602), .B2(n_605), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_610), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_625), .C(n_629), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_618), .B(n_621), .Y(n_617) );
BUFx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_632), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_697), .B1(n_778), .B2(n_779), .Y(n_636) );
INVx1_ASAP7_75t_L g778 ( .A(n_637), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_659), .B1(n_695), .B2(n_696), .Y(n_637) );
INVx1_ASAP7_75t_L g695 ( .A(n_638), .Y(n_695) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g657 ( .A(n_640), .Y(n_657) );
NOR2xp67_ASAP7_75t_L g640 ( .A(n_641), .B(n_651), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .C(n_645), .D(n_649), .Y(n_641) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_644), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g1031 ( .A(n_648), .B(n_1032), .Y(n_1031) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .C(n_655), .D(n_656), .Y(n_651) );
INVx2_ASAP7_75t_SL g696 ( .A(n_659), .Y(n_696) );
AO22x2_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_677), .B1(n_678), .B2(n_693), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_670), .C(n_677), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND4xp75_ASAP7_75t_SL g693 ( .A(n_662), .B(n_679), .C(n_685), .D(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_R g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_685), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .Y(n_685) );
BUFx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g759 ( .A(n_691), .Y(n_759) );
INVx1_ASAP7_75t_L g779 ( .A(n_697), .Y(n_779) );
XOR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_748), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_728), .B1(n_729), .B2(n_747), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_713), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_708), .C(n_709), .D(n_711), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_721), .C(n_725), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_719), .Y(n_716) );
BUFx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B(n_744), .Y(n_730) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_731), .B(n_745), .C(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_739), .Y(n_733) );
INVx1_ASAP7_75t_L g746 ( .A(n_734), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .C(n_737), .D(n_738), .Y(n_734) );
INVxp67_ASAP7_75t_L g745 ( .A(n_739), .Y(n_745) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .C(n_742), .D(n_743), .Y(n_739) );
AO211x2_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_760), .B(n_776), .C(n_777), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_754), .Y(n_749) );
AO22x2_ASAP7_75t_L g777 ( .A1(n_750), .A2(n_761), .B1(n_775), .B2(n_1077), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_753), .Y(n_750) );
AO22x1_ASAP7_75t_L g776 ( .A1(n_754), .A2(n_770), .B1(n_775), .B2(n_1076), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_770), .C(n_775), .Y(n_760) );
NAND2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_768), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_1020), .B1(n_1023), .B2(n_1047), .C(n_1051), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_943), .C(n_986), .Y(n_781) );
NAND5xp2_ASAP7_75t_L g782 ( .A(n_783), .B(n_883), .C(n_913), .D(n_922), .E(n_938), .Y(n_782) );
OAI31xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_836), .A3(n_857), .B(n_873), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_803), .Y(n_784) );
INVx1_ASAP7_75t_L g961 ( .A(n_785), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_800), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_786), .Y(n_844) );
AND2x2_ASAP7_75t_L g868 ( .A(n_786), .B(n_840), .Y(n_868) );
AND2x2_ASAP7_75t_L g888 ( .A(n_786), .B(n_847), .Y(n_888) );
OR2x2_ASAP7_75t_L g985 ( .A(n_786), .B(n_800), .Y(n_985) );
AND2x4_ASAP7_75t_SL g786 ( .A(n_787), .B(n_794), .Y(n_786) );
INVx1_ASAP7_75t_L g808 ( .A(n_788), .Y(n_808) );
AND2x4_ASAP7_75t_L g792 ( .A(n_789), .B(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_789), .B(n_793), .Y(n_810) );
AND2x4_ASAP7_75t_L g821 ( .A(n_789), .B(n_796), .Y(n_821) );
AND2x4_ASAP7_75t_L g835 ( .A(n_789), .B(n_793), .Y(n_835) );
INVx2_ASAP7_75t_SL g882 ( .A(n_792), .Y(n_882) );
AND2x2_ASAP7_75t_L g799 ( .A(n_793), .B(n_798), .Y(n_799) );
AND2x4_ASAP7_75t_L g830 ( .A(n_793), .B(n_798), .Y(n_830) );
AND2x2_ASAP7_75t_L g833 ( .A(n_793), .B(n_798), .Y(n_833) );
INVx1_ASAP7_75t_L g816 ( .A(n_795), .Y(n_816) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .Y(n_795) );
AND2x4_ASAP7_75t_L g827 ( .A(n_796), .B(n_798), .Y(n_827) );
AND2x2_ASAP7_75t_L g842 ( .A(n_796), .B(n_798), .Y(n_842) );
INVx1_ASAP7_75t_L g814 ( .A(n_799), .Y(n_814) );
AND2x2_ASAP7_75t_L g838 ( .A(n_800), .B(n_839), .Y(n_838) );
CKINVDCx6p67_ASAP7_75t_R g849 ( .A(n_800), .Y(n_849) );
INVx1_ASAP7_75t_L g863 ( .A(n_800), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_800), .B(n_844), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_800), .B(n_846), .Y(n_951) );
AND2x2_ASAP7_75t_L g962 ( .A(n_800), .B(n_953), .Y(n_962) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_817), .Y(n_804) );
AND2x2_ASAP7_75t_L g848 ( .A(n_805), .B(n_849), .Y(n_848) );
AND2x2_ASAP7_75t_L g861 ( .A(n_805), .B(n_862), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_805), .B(n_887), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g903 ( .A(n_805), .B(n_904), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_805), .B(n_909), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_805), .B(n_868), .Y(n_976) );
NOR2x1p5_ASAP7_75t_L g984 ( .A(n_805), .B(n_985), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_805), .B(n_855), .Y(n_995) );
INVx1_ASAP7_75t_L g1004 ( .A(n_805), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_805), .B(n_858), .Y(n_1012) );
CKINVDCx6p67_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g854 ( .A(n_806), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g871 ( .A(n_806), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_806), .B(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g928 ( .A(n_806), .B(n_846), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_806), .B(n_818), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_806), .B(n_933), .Y(n_932) );
AND2x2_ASAP7_75t_L g953 ( .A(n_806), .B(n_868), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_806), .B(n_849), .Y(n_1019) );
OR2x6_ASAP7_75t_SL g806 ( .A(n_807), .B(n_812), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_810), .A2(n_820), .B1(n_822), .B2(n_823), .Y(n_819) );
OAI221xp5_ASAP7_75t_L g894 ( .A1(n_810), .A2(n_820), .B1(n_895), .B2(n_896), .C(n_897), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .B1(n_815), .B2(n_816), .Y(n_812) );
OAI221xp5_ASAP7_75t_L g901 ( .A1(n_817), .A2(n_902), .B1(n_908), .B2(n_910), .C(n_911), .Y(n_901) );
INVx1_ASAP7_75t_L g921 ( .A(n_817), .Y(n_921) );
OR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_831), .Y(n_817) );
AND2x2_ASAP7_75t_L g851 ( .A(n_818), .B(n_852), .Y(n_851) );
INVx3_ASAP7_75t_L g855 ( .A(n_818), .Y(n_855) );
INVx2_ASAP7_75t_L g866 ( .A(n_818), .Y(n_866) );
AND2x2_ASAP7_75t_L g909 ( .A(n_818), .B(n_831), .Y(n_909) );
OR2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .Y(n_818) );
INVx1_ASAP7_75t_L g1022 ( .A(n_820), .Y(n_1022) );
INVx3_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_826), .B1(n_828), .B2(n_829), .Y(n_824) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g852 ( .A(n_831), .Y(n_852) );
AND2x2_ASAP7_75t_L g937 ( .A(n_831), .B(n_855), .Y(n_937) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_831), .B(n_878), .Y(n_1001) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_834), .Y(n_831) );
A2O1A1Ixp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_845), .B(n_850), .C(n_853), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_SL g856 ( .A(n_839), .B(n_849), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_839), .B(n_870), .Y(n_910) );
AND2x2_ASAP7_75t_L g954 ( .A(n_839), .B(n_861), .Y(n_954) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
INVx1_ASAP7_75t_L g847 ( .A(n_840), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
AND2x2_ASAP7_75t_L g846 ( .A(n_844), .B(n_847), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_844), .B(n_862), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_844), .B(n_861), .Y(n_998) );
INVx1_ASAP7_75t_L g919 ( .A(n_845), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .Y(n_845) );
AND2x2_ASAP7_75t_L g860 ( .A(n_846), .B(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g917 ( .A(n_846), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_L g947 ( .A1(n_846), .A2(n_948), .B(n_949), .C(n_950), .Y(n_947) );
OAI211xp5_ASAP7_75t_L g973 ( .A1(n_846), .A2(n_974), .B(n_975), .C(n_976), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_847), .B(n_862), .Y(n_892) );
AND2x2_ASAP7_75t_L g907 ( .A(n_847), .B(n_862), .Y(n_907) );
AND2x2_ASAP7_75t_L g933 ( .A(n_847), .B(n_849), .Y(n_933) );
INVx1_ASAP7_75t_L g972 ( .A(n_847), .Y(n_972) );
AND2x2_ASAP7_75t_L g887 ( .A(n_849), .B(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_849), .B(n_868), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_849), .B(n_899), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_849), .B(n_928), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_850), .B(n_874), .Y(n_958) );
AOI21xp33_ASAP7_75t_L g997 ( .A1(n_850), .A2(n_869), .B(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_851), .B(n_870), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_851), .B(n_887), .Y(n_1015) );
INVx3_ASAP7_75t_L g858 ( .A(n_852), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_852), .B(n_878), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_852), .B(n_877), .Y(n_978) );
OR2x2_ASAP7_75t_L g982 ( .A(n_852), .B(n_878), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_854), .B(n_888), .Y(n_975) );
INVx1_ASAP7_75t_L g890 ( .A(n_855), .Y(n_890) );
AOI21xp33_ASAP7_75t_L g950 ( .A1(n_855), .A2(n_906), .B(n_951), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_855), .B(n_876), .Y(n_965) );
AND2x2_ASAP7_75t_L g983 ( .A(n_855), .B(n_877), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_856), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g1010 ( .A(n_856), .Y(n_1010) );
AOI32xp33_ASAP7_75t_SL g857 ( .A1(n_858), .A2(n_859), .A3(n_864), .B1(n_869), .B2(n_872), .Y(n_857) );
INVx3_ASAP7_75t_L g872 ( .A(n_858), .Y(n_872) );
AOI31xp33_ASAP7_75t_L g943 ( .A1(n_858), .A2(n_944), .A3(n_955), .B(n_956), .Y(n_943) );
INVx1_ASAP7_75t_L g1013 ( .A(n_858), .Y(n_1013) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_859), .A2(n_925), .B(n_1015), .C(n_1016), .Y(n_1014) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AND2x2_ASAP7_75t_L g867 ( .A(n_861), .B(n_868), .Y(n_867) );
INVxp67_ASAP7_75t_SL g974 ( .A(n_861), .Y(n_974) );
AND2x2_ASAP7_75t_L g927 ( .A(n_862), .B(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g884 ( .A(n_864), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_865), .B(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
BUFx2_ASAP7_75t_L g926 ( .A(n_866), .Y(n_926) );
INVx1_ASAP7_75t_L g899 ( .A(n_868), .Y(n_899) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_868), .B(n_1018), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_870), .B(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_870), .B(n_937), .Y(n_969) );
INVx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_872), .B(n_893), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_872), .A2(n_920), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI32xp33_ASAP7_75t_L g967 ( .A1(n_873), .A2(n_968), .A3(n_970), .B1(n_973), .B2(n_977), .Y(n_967) );
INVx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_874), .A2(n_945), .B1(n_957), .B2(n_966), .Y(n_956) );
INVx3_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_877), .B(n_914), .Y(n_955) );
NOR3xp33_ASAP7_75t_L g993 ( .A(n_877), .B(n_994), .C(n_996), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_877), .B(n_914), .Y(n_1006) );
INVx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AND2x2_ASAP7_75t_L g920 ( .A(n_878), .B(n_921), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_878), .B(n_909), .Y(n_991) );
AND2x4_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
OAI321xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .A3(n_889), .B1(n_898), .B2(n_901), .C(n_912), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_885), .A2(n_1008), .B1(n_1011), .B2(n_1013), .C(n_1014), .Y(n_1007) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_888), .B(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g996 ( .A(n_888), .Y(n_996) );
OAI21xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_891), .B(n_893), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_892), .B(n_931), .Y(n_930) );
CKINVDCx16_ASAP7_75t_R g911 ( .A(n_893), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_893), .B(n_936), .Y(n_935) );
AOI221xp5_ASAP7_75t_SL g963 ( .A1(n_893), .A2(n_923), .B1(n_941), .B2(n_954), .C(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
BUFx3_ASAP7_75t_L g914 ( .A(n_894), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g946 ( .A(n_903), .Y(n_946) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
OAI21xp33_ASAP7_75t_L g999 ( .A1(n_906), .A2(n_1000), .B(n_1002), .Y(n_999) );
INVx1_ASAP7_75t_L g1009 ( .A(n_907), .Y(n_1009) );
OAI211xp5_ASAP7_75t_L g945 ( .A1(n_908), .A2(n_946), .B(n_947), .C(n_952), .Y(n_945) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
O2A1O1Ixp33_ASAP7_75t_L g980 ( .A1(n_911), .A2(n_981), .B(n_983), .C(n_984), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_912), .A2(n_930), .B1(n_932), .B2(n_934), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_919), .B2(n_920), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_914), .A2(n_987), .B1(n_1006), .B2(n_1007), .Y(n_986) );
AOI21xp33_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_917), .B(n_918), .Y(n_915) );
INVx1_ASAP7_75t_L g1005 ( .A(n_916), .Y(n_1005) );
INVx1_ASAP7_75t_L g949 ( .A(n_918), .Y(n_949) );
INVx1_ASAP7_75t_L g942 ( .A(n_920), .Y(n_942) );
O2A1O1Ixp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_925), .B(n_927), .C(n_929), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
OAI211xp5_ASAP7_75t_L g988 ( .A1(n_924), .A2(n_951), .B(n_989), .C(n_992), .Y(n_988) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVxp67_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g952 ( .A1(n_937), .A2(n_953), .B(n_954), .Y(n_952) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVxp67_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g1002 ( .A1(n_948), .A2(n_964), .B(n_1003), .C(n_1005), .Y(n_1002) );
OAI211xp5_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_959), .B(n_960), .C(n_963), .Y(n_957) );
INVx1_ASAP7_75t_L g979 ( .A(n_962), .Y(n_979) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_979), .C(n_980), .Y(n_966) );
INVxp67_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
NOR3xp33_ASAP7_75t_L g987 ( .A(n_988), .B(n_997), .C(n_999), .Y(n_987) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
CKINVDCx14_ASAP7_75t_R g1003 ( .A(n_1004), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_1021), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
OAI21x1_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1026), .B(n_1044), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1036), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_1027), .B(n_1045), .C(n_1046), .Y(n_1044) );
AND4x1_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .C(n_1033), .D(n_1034), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1041), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_1037), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1040), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
CKINVDCx16_ASAP7_75t_R g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1054), .Y(n_1068) );
INVxp33_ASAP7_75t_SL g1054 ( .A(n_1055), .Y(n_1054) );
NOR2x1_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1061), .Y(n_1055) );
NAND4xp25_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .C(n_1059), .D(n_1060), .Y(n_1056) );
NAND4xp25_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .C(n_1064), .D(n_1067), .Y(n_1061) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
endmodule