module real_aes_258_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_832, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_833, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_832;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_833;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g233 ( .A(n_0), .B(n_155), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_1), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g148 ( .A(n_2), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_3), .B(n_161), .Y(n_174) );
NAND2xp33_ASAP7_75t_SL g225 ( .A(n_4), .B(n_159), .Y(n_225) );
INVx1_ASAP7_75t_L g206 ( .A(n_5), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_6), .B(n_179), .Y(n_552) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_7), .A2(n_122), .B1(n_123), .B2(n_125), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g532 ( .A(n_8), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_9), .Y(n_112) );
AND2x2_ASAP7_75t_L g172 ( .A(n_10), .B(n_165), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_11), .Y(n_499) );
INVxp33_ASAP7_75t_L g830 ( .A(n_12), .Y(n_830) );
INVx2_ASAP7_75t_L g166 ( .A(n_13), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_14), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_15), .B(n_111), .C(n_113), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_15), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_15), .B(n_28), .Y(n_728) );
INVx1_ASAP7_75t_L g560 ( .A(n_16), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g817 ( .A1(n_17), .A2(n_28), .B1(n_782), .B2(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_17), .Y(n_818) );
AOI221x1_ASAP7_75t_L g219 ( .A1(n_18), .A2(n_143), .B1(n_220), .B2(n_222), .C(n_224), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_19), .B(n_161), .Y(n_194) );
INVx1_ASAP7_75t_L g116 ( .A(n_20), .Y(n_116) );
INVx1_ASAP7_75t_L g558 ( .A(n_21), .Y(n_558) );
INVx1_ASAP7_75t_SL g481 ( .A(n_22), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_23), .B(n_162), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_24), .A2(n_143), .B(n_176), .Y(n_175) );
AOI221xp5_ASAP7_75t_SL g186 ( .A1(n_25), .A2(n_41), .B1(n_143), .B2(n_161), .C(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_26), .B(n_155), .Y(n_177) );
AOI33xp33_ASAP7_75t_L g518 ( .A1(n_27), .A2(n_54), .A3(n_209), .B1(n_215), .B2(n_519), .B3(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g782 ( .A(n_28), .Y(n_782) );
INVx1_ASAP7_75t_L g492 ( .A(n_29), .Y(n_492) );
OR2x2_ASAP7_75t_L g167 ( .A(n_30), .B(n_94), .Y(n_167) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_30), .A2(n_94), .B(n_166), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_31), .B(n_151), .Y(n_198) );
INVxp67_ASAP7_75t_L g218 ( .A(n_32), .Y(n_218) );
AND2x2_ASAP7_75t_L g249 ( .A(n_33), .B(n_164), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_34), .B(n_207), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_35), .A2(n_143), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_36), .B(n_151), .Y(n_188) );
AND2x2_ASAP7_75t_L g144 ( .A(n_37), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g159 ( .A(n_37), .B(n_148), .Y(n_159) );
INVx1_ASAP7_75t_L g214 ( .A(n_37), .Y(n_214) );
INVxp67_ASAP7_75t_L g113 ( .A(n_38), .Y(n_113) );
OR2x6_ASAP7_75t_L g792 ( .A(n_38), .B(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_39), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_40), .B(n_207), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_42), .A2(n_179), .B1(n_223), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_43), .B(n_550), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_44), .A2(n_84), .B1(n_143), .B2(n_212), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_45), .B(n_162), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_46), .B(n_155), .Y(n_247) );
INVx1_ASAP7_75t_L g790 ( .A(n_47), .Y(n_790) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_48), .B(n_88), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_49), .B(n_199), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_50), .B(n_162), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_51), .Y(n_545) );
AND2x2_ASAP7_75t_L g236 ( .A(n_52), .B(n_164), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_53), .B(n_164), .Y(n_190) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_53), .B(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_55), .B(n_162), .Y(n_510) );
INVx1_ASAP7_75t_L g147 ( .A(n_56), .Y(n_147) );
INVx1_ASAP7_75t_L g157 ( .A(n_56), .Y(n_157) );
AND2x2_ASAP7_75t_L g511 ( .A(n_57), .B(n_164), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_58), .A2(n_77), .B1(n_207), .B2(n_212), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_59), .B(n_207), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_60), .B(n_161), .Y(n_248) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_61), .A2(n_121), .B1(n_126), .B2(n_127), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_61), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_62), .B(n_223), .Y(n_501) );
AOI21xp5_ASAP7_75t_SL g470 ( .A1(n_63), .A2(n_212), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g168 ( .A(n_64), .B(n_164), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_65), .B(n_151), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_66), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_67), .B(n_165), .Y(n_201) );
INVx1_ASAP7_75t_L g555 ( .A(n_68), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_69), .B(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_70), .A2(n_143), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g509 ( .A(n_71), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_72), .B(n_151), .Y(n_178) );
AND2x2_ASAP7_75t_SL g286 ( .A(n_73), .B(n_199), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_74), .A2(n_212), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g145 ( .A(n_75), .Y(n_145) );
INVx1_ASAP7_75t_L g153 ( .A(n_75), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_76), .B(n_207), .Y(n_521) );
AND2x2_ASAP7_75t_L g483 ( .A(n_78), .B(n_222), .Y(n_483) );
INVx1_ASAP7_75t_L g556 ( .A(n_79), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_80), .A2(n_212), .B(n_480), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_81), .A2(n_212), .B(n_282), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_82), .B(n_161), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_83), .A2(n_87), .B1(n_161), .B2(n_207), .Y(n_284) );
INVx1_ASAP7_75t_L g115 ( .A(n_85), .Y(n_115) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_86), .B(n_222), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_89), .A2(n_212), .B1(n_516), .B2(n_517), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_90), .B(n_155), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_91), .B(n_155), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_92), .B(n_795), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_93), .A2(n_143), .B(n_149), .Y(n_142) );
INVx1_ASAP7_75t_L g472 ( .A(n_95), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_96), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g522 ( .A(n_97), .B(n_222), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_98), .A2(n_490), .B(n_491), .C(n_493), .Y(n_489) );
INVxp67_ASAP7_75t_L g221 ( .A(n_99), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_100), .B(n_161), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_101), .B(n_151), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_102), .A2(n_143), .B(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_SL g788 ( .A(n_103), .Y(n_788) );
BUFx2_ASAP7_75t_L g804 ( .A(n_103), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_104), .B(n_162), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_117), .B(n_829), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_108), .B(n_830), .Y(n_829) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_114), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_115), .B(n_116), .Y(n_793) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_805), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_784), .B(n_799), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_128), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_120), .Y(n_828) );
INVxp33_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
INVx1_ASAP7_75t_L g125 ( .A(n_123), .Y(n_125) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_129), .Y(n_827) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_132), .B(n_458), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g783 ( .A(n_131), .Y(n_783) );
OR2x2_ASAP7_75t_L g791 ( .A(n_131), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_131), .B(n_798), .Y(n_797) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_397), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_290), .C(n_341), .Y(n_133) );
OAI211xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_180), .B(n_237), .C(n_268), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_169), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_139), .B(n_242), .Y(n_405) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g250 ( .A(n_140), .B(n_171), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_140), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g267 ( .A(n_140), .B(n_257), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_140), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g304 ( .A(n_140), .B(n_280), .Y(n_304) );
INVx2_ASAP7_75t_L g330 ( .A(n_140), .Y(n_330) );
AND2x4_ASAP7_75t_L g339 ( .A(n_140), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g444 ( .A(n_140), .B(n_311), .Y(n_444) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_163), .B(n_168), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_160), .Y(n_141) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
BUFx3_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
AND2x6_ASAP7_75t_L g155 ( .A(n_145), .B(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
AND2x4_ASAP7_75t_L g212 ( .A(n_146), .B(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g151 ( .A(n_147), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_154), .B(n_158), .Y(n_149) );
INVxp67_ASAP7_75t_L g561 ( .A(n_151), .Y(n_561) );
AND2x4_ASAP7_75t_L g162 ( .A(n_152), .B(n_156), .Y(n_162) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVxp67_ASAP7_75t_L g559 ( .A(n_155), .Y(n_559) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_158), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_158), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_158), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_158), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_158), .A2(n_246), .B(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_158), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_158), .A2(n_473), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_158), .A2(n_473), .B(n_509), .C(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g516 ( .A(n_158), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_158), .A2(n_473), .B(n_532), .C(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_158), .A2(n_548), .B(n_549), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_158), .B(n_179), .Y(n_562) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g161 ( .A(n_159), .B(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_159), .Y(n_493) );
INVx1_ASAP7_75t_L g226 ( .A(n_162), .Y(n_226) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_163), .A2(n_243), .B(n_249), .Y(n_242) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_163), .A2(n_243), .B(n_249), .Y(n_257) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_163), .A2(n_477), .B(n_483), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_164), .Y(n_163) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_164), .A2(n_186), .B(n_190), .Y(n_185) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AND2x4_ASAP7_75t_L g179 ( .A(n_166), .B(n_167), .Y(n_179) );
AND2x2_ASAP7_75t_L g328 ( .A(n_169), .B(n_329), .Y(n_328) );
OAI32xp33_ASAP7_75t_L g411 ( .A1(n_169), .A2(n_333), .A3(n_337), .B1(n_344), .B2(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_169), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g265 ( .A(n_170), .B(n_266), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_170), .B(n_260), .C(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g364 ( .A(n_170), .B(n_267), .Y(n_364) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_171), .Y(n_254) );
INVx5_ASAP7_75t_L g289 ( .A(n_171), .Y(n_289) );
AND2x4_ASAP7_75t_L g345 ( .A(n_171), .B(n_257), .Y(n_345) );
OR2x2_ASAP7_75t_L g360 ( .A(n_171), .B(n_280), .Y(n_360) );
OR2x2_ASAP7_75t_L g386 ( .A(n_171), .B(n_242), .Y(n_386) );
AND2x2_ASAP7_75t_L g394 ( .A(n_171), .B(n_340), .Y(n_394) );
AND2x4_ASAP7_75t_SL g419 ( .A(n_171), .B(n_339), .Y(n_419) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_179), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_179), .B(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_179), .B(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_179), .B(n_221), .Y(n_220) );
NOR3xp33_ASAP7_75t_L g224 ( .A(n_179), .B(n_225), .C(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_179), .A2(n_470), .B(n_475), .Y(n_469) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_181), .B(n_339), .Y(n_415) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_182), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x6_ASAP7_75t_SL g239 ( .A(n_183), .B(n_240), .Y(n_239) );
INVxp67_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g264 ( .A(n_184), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_184), .B(n_299), .Y(n_317) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_184), .Y(n_455) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
AND2x2_ASAP7_75t_L g297 ( .A(n_185), .B(n_228), .Y(n_297) );
INVx2_ASAP7_75t_L g325 ( .A(n_185), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_185), .B(n_192), .Y(n_366) );
BUFx3_ASAP7_75t_L g390 ( .A(n_185), .Y(n_390) );
OR2x2_ASAP7_75t_L g402 ( .A(n_185), .B(n_192), .Y(n_402) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_185), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_191), .A2(n_433), .B1(n_436), .B2(n_437), .Y(n_432) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
INVx1_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
OR2x2_ASAP7_75t_L g271 ( .A(n_192), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g278 ( .A(n_192), .Y(n_278) );
AND2x4_ASAP7_75t_SL g295 ( .A(n_192), .B(n_203), .Y(n_295) );
AND2x4_ASAP7_75t_L g300 ( .A(n_192), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g309 ( .A(n_192), .Y(n_309) );
OR2x2_ASAP7_75t_L g315 ( .A(n_192), .B(n_203), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_192), .B(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_192), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_192), .B(n_297), .Y(n_431) );
OR2x2_ASAP7_75t_L g447 ( .A(n_192), .B(n_350), .Y(n_447) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_199), .Y(n_193) );
INVx2_ASAP7_75t_SL g282 ( .A(n_199), .Y(n_282) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_199), .A2(n_530), .B(n_534), .Y(n_529) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g223 ( .A(n_200), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_202), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_202), .B(n_264), .Y(n_380) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_227), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_203), .B(n_228), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_203), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_203), .B(n_272), .Y(n_276) );
INVx3_ASAP7_75t_L g301 ( .A(n_203), .Y(n_301) );
INVx1_ASAP7_75t_L g334 ( .A(n_203), .Y(n_334) );
AND2x2_ASAP7_75t_L g414 ( .A(n_203), .B(n_278), .Y(n_414) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_219), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B1(n_212), .B2(n_217), .Y(n_204) );
INVx1_ASAP7_75t_L g502 ( .A(n_207), .Y(n_502) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_211), .Y(n_207) );
INVx1_ASAP7_75t_L g543 ( .A(n_208), .Y(n_543) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
OR2x6_ASAP7_75t_L g473 ( .A(n_209), .B(n_216), .Y(n_473) );
INVxp33_ASAP7_75t_L g519 ( .A(n_209), .Y(n_519) );
INVx1_ASAP7_75t_L g544 ( .A(n_211), .Y(n_544) );
INVxp67_ASAP7_75t_L g500 ( .A(n_212), .Y(n_500) );
NOR2x1p5_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g520 ( .A(n_215), .Y(n_520) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_222), .A2(n_489), .B1(n_494), .B2(n_495), .Y(n_488) );
INVx3_ASAP7_75t_L g495 ( .A(n_222), .Y(n_495) );
INVx4_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_223), .A2(n_230), .B(n_236), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_223), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_226), .B(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_226), .A2(n_473), .B1(n_555), .B2(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_228), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g299 ( .A(n_228), .Y(n_299) );
AND2x2_ASAP7_75t_L g324 ( .A(n_228), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g350 ( .A(n_228), .B(n_272), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_228), .B(n_301), .Y(n_367) );
INVx1_ASAP7_75t_L g373 ( .A(n_228), .Y(n_373) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AOI222xp33_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_241), .B1(n_251), .B2(n_258), .C1(n_261), .C2(n_265), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_250), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_242), .B(n_311), .Y(n_362) );
AND2x4_ASAP7_75t_L g378 ( .A(n_242), .B(n_289), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g303 ( .A(n_254), .B(n_304), .Y(n_303) );
AOI222xp33_ASAP7_75t_L g268 ( .A1(n_255), .A2(n_269), .B1(n_274), .B2(n_279), .C1(n_287), .C2(n_832), .Y(n_268) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g407 ( .A(n_256), .B(n_311), .Y(n_407) );
OR2x2_ASAP7_75t_L g450 ( .A(n_256), .B(n_356), .Y(n_450) );
AND2x2_ASAP7_75t_L g279 ( .A(n_257), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_257), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_L g368 ( .A1(n_258), .A2(n_369), .B(n_374), .C(n_375), .Y(n_368) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g396 ( .A(n_260), .Y(n_396) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g326 ( .A(n_265), .Y(n_326) );
AND2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g319 ( .A(n_266), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI31xp33_ASAP7_75t_L g361 ( .A1(n_269), .A2(n_287), .A3(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_270), .A2(n_320), .B(n_364), .C(n_365), .Y(n_363) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
OR2x2_ASAP7_75t_L g352 ( .A(n_271), .B(n_301), .Y(n_352) );
INVx2_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
BUFx2_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
AND2x2_ASAP7_75t_L g329 ( .A(n_280), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
AOI21x1_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_286), .Y(n_281) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_282), .A2(n_514), .B(n_522), .Y(n_513) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_282), .A2(n_514), .B(n_522), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_289), .B(n_346), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_302), .B(n_305), .C(n_327), .Y(n_290) );
INVxp33_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_298), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g331 ( .A(n_295), .B(n_324), .Y(n_331) );
OR2x2_ASAP7_75t_L g307 ( .A(n_296), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g337 ( .A(n_296), .B(n_311), .Y(n_337) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g413 ( .A(n_297), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g436 ( .A(n_298), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_300), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_300), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g448 ( .A(n_300), .B(n_324), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_300), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g391 ( .A(n_301), .B(n_373), .Y(n_391) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AOI322xp5_ASAP7_75t_L g445 ( .A1(n_304), .A2(n_324), .A3(n_378), .B1(n_403), .B2(n_446), .C1(n_448), .C2(n_449), .Y(n_445) );
AOI211xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_310), .B(n_312), .C(n_321), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_308), .B(n_336), .Y(n_358) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g323 ( .A(n_309), .B(n_324), .Y(n_323) );
NOR2x1p5_ASAP7_75t_L g389 ( .A(n_309), .B(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_309), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_310), .A2(n_328), .B(n_331), .C(n_332), .Y(n_327) );
AND2x4_ASAP7_75t_L g346 ( .A(n_311), .B(n_330), .Y(n_346) );
INVx2_ASAP7_75t_L g356 ( .A(n_311), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_311), .B(n_345), .Y(n_376) );
AND2x2_ASAP7_75t_L g418 ( .A(n_311), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_311), .B(n_435), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_311), .B(n_339), .Y(n_457) );
AOI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B(n_318), .Y(n_312) );
AND2x2_ASAP7_75t_L g408 ( .A(n_314), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_329), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g423 ( .A(n_329), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_335), .B(n_337), .C(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_336), .Y(n_420) );
INVx3_ASAP7_75t_SL g435 ( .A(n_339), .Y(n_435) );
NAND5xp2_ASAP7_75t_L g341 ( .A(n_342), .B(n_361), .C(n_368), .D(n_381), .E(n_392), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_351), .B2(n_353), .C1(n_357), .C2(n_359), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_344), .A2(n_425), .B1(n_429), .B2(n_430), .Y(n_424) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g374 ( .A(n_345), .B(n_346), .Y(n_374) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_355), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_356), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g393 ( .A(n_356), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g404 ( .A(n_356), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g434 ( .A(n_360), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g382 ( .A(n_367), .Y(n_382) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_379), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_378), .A2(n_382), .B1(n_383), .B2(n_387), .Y(n_381) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g395 ( .A(n_380), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g400 ( .A(n_382), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_SL g428 ( .A(n_391), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_416), .C(n_439), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_415), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B1(n_406), .B2(n_408), .C(n_411), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g440 ( .A(n_402), .B(n_428), .Y(n_440) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
OAI321xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .A3(n_421), .B1(n_423), .B2(n_424), .C(n_432), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_430), .A2(n_452), .B1(n_456), .B2(n_457), .Y(n_451) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_441), .B(n_445), .C(n_451), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_779), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_729), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_669), .B(n_728), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_461), .B(n_730), .C(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g823 ( .A(n_461), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_633), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_574), .C(n_603), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_464), .B(n_563), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_484), .B1(n_523), .B2(n_535), .Y(n_464) );
NAND2x1_ASAP7_75t_L g765 ( .A(n_465), .B(n_564), .Y(n_765) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
INVx2_ASAP7_75t_L g537 ( .A(n_467), .Y(n_537) );
INVx4_ASAP7_75t_L g579 ( .A(n_467), .Y(n_579) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_467), .Y(n_599) );
AND2x4_ASAP7_75t_L g610 ( .A(n_467), .B(n_578), .Y(n_610) );
AND2x2_ASAP7_75t_L g616 ( .A(n_467), .B(n_540), .Y(n_616) );
NOR2x1_ASAP7_75t_SL g689 ( .A(n_467), .B(n_551), .Y(n_689) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVxp67_ASAP7_75t_L g490 ( .A(n_473), .Y(n_490) );
INVx2_ASAP7_75t_L g550 ( .A(n_473), .Y(n_550) );
INVx2_ASAP7_75t_L g582 ( .A(n_476), .Y(n_582) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_476), .Y(n_596) );
INVx1_ASAP7_75t_L g607 ( .A(n_476), .Y(n_607) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_476), .Y(n_619) );
AND2x2_ASAP7_75t_L g651 ( .A(n_476), .B(n_551), .Y(n_651) );
INVx1_ASAP7_75t_L g677 ( .A(n_476), .Y(n_677) );
AND2x2_ASAP7_75t_L g739 ( .A(n_476), .B(n_567), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_503), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g632 ( .A(n_486), .B(n_571), .Y(n_632) );
INVx2_ASAP7_75t_L g674 ( .A(n_486), .Y(n_674) );
AND2x2_ASAP7_75t_L g776 ( .A(n_486), .B(n_503), .Y(n_776) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_487), .B(n_526), .Y(n_570) );
INVx2_ASAP7_75t_L g591 ( .A(n_487), .Y(n_591) );
AND2x4_ASAP7_75t_L g613 ( .A(n_487), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g648 ( .A(n_487), .Y(n_648) );
AND2x2_ASAP7_75t_L g772 ( .A(n_487), .B(n_529), .Y(n_772) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_495), .A2(n_505), .B(n_511), .Y(n_504) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_495), .A2(n_505), .B(n_511), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g746 ( .A(n_503), .Y(n_746) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_512), .Y(n_503) );
NOR2xp67_ASAP7_75t_L g621 ( .A(n_504), .B(n_591), .Y(n_621) );
AND2x2_ASAP7_75t_L g626 ( .A(n_504), .B(n_591), .Y(n_626) );
INVx2_ASAP7_75t_L g639 ( .A(n_504), .Y(n_639) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_504), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AND2x4_ASAP7_75t_L g612 ( .A(n_512), .B(n_525), .Y(n_612) );
AND2x2_ASAP7_75t_L g627 ( .A(n_512), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g682 ( .A(n_512), .Y(n_682) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_513), .B(n_529), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_513), .B(n_526), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_515), .B(n_521), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVxp33_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
INVx3_ASAP7_75t_L g588 ( .A(n_525), .Y(n_588) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_526), .Y(n_586) );
AND2x2_ASAP7_75t_L g700 ( .A(n_526), .B(n_701), .Y(n_700) );
INVx3_ASAP7_75t_L g643 ( .A(n_527), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_527), .B(n_682), .Y(n_723) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g590 ( .A(n_528), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g571 ( .A(n_529), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g614 ( .A(n_529), .Y(n_614) );
INVxp67_ASAP7_75t_L g628 ( .A(n_529), .Y(n_628) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_529), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_529), .Y(n_705) );
INVx1_ASAP7_75t_L g683 ( .A(n_535), .Y(n_683) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_536), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g725 ( .A(n_537), .B(n_566), .Y(n_725) );
OR2x2_ASAP7_75t_L g777 ( .A(n_538), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g676 ( .A(n_539), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g712 ( .A(n_539), .B(n_599), .Y(n_712) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_551), .Y(n_539) );
AND2x4_ASAP7_75t_L g566 ( .A(n_540), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g578 ( .A(n_540), .Y(n_578) );
INVx2_ASAP7_75t_L g595 ( .A(n_540), .Y(n_595) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_540), .Y(n_721) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_546), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .C(n_545), .Y(n_542) );
INVx3_ASAP7_75t_L g567 ( .A(n_551), .Y(n_567) );
INVx2_ASAP7_75t_L g661 ( .A(n_551), .Y(n_661) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_557), .B(n_562), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_565), .B(n_641), .Y(n_658) );
NOR2x1_ASAP7_75t_L g750 ( .A(n_565), .B(n_579), .Y(n_750) );
INVx4_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_566), .B(n_641), .Y(n_727) );
AND2x2_ASAP7_75t_L g594 ( .A(n_567), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g608 ( .A(n_567), .Y(n_608) );
AOI22xp5_ASAP7_75t_SL g656 ( .A1(n_568), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_569), .B(n_627), .Y(n_653) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g761 ( .A(n_570), .B(n_602), .Y(n_761) );
AND2x2_ASAP7_75t_L g584 ( .A(n_571), .B(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g620 ( .A(n_571), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g763 ( .A(n_571), .B(n_674), .Y(n_763) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g638 ( .A(n_573), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g664 ( .A(n_573), .Y(n_664) );
AND2x2_ASAP7_75t_L g699 ( .A(n_573), .B(n_591), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_583), .B1(n_587), .B2(n_592), .C(n_597), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_L g655 ( .A(n_577), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_577), .B(n_651), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_577), .B(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NOR2xp67_ASAP7_75t_SL g623 ( .A(n_579), .B(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_579), .Y(n_636) );
AND2x4_ASAP7_75t_SL g720 ( .A(n_579), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g767 ( .A(n_579), .B(n_768), .Y(n_767) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_582), .Y(n_778) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI221x1_ASAP7_75t_L g731 ( .A1(n_584), .A2(n_732), .B1(n_734), .B2(n_735), .C(n_737), .Y(n_731) );
AND2x2_ASAP7_75t_L g657 ( .A(n_585), .B(n_613), .Y(n_657) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g600 ( .A(n_588), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_588), .B(n_590), .Y(n_774) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
AND2x2_ASAP7_75t_SL g598 ( .A(n_594), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_594), .B(n_607), .Y(n_624) );
INVx2_ASAP7_75t_L g631 ( .A(n_594), .Y(n_631) );
INVx1_ASAP7_75t_L g693 ( .A(n_595), .Y(n_693) );
BUFx2_ASAP7_75t_L g713 ( .A(n_596), .Y(n_713) );
NAND2xp33_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
OR2x6_ASAP7_75t_L g630 ( .A(n_599), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g759 ( .A(n_599), .B(n_651), .Y(n_759) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_622), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_611), .B1(n_615), .B2(n_620), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
AND2x2_ASAP7_75t_SL g668 ( .A(n_606), .B(n_610), .Y(n_668) );
AND2x4_ASAP7_75t_L g734 ( .A(n_606), .B(n_692), .Y(n_734) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_607), .B(n_608), .Y(n_606) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_607), .Y(n_749) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_610), .B(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_610), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_610), .B(n_641), .Y(n_733) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g754 ( .A(n_612), .B(n_673), .Y(n_754) );
INVx3_ASAP7_75t_L g665 ( .A(n_613), .Y(n_665) );
AND2x2_ASAP7_75t_L g686 ( .A(n_613), .B(n_638), .Y(n_686) );
NAND2x1_ASAP7_75t_SL g757 ( .A(n_613), .B(n_664), .Y(n_757) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B1(n_629), .B2(n_632), .Y(n_622) );
BUFx2_ASAP7_75t_L g678 ( .A(n_624), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_625), .A2(n_716), .B1(n_725), .B2(n_726), .Y(n_724) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g681 ( .A(n_626), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g646 ( .A(n_627), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_631), .B(n_711), .C(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g666 ( .A(n_632), .Y(n_666) );
AOI211x1_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_642), .B(n_644), .C(n_662), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_637), .B(n_725), .Y(n_744) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_638), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g716 ( .A(n_638), .B(n_674), .Y(n_716) );
AND2x2_ASAP7_75t_L g771 ( .A(n_638), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g694 ( .A(n_641), .Y(n_694) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g736 ( .A(n_643), .B(n_681), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_656), .Y(n_644) );
AOI22xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_649), .B1(n_652), .B2(n_654), .Y(n_645) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g709 ( .A(n_648), .B(n_704), .Y(n_709) );
INVx1_ASAP7_75t_SL g751 ( .A(n_648), .Y(n_751) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_651), .B(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g755 ( .A(n_660), .B(n_677), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_667), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_664), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g679 ( .A(n_665), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_669), .Y(n_825) );
NAND3x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_706), .C(n_714), .Y(n_669) );
NAND4xp25_ASAP7_75t_L g780 ( .A(n_670), .B(n_706), .C(n_714), .D(n_781), .Y(n_780) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_684), .Y(n_670) );
OAI222xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .B1(n_678), .B2(n_679), .C1(n_681), .C2(n_683), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g758 ( .A1(n_676), .A2(n_759), .B(n_760), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_677), .B(n_692), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_680), .A2(n_738), .B1(n_740), .B2(n_741), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_695), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_688), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_692), .B(n_694), .Y(n_697) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_702), .B2(n_703), .Y(n_695) );
AND2x4_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_L g703 ( .A(n_699), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_707), .B(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g740 ( .A(n_709), .Y(n_740) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_724), .Y(n_714) );
AOI22xp5_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_722), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp33_ASAP7_75t_L g729 ( .A(n_728), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g824 ( .A(n_730), .Y(n_824) );
NAND3x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_742), .C(n_762), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_734), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g768 ( .A(n_739), .Y(n_768) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_752), .Y(n_742) );
AOI21xp5_ASAP7_75t_SL g743 ( .A1(n_744), .A2(n_745), .B(n_751), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_758), .Y(n_752) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_757), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_766), .B2(n_769), .C(n_773), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVxp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B(n_777), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVxp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_785), .B(n_827), .C(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_794), .Y(n_785) );
INVxp33_ASAP7_75t_L g801 ( .A(n_786), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
CKINVDCx8_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_792), .Y(n_798) );
OAI32xp33_ASAP7_75t_L g799 ( .A1(n_792), .A2(n_800), .A3(n_801), .B1(n_802), .B2(n_833), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_794), .Y(n_800) );
INVx1_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NOR2x1_ASAP7_75t_R g803 ( .A(n_797), .B(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_800), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_804), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_812), .B(n_826), .Y(n_805) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_815), .B1(n_821), .B2(n_822), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AND3x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .C(n_825), .Y(n_822) );
endmodule