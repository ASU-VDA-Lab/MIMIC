module real_jpeg_14168_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_38),
.B(n_39),
.C(n_45),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_42),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_42),
.B(n_113),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_26),
.C(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_3),
.A2(n_41),
.B1(n_62),
.B2(n_66),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_62),
.B1(n_66),
.B2(n_71),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_71),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_62),
.B1(n_66),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_9),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_97),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_12),
.A2(n_54),
.B1(n_62),
.B2(n_66),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_69),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_14),
.A2(n_62),
.B1(n_66),
.B2(n_85),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_14),
.A2(n_26),
.B1(n_33),
.B2(n_85),
.Y(n_147)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_102),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_102),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_49),
.B1(n_72),
.B2(n_73),
.Y(n_20)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_36),
.B2(n_37),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_24),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_24),
.A2(n_30),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_25),
.A2(n_29),
.B1(n_145),
.B2(n_153),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_25),
.A2(n_147),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_26),
.A2(n_33),
.B1(n_91),
.B2(n_92),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_29),
.B(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_29),
.B(n_41),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_31),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_30),
.B(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_33),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_42),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_41),
.B(n_94),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_67)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_SL g114 ( 
.A(n_43),
.B(n_64),
.C(n_66),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_59),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_59),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_61),
.B1(n_70),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_61),
.B1(n_68),
.B2(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_66),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_65),
.B(n_112),
.C(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_139),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_82),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_101),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_95),
.B(n_98),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_100),
.B1(n_107),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_100),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_89),
.A2(n_100),
.B1(n_132),
.B2(n_142),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_109),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_133),
.B(n_177),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_125),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.C(n_131),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_171),
.B(n_176),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_159),
.B(n_170),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_148),
.B(n_158),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_143),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_140),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_154),
.B(n_157),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_175),
.Y(n_176)
);


endmodule