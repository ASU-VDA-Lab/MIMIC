module fake_jpeg_10248_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_30),
.Y(n_64)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_26),
.Y(n_53)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_21),
.C(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_26),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AND2x4_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_18),
.B1(n_28),
.B2(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_30),
.B1(n_31),
.B2(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_18),
.B1(n_34),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_34),
.B1(n_20),
.B2(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_83),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_89),
.B1(n_57),
.B2(n_56),
.Y(n_120)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_84),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_17),
.B1(n_22),
.B2(n_11),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_86),
.B(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_17),
.B1(n_22),
.B2(n_10),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_10),
.C(n_16),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_8),
.C(n_15),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_22),
.B1(n_25),
.B2(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_33),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_33),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_65),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_95),
.B(n_89),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_89),
.B1(n_87),
.B2(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_60),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_121),
.C(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_106),
.Y(n_128)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_117),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_115),
.Y(n_150)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_50),
.B1(n_52),
.B2(n_67),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_58),
.C(n_62),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_19),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_22),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_68),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_123),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_80),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_146),
.C(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_135),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_144),
.B(n_110),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_72),
.B1(n_57),
.B2(n_59),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_148),
.B1(n_106),
.B2(n_100),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_89),
.B1(n_56),
.B2(n_77),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_102),
.B1(n_115),
.B2(n_96),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_101),
.B(n_110),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_123),
.B(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_15),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_66),
.B1(n_77),
.B2(n_70),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_106),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_176),
.B1(n_178),
.B2(n_127),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_97),
.B1(n_112),
.B2(n_117),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_183),
.B1(n_176),
.B2(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_169),
.Y(n_197)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_175),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_123),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_178),
.B(n_164),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_174),
.C(n_151),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_101),
.B(n_100),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_164),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_135),
.B1(n_138),
.B2(n_127),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_173),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_101),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_152),
.Y(n_175)
);

OAI22x1_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_96),
.B1(n_122),
.B2(n_22),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_78),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_181),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_136),
.B1(n_125),
.B2(n_134),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_132),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_130),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_19),
.B(n_25),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_144),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_196),
.B1(n_199),
.B2(n_206),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_7),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_201),
.C(n_205),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_25),
.B(n_8),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_140),
.B1(n_141),
.B2(n_119),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_153),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_172),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_103),
.B1(n_152),
.B2(n_145),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_163),
.C(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_210),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_22),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_103),
.B1(n_79),
.B2(n_81),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_179),
.B1(n_170),
.B2(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_168),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_158),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_211),
.B(n_217),
.C(n_221),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_224),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_165),
.B1(n_160),
.B2(n_182),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_215),
.B1(n_196),
.B2(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_160),
.B1(n_158),
.B2(n_166),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_159),
.B(n_9),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_234),
.B(n_184),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_45),
.C(n_33),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_225),
.C(n_232),
.Y(n_240)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_33),
.C(n_25),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_25),
.CI(n_1),
.CON(n_226),
.SN(n_226)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_233),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_235),
.B(n_2),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_25),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_230),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_7),
.B(n_14),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_189),
.A2(n_6),
.B(n_14),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_204),
.B1(n_195),
.B2(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_185),
.CI(n_187),
.CON(n_239),
.SN(n_239)
);

AOI321xp33_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_228),
.A3(n_222),
.B1(n_232),
.B2(n_225),
.C(n_223),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_185),
.B1(n_208),
.B2(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_6),
.C(n_13),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_236),
.C(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_215),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_254),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_15),
.B(n_12),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_248),
.A2(n_253),
.B(n_243),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_0),
.C(n_2),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_255),
.C(n_222),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_234),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_252),
.A2(n_256),
.B(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_2),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_3),
.C(n_4),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_6),
.B1(n_9),
.B2(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

BUFx12_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_221),
.B(n_226),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_248),
.B(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_266),
.C(n_245),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_256),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_212),
.C(n_4),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_267),
.C(n_254),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_3),
.B(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_3),
.C(n_5),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_247),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_283),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_285),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_284),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_238),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_279),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_244),
.B1(n_242),
.B2(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_274),
.Y(n_294)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_239),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_262),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_249),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_258),
.B(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_267),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_264),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_287),
.B(n_298),
.C(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_269),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_259),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_313),
.B1(n_305),
.B2(n_306),
.C(n_301),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_288),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_311),
.B(n_308),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_317),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.C(n_314),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_309),
.B(n_255),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_239),
.B(n_3),
.Y(n_321)
);


endmodule