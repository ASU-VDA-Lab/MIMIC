module fake_aes_4439_n_508 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_508);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_508;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g67 ( .A(n_38), .Y(n_67) );
CKINVDCx14_ASAP7_75t_R g68 ( .A(n_14), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_28), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_57), .Y(n_70) );
INVxp67_ASAP7_75t_SL g71 ( .A(n_23), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_8), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_18), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_5), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_55), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_15), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_50), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_8), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_20), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_13), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_22), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_63), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_10), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_21), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_45), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_61), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_49), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_64), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_34), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_27), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_4), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_3), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_32), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_35), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_14), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_67), .B(n_31), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g103 ( .A1(n_101), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g104 ( .A(n_101), .B(n_0), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_79), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_68), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_99), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_69), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_79), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_88), .B(n_5), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_94), .B(n_6), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_70), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_72), .B(n_6), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_92), .B(n_7), .Y(n_116) );
BUFx8_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_75), .B(n_7), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_92), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_93), .B(n_9), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_108), .B(n_67), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_124), .Y(n_130) );
AO22x2_ASAP7_75t_L g131 ( .A1(n_115), .A2(n_100), .B1(n_90), .B2(n_97), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_106), .B(n_91), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_102), .B(n_91), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_126), .Y(n_134) );
INVx4_ASAP7_75t_L g135 ( .A(n_115), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_124), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_106), .B(n_96), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_105), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_115), .B(n_74), .Y(n_140) );
INVx2_ASAP7_75t_SL g141 ( .A(n_109), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_109), .B(n_82), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
BUFx4f_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_124), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_124), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_124), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g149 ( .A(n_102), .B(n_100), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_113), .B(n_72), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_110), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_114), .B(n_74), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_114), .B(n_84), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_118), .B(n_95), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_158), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_148), .B(n_117), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_131), .A2(n_117), .B1(n_104), .B2(n_112), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_132), .B(n_127), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_141), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
BUFx8_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_144), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_133), .B(n_120), .C(n_116), .Y(n_173) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_135), .B(n_119), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_159), .B(n_127), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_137), .B(n_122), .Y(n_180) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_135), .B(n_119), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_142), .B(n_121), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_140), .B(n_122), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_135), .B(n_121), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_139), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_131), .A2(n_128), .B1(n_107), .B2(n_76), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_155), .B(n_85), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_131), .A2(n_84), .B1(n_81), .B2(n_76), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_140), .B(n_80), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_174), .B(n_149), .Y(n_200) );
NOR2x1_ASAP7_75t_L g201 ( .A(n_173), .B(n_156), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_195), .A2(n_131), .B1(n_149), .B2(n_140), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_178), .B(n_140), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_175), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_196), .A2(n_149), .B1(n_144), .B2(n_155), .Y(n_205) );
BUFx10_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_174), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_196), .A2(n_144), .B1(n_156), .B2(n_155), .Y(n_208) );
INVx1_ASAP7_75t_SL g209 ( .A(n_168), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_174), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_169), .Y(n_212) );
BUFx8_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_175), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_172), .B(n_156), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_179), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_181), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_156), .B(n_155), .C(n_154), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_181), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_167), .A2(n_157), .B(n_154), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_175), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_181), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_198), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_189), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_182), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_180), .B(n_157), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_214), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g238 ( .A1(n_212), .A2(n_191), .B1(n_103), .B2(n_165), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_213), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_196), .B1(n_162), .B2(n_163), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_233), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_233), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_214), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_202), .A2(n_192), .B1(n_176), .B2(n_186), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_209), .A2(n_177), .B1(n_188), .B2(n_184), .C(n_199), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_203), .B(n_171), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_233), .B(n_198), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_219), .B(n_203), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_202), .A2(n_199), .B1(n_182), .B2(n_183), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g250 ( .A1(n_200), .A2(n_83), .B1(n_77), .B2(n_190), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_234), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_219), .B(n_190), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_230), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_203), .B(n_171), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_217), .B(n_187), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_227), .B(n_187), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_183), .B1(n_170), .B2(n_167), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_200), .A2(n_197), .B1(n_194), .B2(n_185), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_230), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_218), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_223), .B1(n_235), .B2(n_205), .C(n_97), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_213), .B1(n_206), .B2(n_200), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_245), .A2(n_213), .B1(n_206), .B2(n_200), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g266 ( .A1(n_239), .A2(n_206), .B1(n_232), .B2(n_207), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_262), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_241), .B(n_207), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_249), .A2(n_227), .B1(n_200), .B2(n_232), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_250), .A2(n_206), .B1(n_201), .B2(n_224), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_201), .B1(n_222), .B2(n_228), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_230), .B1(n_211), .B2(n_236), .Y(n_272) );
AOI21x1_ASAP7_75t_L g273 ( .A1(n_237), .A2(n_220), .B(n_218), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_248), .A2(n_230), .B1(n_211), .B2(n_236), .Y(n_274) );
AOI222xp33_ASAP7_75t_L g275 ( .A1(n_239), .A2(n_89), .B1(n_80), .B2(n_81), .C1(n_218), .C2(n_220), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_257), .B(n_231), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_237), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_256), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_243), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_256), .A2(n_230), .B1(n_210), .B2(n_220), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_252), .A2(n_89), .B1(n_225), .B2(n_231), .C(n_221), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_246), .A2(n_230), .B1(n_236), .B2(n_211), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_257), .B(n_231), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_247), .B(n_226), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_273), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_276), .B(n_262), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_277), .B(n_243), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_278), .B(n_242), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_277), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_269), .A2(n_210), .B(n_254), .C(n_247), .Y(n_290) );
OAI22xp5_ASAP7_75t_SL g291 ( .A1(n_264), .A2(n_242), .B1(n_241), .B2(n_253), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_263), .A2(n_251), .B1(n_258), .B2(n_241), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_265), .A2(n_247), .B1(n_258), .B2(n_251), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_279), .B(n_253), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_276), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
AOI222xp33_ASAP7_75t_L g300 ( .A1(n_270), .A2(n_240), .B1(n_259), .B2(n_247), .C1(n_253), .C2(n_260), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_275), .A2(n_253), .B1(n_261), .B2(n_71), .C(n_98), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_281), .A2(n_261), .B(n_170), .Y(n_302) );
INVx3_ASAP7_75t_SL g303 ( .A(n_268), .Y(n_303) );
OAI31xp33_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_93), .A3(n_221), .B(n_211), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_283), .B(n_185), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_267), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_275), .A2(n_236), .B1(n_221), .B2(n_194), .C(n_197), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_283), .B(n_229), .Y(n_309) );
INVx4_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_297), .B(n_267), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_303), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_303), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_267), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_301), .A2(n_271), .B1(n_266), .B2(n_284), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_286), .B(n_86), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_306), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
OAI31xp33_ASAP7_75t_L g319 ( .A1(n_301), .A2(n_272), .A3(n_274), .B(n_282), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_286), .B(n_10), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_309), .B(n_86), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_308), .A2(n_221), .B1(n_226), .B2(n_229), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_288), .B(n_11), .Y(n_324) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_300), .A2(n_86), .B(n_229), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_306), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_289), .B(n_11), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_86), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_308), .A2(n_153), .B(n_136), .C(n_145), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_303), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_292), .A2(n_229), .B1(n_216), .B2(n_215), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_293), .A2(n_125), .B1(n_193), .B2(n_153), .C(n_136), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_292), .A2(n_226), .B1(n_229), .B2(n_216), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_12), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_288), .B(n_12), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_299), .B(n_13), .Y(n_338) );
AOI33xp33_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_16), .A3(n_17), .B1(n_153), .B2(n_147), .B3(n_136), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_295), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_285), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_296), .B(n_16), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_287), .B(n_17), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_287), .B(n_193), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_310), .B(n_226), .Y(n_345) );
OAI221xp5_ASAP7_75t_L g346 ( .A1(n_304), .A2(n_193), .B1(n_226), .B2(n_125), .C(n_215), .Y(n_346) );
AO21x2_ASAP7_75t_L g347 ( .A1(n_298), .A2(n_145), .B(n_147), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_293), .A2(n_226), .B1(n_229), .B2(n_216), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_337), .B(n_298), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_325), .A2(n_300), .B1(n_295), .B2(n_307), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_312), .B(n_310), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_312), .B(n_310), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_333), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_321), .B(n_298), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_325), .A2(n_290), .B(n_304), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_313), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_310), .Y(n_358) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_339), .B(n_125), .C(n_302), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_324), .B(n_291), .C(n_302), .Y(n_361) );
AND4x1_ASAP7_75t_L g362 ( .A(n_336), .B(n_309), .C(n_305), .D(n_291), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_341), .Y(n_364) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_327), .B(n_305), .C(n_307), .Y(n_365) );
AOI31xp33_ASAP7_75t_L g366 ( .A1(n_335), .A2(n_307), .A3(n_295), .B(n_24), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_316), .B(n_125), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_312), .Y(n_368) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_312), .B(n_216), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_311), .B(n_193), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_328), .B(n_19), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_313), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_328), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_314), .B(n_25), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_314), .B(n_26), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_317), .B(n_29), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_318), .B(n_30), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_318), .B(n_33), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_326), .B(n_36), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_326), .B(n_37), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_335), .A2(n_193), .B(n_147), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_340), .B(n_40), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_338), .B(n_130), .C(n_215), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_347), .Y(n_385) );
AND4x1_ASAP7_75t_L g386 ( .A(n_323), .B(n_41), .C(n_42), .D(n_44), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_330), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_340), .B(n_46), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_330), .B(n_216), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_347), .Y(n_391) );
NAND2xp33_ASAP7_75t_L g392 ( .A(n_345), .B(n_204), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_348), .B(n_47), .Y(n_393) );
AND4x1_ASAP7_75t_L g394 ( .A(n_315), .B(n_48), .C(n_51), .D(n_52), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_374), .B(n_342), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_352), .B(n_348), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_363), .B(n_342), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_357), .B(n_343), .Y(n_398) );
OAI32xp33_ASAP7_75t_L g399 ( .A1(n_351), .A2(n_345), .A3(n_320), .B1(n_346), .B2(n_334), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_349), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_365), .B(n_315), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_360), .B(n_331), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_360), .B(n_334), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_358), .B(n_344), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_356), .B(n_319), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_373), .B(n_53), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_364), .B(n_332), .Y(n_409) );
AOI32xp33_ASAP7_75t_L g410 ( .A1(n_361), .A2(n_319), .A3(n_329), .B1(n_145), .B2(n_146), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_388), .B(n_54), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_354), .B(n_56), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_383), .B(n_215), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_372), .B(n_58), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_354), .B(n_59), .Y(n_415) );
AND3x2_ASAP7_75t_L g416 ( .A(n_368), .B(n_62), .C(n_65), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_353), .B(n_66), .Y(n_417) );
AOI21xp33_ASAP7_75t_SL g418 ( .A1(n_366), .A2(n_146), .B(n_204), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_372), .B(n_204), .Y(n_419) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_383), .B(n_204), .Y(n_420) );
AND4x1_ASAP7_75t_L g421 ( .A(n_359), .B(n_215), .C(n_204), .D(n_130), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_369), .B(n_215), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_350), .B(n_130), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_375), .B(n_204), .Y(n_424) );
NAND2x2_ASAP7_75t_L g425 ( .A(n_362), .B(n_130), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_394), .B(n_130), .C(n_362), .Y(n_426) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_383), .B(n_376), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_385), .B(n_387), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_385), .B(n_387), .Y(n_429) );
AND3x2_ASAP7_75t_L g430 ( .A(n_393), .B(n_383), .C(n_355), .Y(n_430) );
AOI21xp5_ASAP7_75t_SL g431 ( .A1(n_371), .A2(n_379), .B(n_359), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_400), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_408), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_395), .B(n_375), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_405), .B(n_376), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_431), .A2(n_392), .B(n_390), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_406), .B(n_367), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_401), .B(n_394), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_428), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_427), .Y(n_440) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_430), .B(n_386), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_418), .B(n_384), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_398), .B(n_370), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_391), .Y(n_445) );
XOR2xp5_ASAP7_75t_L g446 ( .A(n_404), .B(n_371), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_425), .A2(n_393), .B1(n_389), .B2(n_379), .Y(n_447) );
OA22x2_ASAP7_75t_L g448 ( .A1(n_396), .A2(n_382), .B1(n_389), .B2(n_379), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_429), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_429), .Y(n_452) );
AOI32xp33_ASAP7_75t_L g453 ( .A1(n_411), .A2(n_379), .A3(n_378), .B1(n_377), .B2(n_380), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_403), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_426), .A2(n_384), .B1(n_378), .B2(n_380), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_399), .A2(n_381), .B(n_386), .C(n_407), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_410), .A2(n_420), .B(n_415), .C(n_412), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_424), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_413), .Y(n_460) );
XNOR2x1_ASAP7_75t_L g461 ( .A(n_416), .B(n_413), .Y(n_461) );
AO22x2_ASAP7_75t_L g462 ( .A1(n_409), .A2(n_422), .B1(n_417), .B2(n_419), .Y(n_462) );
AO22x2_ASAP7_75t_L g463 ( .A1(n_409), .A2(n_414), .B1(n_423), .B2(n_421), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
NOR3x1_ASAP7_75t_L g465 ( .A(n_401), .B(n_405), .C(n_368), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_427), .A2(n_368), .B1(n_352), .B2(n_425), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_418), .A2(n_366), .B(n_401), .C(n_250), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_406), .Y(n_468) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_430), .B(n_212), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_405), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_400), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_405), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_400), .Y(n_474) );
XOR2xp5_ASAP7_75t_L g475 ( .A(n_404), .B(n_212), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_451), .Y(n_476) );
OAI22xp33_ASAP7_75t_SL g477 ( .A1(n_468), .A2(n_440), .B1(n_465), .B2(n_436), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_452), .Y(n_478) );
O2A1O1Ixp5_ASAP7_75t_L g479 ( .A1(n_450), .A2(n_438), .B(n_459), .C(n_454), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_452), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_467), .A2(n_457), .B(n_438), .C(n_466), .Y(n_481) );
CKINVDCx6p67_ASAP7_75t_R g482 ( .A(n_475), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_461), .B(n_460), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_448), .A2(n_441), .B1(n_444), .B2(n_469), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_473), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_444), .A2(n_448), .B1(n_441), .B2(n_464), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_449), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_476), .Y(n_489) );
NOR2x1p5_ASAP7_75t_L g490 ( .A(n_482), .B(n_443), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_481), .A2(n_467), .B(n_474), .C(n_472), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_477), .A2(n_481), .B(n_483), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_484), .A2(n_455), .B1(n_458), .B2(n_460), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_487), .B(n_456), .C(n_447), .D(n_442), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_483), .A2(n_471), .B1(n_470), .B2(n_434), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_494), .A2(n_492), .B1(n_493), .B2(n_487), .Y(n_496) );
NAND4xp25_ASAP7_75t_SL g497 ( .A(n_491), .B(n_490), .C(n_453), .D(n_495), .Y(n_497) );
OAI222xp33_ASAP7_75t_L g498 ( .A1(n_489), .A2(n_488), .B1(n_486), .B2(n_485), .C1(n_446), .C2(n_433), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g499 ( .A1(n_491), .A2(n_479), .B(n_488), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_497), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_496), .A2(n_462), .B1(n_478), .B2(n_437), .Y(n_501) );
NAND3xp33_ASAP7_75t_SL g502 ( .A(n_498), .B(n_478), .C(n_480), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_500), .A2(n_499), .B1(n_463), .B2(n_462), .Y(n_503) );
XOR2xp5_ASAP7_75t_L g504 ( .A(n_501), .B(n_462), .Y(n_504) );
AOI22xp5_ASAP7_75t_SL g505 ( .A1(n_504), .A2(n_502), .B1(n_435), .B2(n_449), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_505), .A2(n_503), .B1(n_463), .B2(n_445), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_506), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_507), .A2(n_463), .B(n_439), .Y(n_508) );
endmodule