module fake_jpeg_1618_n_224 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_224);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_92),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_71),
.B1(n_74),
.B2(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_68),
.B1(n_76),
.B2(n_59),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_113),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_73),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_87),
.B1(n_71),
.B2(n_74),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_141)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_77),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_4),
.C(n_5),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_83),
.B1(n_58),
.B2(n_62),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_51),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_67),
.B1(n_78),
.B2(n_75),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_75),
.B1(n_67),
.B2(n_78),
.Y(n_118)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_73),
.B1(n_72),
.B2(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_104),
.B1(n_115),
.B2(n_6),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_60),
.A3(n_67),
.B1(n_75),
.B2(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_109),
.B(n_108),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_131),
.B(n_136),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_80),
.B(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_135),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_60),
.B(n_64),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_1),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_1),
.B(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_138),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_8),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_130),
.C(n_139),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_157),
.C(n_15),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_117),
.B(n_119),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_35),
.B(n_32),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_164),
.Y(n_179)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_154),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_150),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_115),
.C(n_40),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_18),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_19),
.B(n_20),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_24),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_178),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_173),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_151),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_176),
.B(n_177),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_28),
.B(n_27),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_16),
.B(n_17),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_26),
.B(n_23),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_21),
.B(n_171),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_185),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_154),
.C(n_163),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_19),
.B1(n_21),
.B2(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_142),
.B1(n_157),
.B2(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_166),
.B1(n_165),
.B2(n_22),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_191),
.A2(n_179),
.B1(n_172),
.B2(n_167),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_194),
.Y(n_201)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_175),
.B(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_175),
.C(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_206),
.C(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_185),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_188),
.B1(n_192),
.B2(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_190),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_189),
.B(n_203),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_189),
.C(n_194),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_217),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_212),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_169),
.B(n_184),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_204),
.C(n_201),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_168),
.CI(n_200),
.CON(n_224),
.SN(n_224)
);


endmodule