module real_aes_14515_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_954;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
OA21x2_ASAP7_75t_L g141 ( .A1(n_0), .A2(n_51), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g254 ( .A(n_0), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_1), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g296 ( .A(n_2), .B(n_212), .Y(n_296) );
NAND2xp33_ASAP7_75t_L g646 ( .A(n_3), .B(n_210), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_4), .A2(n_98), .B1(n_181), .B2(n_230), .C(n_250), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_5), .A2(n_124), .B1(n_568), .B2(n_569), .Y(n_123) );
INVx1_ASAP7_75t_L g568 ( .A(n_5), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_5), .A2(n_101), .B1(n_954), .B2(n_956), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_6), .B(n_197), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_7), .B(n_657), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_8), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_9), .B(n_146), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_10), .B(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_11), .Y(n_650) );
BUFx3_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g159 ( .A(n_12), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_13), .B(n_161), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_14), .A2(n_187), .B(n_635), .C(n_636), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g949 ( .A1(n_15), .A2(n_54), .B1(n_950), .B2(n_951), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_15), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_16), .Y(n_239) );
BUFx10_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_18), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_19), .B(n_286), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_20), .B(n_180), .Y(n_179) );
OAI21xp33_ASAP7_75t_L g257 ( .A1(n_21), .A2(n_68), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_21), .B(n_169), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_22), .B(n_284), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_23), .A2(n_626), .B(n_627), .C(n_629), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_24), .B(n_680), .Y(n_679) );
O2A1O1Ixp5_ASAP7_75t_L g262 ( .A1(n_25), .A2(n_186), .B(n_188), .C(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g711 ( .A(n_26), .B(n_197), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_27), .B(n_169), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_28), .A2(n_79), .B1(n_146), .B2(n_150), .Y(n_659) );
INVx1_ASAP7_75t_L g167 ( .A(n_29), .Y(n_167) );
INVx1_ASAP7_75t_L g620 ( .A(n_30), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_31), .B(n_151), .Y(n_242) );
XOR2xp5_ASAP7_75t_L g947 ( .A(n_32), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g468 ( .A(n_33), .Y(n_468) );
NAND2xp33_ASAP7_75t_L g528 ( .A(n_33), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_33), .A2(n_565), .B(n_567), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_34), .B(n_150), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_35), .B(n_169), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_36), .B(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
AND3x2_ASAP7_75t_L g955 ( .A(n_37), .B(n_585), .C(n_586), .Y(n_955) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_38), .B(n_181), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_39), .B(n_169), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_40), .B(n_186), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_41), .B(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_42), .Y(n_637) );
AND2x4_ASAP7_75t_L g166 ( .A(n_43), .B(n_167), .Y(n_166) );
NAND2x1_ASAP7_75t_L g211 ( .A(n_44), .B(n_212), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_45), .Y(n_246) );
INVx1_ASAP7_75t_L g206 ( .A(n_46), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_47), .Y(n_278) );
AND2x2_ASAP7_75t_L g295 ( .A(n_48), .B(n_157), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_49), .B(n_150), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_50), .A2(n_93), .B1(n_150), .B2(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g255 ( .A(n_51), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_52), .B(n_197), .Y(n_288) );
INVx1_ASAP7_75t_L g142 ( .A(n_53), .Y(n_142) );
INVx1_ASAP7_75t_L g951 ( .A(n_54), .Y(n_951) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_55), .B(n_157), .Y(n_302) );
AND2x4_ASAP7_75t_L g109 ( .A(n_56), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_57), .B(n_169), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_58), .B(n_210), .Y(n_209) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_59), .B(n_81), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_60), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g685 ( .A(n_61), .B(n_170), .Y(n_685) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_63), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_64), .B(n_680), .Y(n_718) );
NAND2x1_ASAP7_75t_L g698 ( .A(n_65), .B(n_635), .Y(n_698) );
AND2x2_ASAP7_75t_L g300 ( .A(n_66), .B(n_197), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_67), .B(n_161), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_68), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_69), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_70), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_71), .B(n_150), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_72), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_73), .A2(n_100), .B1(n_126), .B2(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_74), .B(n_275), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_75), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g119 ( .A(n_76), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_77), .B(n_178), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_78), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_80), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_82), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_83), .B(n_181), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_84), .B(n_170), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_85), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_86), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_87), .B(n_286), .Y(n_695) );
NAND2xp33_ASAP7_75t_SL g615 ( .A(n_88), .B(n_245), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_89), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_90), .B(n_157), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_91), .B(n_180), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_92), .B(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g154 ( .A(n_94), .Y(n_154) );
BUFx3_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
INVx1_ASAP7_75t_L g189 ( .A(n_94), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_95), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_96), .B(n_247), .Y(n_683) );
NAND2xp33_ASAP7_75t_L g643 ( .A(n_97), .B(n_207), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_99), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_102), .B(n_157), .Y(n_715) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_111), .B(n_578), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g957 ( .A(n_106), .B(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_109), .B(n_115), .Y(n_590) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_123), .B(n_570), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
CKINVDCx11_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx3_ASAP7_75t_L g574 ( .A(n_115), .Y(n_574) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_116), .Y(n_577) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g588 ( .A(n_117), .Y(n_588) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_117), .Y(n_960) );
NOR2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g586 ( .A(n_119), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
BUFx2_ASAP7_75t_L g597 ( .A(n_121), .Y(n_597) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_122), .Y(n_585) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_124), .Y(n_569) );
XNOR2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_128), .A2(n_593), .B(n_598), .Y(n_592) );
OA21x2_ASAP7_75t_L g952 ( .A1(n_128), .A2(n_593), .B(n_598), .Y(n_952) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_469), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_385), .B(n_468), .Y(n_129) );
NOR2xp67_ASAP7_75t_SL g470 ( .A(n_130), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_352), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_317), .C(n_342), .Y(n_131) );
OAI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_214), .B1(n_289), .B2(n_309), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_133), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_172), .Y(n_134) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_135), .Y(n_308) );
INVx1_ASAP7_75t_L g351 ( .A(n_135), .Y(n_351) );
AND2x2_ASAP7_75t_L g391 ( .A(n_135), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g412 ( .A(n_135), .B(n_173), .Y(n_412) );
INVx1_ASAP7_75t_L g535 ( .A(n_135), .Y(n_535) );
INVx1_ASAP7_75t_L g542 ( .A(n_135), .Y(n_542) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g383 ( .A(n_136), .B(n_193), .Y(n_383) );
AND2x2_ASAP7_75t_L g447 ( .A(n_136), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g475 ( .A(n_136), .B(n_434), .Y(n_475) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g403 ( .A(n_137), .Y(n_403) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_143), .B(n_168), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_139), .A2(n_165), .B(n_619), .Y(n_622) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g258 ( .A(n_140), .Y(n_258) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
INVxp33_ASAP7_75t_L g621 ( .A(n_141), .Y(n_621) );
INVx1_ASAP7_75t_L g256 ( .A(n_142), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_155), .B(n_165), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B(n_152), .Y(n_144) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g247 ( .A(n_147), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_147), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g275 ( .A(n_147), .Y(n_275) );
INVx2_ASAP7_75t_L g284 ( .A(n_147), .Y(n_284) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_148), .Y(n_162) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
INVx2_ASAP7_75t_L g210 ( .A(n_151), .Y(n_210) );
INVx2_ASAP7_75t_L g241 ( .A(n_151), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_152), .A2(n_177), .B(n_179), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_152), .A2(n_228), .B(n_231), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_152), .A2(n_282), .B(n_285), .Y(n_281) );
AO21x1_ASAP7_75t_L g611 ( .A1(n_152), .A2(n_612), .B(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_152), .A2(n_670), .B(n_672), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_152), .A2(n_694), .B(n_695), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_152), .A2(n_717), .B(n_718), .Y(n_716) );
BUFx10_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g250 ( .A(n_154), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B(n_163), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx1_ASAP7_75t_L g207 ( .A(n_158), .Y(n_207) );
INVx2_ASAP7_75t_L g245 ( .A(n_158), .Y(n_245) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx3_ASAP7_75t_L g212 ( .A(n_162), .Y(n_212) );
INVx2_ASAP7_75t_L g617 ( .A(n_162), .Y(n_617) );
INVx2_ASAP7_75t_L g657 ( .A(n_162), .Y(n_657) );
INVx2_ASAP7_75t_L g680 ( .A(n_162), .Y(n_680) );
AO21x1_ASAP7_75t_L g614 ( .A1(n_163), .A2(n_615), .B(n_616), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_163), .A2(n_667), .B(n_668), .Y(n_666) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g201 ( .A(n_164), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_164), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g243 ( .A(n_164), .Y(n_243) );
AOI211x1_ASAP7_75t_L g712 ( .A1(n_164), .A2(n_711), .B(n_713), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_199), .B(n_208), .Y(n_198) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_165), .A2(n_641), .B(n_644), .Y(n_640) );
OAI21x1_ASAP7_75t_L g665 ( .A1(n_165), .A2(n_666), .B(n_669), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_165), .A2(n_710), .B(n_711), .Y(n_709) );
BUFx6f_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g233 ( .A(n_166), .Y(n_233) );
INVx1_ASAP7_75t_L g252 ( .A(n_166), .Y(n_252) );
INVx3_ASAP7_75t_L g265 ( .A(n_166), .Y(n_265) );
INVx1_ASAP7_75t_L g654 ( .A(n_166), .Y(n_654) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_170), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g440 ( .A(n_172), .Y(n_440) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_192), .Y(n_172) );
INVx1_ASAP7_75t_L g325 ( .A(n_173), .Y(n_325) );
INVx3_ASAP7_75t_L g347 ( .A(n_173), .Y(n_347) );
INVx1_ASAP7_75t_L g372 ( .A(n_173), .Y(n_372) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_173), .Y(n_384) );
OR2x2_ASAP7_75t_L g405 ( .A(n_173), .B(n_293), .Y(n_405) );
AND2x2_ASAP7_75t_L g481 ( .A(n_173), .B(n_292), .Y(n_481) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_183), .B(n_190), .Y(n_175) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g626 ( .A(n_181), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_181), .B(n_637), .Y(n_636) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g230 ( .A(n_182), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .Y(n_183) );
AOI21x1_ASAP7_75t_L g208 ( .A1(n_187), .A2(n_209), .B(n_211), .Y(n_208) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx3_ASAP7_75t_L g298 ( .A(n_189), .Y(n_298) );
INVxp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_193), .B(n_293), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_193), .Y(n_324) );
INVx1_ASAP7_75t_L g350 ( .A(n_193), .Y(n_350) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_193), .B(n_292), .Y(n_427) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_193), .Y(n_437) );
INVx2_ASAP7_75t_L g448 ( .A(n_193), .Y(n_448) );
AND2x2_ASAP7_75t_L g486 ( .A(n_193), .B(n_403), .Y(n_486) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_198), .B(n_213), .Y(n_194) );
INVx1_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_197), .Y(n_220) );
INVxp33_ASAP7_75t_L g306 ( .A(n_197), .Y(n_306) );
INVx1_ASAP7_75t_L g336 ( .A(n_197), .Y(n_336) );
NOR2xp67_ASAP7_75t_SL g676 ( .A(n_197), .B(n_252), .Y(n_676) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_197), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_202), .B(n_204), .Y(n_199) );
INVx1_ASAP7_75t_L g629 ( .A(n_201), .Y(n_629) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
INVx1_ASAP7_75t_L g225 ( .A(n_210), .Y(n_225) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_268), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_235), .Y(n_216) );
INVx2_ASAP7_75t_L g456 ( .A(n_217), .Y(n_456) );
INVxp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_221), .B(n_234), .Y(n_218) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_219), .A2(n_272), .B(n_288), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_219), .A2(n_221), .B(n_234), .Y(n_330) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_219), .A2(n_272), .B(n_288), .Y(n_341) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_219), .A2(n_665), .B(n_673), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_219), .A2(n_665), .B(n_673), .Y(n_688) );
OAI21x1_ASAP7_75t_L g691 ( .A1(n_219), .A2(n_692), .B(n_699), .Y(n_691) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_227), .B(n_232), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_226), .Y(n_222) );
INVx1_ASAP7_75t_L g655 ( .A(n_226), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_229), .A2(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_230), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g635 ( .A(n_230), .Y(n_635) );
INVx2_ASAP7_75t_L g671 ( .A(n_230), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_232), .A2(n_693), .B(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_SL g287 ( .A(n_233), .Y(n_287) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g314 ( .A(n_236), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g357 ( .A(n_236), .B(n_316), .Y(n_357) );
INVx1_ASAP7_75t_L g457 ( .A(n_236), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_257), .C(n_259), .Y(n_236) );
AND2x4_ASAP7_75t_L g339 ( .A(n_237), .B(n_340), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .C(n_251), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .C(n_243), .Y(n_238) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_243), .A2(n_642), .B(n_643), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_243), .A2(n_683), .B(n_684), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B1(n_247), .B2(n_248), .C(n_249), .Y(n_244) );
INVx2_ASAP7_75t_L g286 ( .A(n_245), .Y(n_286) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_274), .B1(n_276), .B2(n_280), .Y(n_273) );
INVx2_ASAP7_75t_SL g279 ( .A(n_250), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g267 ( .A(n_253), .Y(n_267) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_256), .Y(n_253) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_254), .A2(n_255), .B(n_256), .Y(n_333) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_258), .A2(n_640), .B(n_647), .Y(n_639) );
NAND2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_266), .Y(n_259) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_260), .A2(n_333), .B(n_334), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .C(n_265), .Y(n_260) );
INVx2_ASAP7_75t_L g307 ( .A(n_265), .Y(n_307) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_267), .B(n_653), .C(n_655), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_267), .B(n_298), .C(n_653), .Y(n_658) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g520 ( .A(n_269), .Y(n_520) );
AND2x4_ASAP7_75t_L g550 ( .A(n_269), .B(n_328), .Y(n_550) );
BUFx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g379 ( .A(n_270), .B(n_339), .Y(n_379) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_281), .B(n_287), .Y(n_272) );
O2A1O1Ixp5_ASAP7_75t_L g696 ( .A1(n_274), .A2(n_298), .B(n_697), .C(n_698), .Y(n_696) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_287), .B(n_333), .Y(n_630) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_308), .Y(n_290) );
INVx1_ASAP7_75t_L g439 ( .A(n_291), .Y(n_439) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_293), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g434 ( .A(n_293), .Y(n_434) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .B(n_305), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g304 ( .A(n_298), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g305 ( .A1(n_300), .A2(n_306), .B(n_307), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_304), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_304), .A2(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g373 ( .A(n_308), .Y(n_373) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2x1p5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVx1_ASAP7_75t_L g502 ( .A(n_311), .Y(n_502) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g398 ( .A(n_312), .B(n_331), .Y(n_398) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g344 ( .A(n_313), .B(n_332), .Y(n_344) );
INVx1_ASAP7_75t_L g458 ( .A(n_314), .Y(n_458) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g408 ( .A(n_316), .Y(n_408) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_316), .Y(n_449) );
AND2x2_ASAP7_75t_L g487 ( .A(n_316), .B(n_398), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_316), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_326), .Y(n_317) );
NOR2xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_322), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g459 ( .A(n_320), .B(n_371), .Y(n_459) );
AND2x2_ASAP7_75t_L g495 ( .A(n_320), .B(n_325), .Y(n_495) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g392 ( .A(n_321), .Y(n_392) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_323), .B(n_346), .Y(n_522) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g474 ( .A(n_324), .B(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g479 ( .A(n_324), .Y(n_479) );
OR2x2_ASAP7_75t_L g537 ( .A(n_324), .B(n_372), .Y(n_537) );
AND2x2_ASAP7_75t_L g451 ( .A(n_325), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g511 ( .A(n_325), .B(n_447), .Y(n_511) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_327), .A2(n_359), .B1(n_561), .B2(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_337), .Y(n_327) );
AND2x2_ASAP7_75t_L g525 ( .A(n_328), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g367 ( .A(n_329), .Y(n_367) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g360 ( .A(n_330), .B(n_332), .Y(n_360) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_331), .Y(n_376) );
AND2x2_ASAP7_75t_L g546 ( .A(n_331), .B(n_397), .Y(n_546) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g443 ( .A(n_332), .Y(n_443) );
INVx2_ASAP7_75t_L g632 ( .A(n_333), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_333), .B(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_R g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x4_ASAP7_75t_SL g418 ( .A(n_337), .B(n_398), .Y(n_418) );
AND2x2_ASAP7_75t_L g421 ( .A(n_337), .B(n_344), .Y(n_421) );
AND2x2_ASAP7_75t_L g441 ( .A(n_337), .B(n_360), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_337), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_337), .B(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
INVx1_ASAP7_75t_L g397 ( .A(n_339), .Y(n_397) );
AND2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_341), .Y(n_424) );
INVx1_ASAP7_75t_L g363 ( .A(n_341), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_344), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g414 ( .A(n_344), .B(n_361), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_344), .B(n_379), .Y(n_416) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g553 ( .A(n_346), .Y(n_553) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g433 ( .A(n_347), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g353 ( .A(n_348), .Y(n_353) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
OR2x2_ASAP7_75t_L g516 ( .A(n_349), .B(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_350), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_364), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_356), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g365 ( .A(n_357), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AND2x2_ASAP7_75t_L g423 ( .A(n_360), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g482 ( .A(n_360), .B(n_408), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_360), .A2(n_484), .B1(n_486), .B2(n_487), .Y(n_483) );
AND2x2_ASAP7_75t_L g505 ( .A(n_360), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g519 ( .A(n_360), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g445 ( .A(n_361), .Y(n_445) );
AND2x2_ASAP7_75t_L g498 ( .A(n_361), .B(n_398), .Y(n_498) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g506 ( .A(n_362), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_374), .B2(n_380), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g530 ( .A1(n_365), .A2(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g476 ( .A(n_366), .B(n_424), .Y(n_476) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g497 ( .A(n_371), .B(n_447), .Y(n_497) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_373), .B(n_439), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g491 ( .A(n_383), .B(n_405), .Y(n_491) );
AND2x2_ASAP7_75t_L g426 ( .A(n_384), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_428), .Y(n_386) );
NOR4xp25_ASAP7_75t_L g527 ( .A(n_387), .B(n_428), .C(n_528), .D(n_551), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_417), .Y(n_387) );
NOR3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_409), .C(n_415), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_390), .B(n_399), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_392), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_395), .B(n_456), .Y(n_490) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_396), .Y(n_559) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_406), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
AND2x2_ASAP7_75t_L g507 ( .A(n_402), .B(n_427), .Y(n_507) );
INVx1_ASAP7_75t_L g517 ( .A(n_402), .Y(n_517) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_402), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g452 ( .A(n_403), .B(n_448), .Y(n_452) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g467 ( .A(n_405), .Y(n_467) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g494 ( .A(n_408), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_412), .B(n_463), .Y(n_549) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_425), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_423), .A2(n_431), .B1(n_438), .B2(n_441), .Y(n_430) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g464 ( .A(n_427), .Y(n_464) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_453), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_442), .Y(n_429) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_432), .B(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_432), .B(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_433), .B(n_534), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g541 ( .A(n_433), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g513 ( .A(n_443), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_449), .B2(n_450), .Y(n_444) );
AND2x2_ASAP7_75t_L g499 ( .A(n_447), .B(n_467), .Y(n_499) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_452), .B(n_481), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_460), .Y(n_453) );
OAI21xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B(n_459), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_455), .A2(n_461), .B1(n_462), .B2(n_465), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_455), .A2(n_533), .B(n_536), .Y(n_532) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_456), .B(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x2_ASAP7_75t_L g563 ( .A(n_467), .B(n_556), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_527), .B(n_564), .Y(n_469) );
INVx1_ASAP7_75t_L g567 ( .A(n_471), .Y(n_567) );
NAND4xp75_ASAP7_75t_L g471 ( .A(n_472), .B(n_488), .C(n_503), .D(n_514), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .B1(n_477), .B2(n_482), .Y(n_473) );
INVx2_ASAP7_75t_L g531 ( .A(n_474), .Y(n_531) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_492), .B2(n_495), .Y(n_489) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_495), .B(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_498), .A2(n_505), .B(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_508), .Y(n_503) );
INVx1_ASAP7_75t_L g526 ( .A(n_506), .Y(n_526) );
AOI21xp5_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_510), .B(n_512), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
OAI21xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_518), .B(n_521), .Y(n_515) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_520), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g566 ( .A(n_529), .Y(n_566) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_538), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B(n_547), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g556 ( .A(n_542), .Y(n_556) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g558 ( .A(n_550), .B(n_559), .Y(n_558) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_551), .B(n_566), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_557), .B(n_560), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_574), .B(n_959), .Y(n_958) );
NOR2x1_ASAP7_75t_SL g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_591), .B(n_953), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx12f_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_587), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AND2x2_ASAP7_75t_L g954 ( .A(n_587), .B(n_955), .Y(n_954) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_946), .B1(n_947), .B2(n_952), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx11_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx8_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_SL g601 ( .A(n_596), .Y(n_601) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_600), .Y(n_599) );
CKINVDCx10_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AND3x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_842), .C(n_908), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_760), .C(n_816), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_733), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_660), .B1(n_700), .B2(n_720), .C1(n_726), .C2(n_731), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_638), .Y(n_607) );
AND2x2_ASAP7_75t_L g875 ( .A(n_608), .B(n_876), .Y(n_875) );
AND2x4_ASAP7_75t_SL g885 ( .A(n_608), .B(n_742), .Y(n_885) );
INVx1_ASAP7_75t_L g900 ( .A(n_608), .Y(n_900) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_623), .Y(n_608) );
AND2x2_ASAP7_75t_L g832 ( .A(n_609), .B(n_732), .Y(n_832) );
INVx1_ASAP7_75t_L g907 ( .A(n_609), .Y(n_907) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g738 ( .A(n_610), .Y(n_738) );
OR2x2_ASAP7_75t_L g740 ( .A(n_610), .B(n_724), .Y(n_740) );
AND2x2_ASAP7_75t_L g765 ( .A(n_610), .B(n_639), .Y(n_765) );
AND2x2_ASAP7_75t_L g790 ( .A(n_610), .B(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g806 ( .A(n_610), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g847 ( .A(n_610), .B(n_724), .Y(n_847) );
AO31x2_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_614), .A3(n_618), .B(n_622), .Y(n_610) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g784 ( .A(n_623), .B(n_785), .Y(n_784) );
BUFx2_ASAP7_75t_L g795 ( .A(n_623), .Y(n_795) );
INVx1_ASAP7_75t_L g807 ( .A(n_623), .Y(n_807) );
INVx1_ASAP7_75t_L g830 ( .A(n_623), .Y(n_830) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_623), .Y(n_918) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_624), .B(n_633), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_624), .B(n_633), .Y(n_724) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_630), .B(n_631), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_629), .A2(n_645), .B(n_646), .Y(n_644) );
OR2x2_ASAP7_75t_L g633 ( .A(n_630), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g736 ( .A(n_638), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g841 ( .A(n_638), .Y(n_841) );
AND2x2_ASAP7_75t_L g911 ( .A(n_638), .B(n_794), .Y(n_911) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_648), .Y(n_638) );
INVx1_ASAP7_75t_L g725 ( .A(n_639), .Y(n_725) );
AND2x2_ASAP7_75t_L g731 ( .A(n_639), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g755 ( .A(n_639), .Y(n_755) );
INVx1_ASAP7_75t_L g791 ( .A(n_639), .Y(n_791) );
AND2x2_ASAP7_75t_L g874 ( .A(n_639), .B(n_723), .Y(n_874) );
INVx1_ASAP7_75t_L g721 ( .A(n_648), .Y(n_721) );
INVx1_ASAP7_75t_L g732 ( .A(n_648), .Y(n_732) );
AND2x2_ASAP7_75t_L g742 ( .A(n_648), .B(n_725), .Y(n_742) );
AND2x2_ASAP7_75t_L g766 ( .A(n_648), .B(n_724), .Y(n_766) );
INVx1_ASAP7_75t_L g772 ( .A(n_648), .Y(n_772) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_648), .Y(n_788) );
INVxp67_ASAP7_75t_L g846 ( .A(n_648), .Y(n_846) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_656), .B1(n_658), .B2(n_659), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_686), .Y(n_661) );
OAI31xp33_ASAP7_75t_L g817 ( .A1(n_662), .A2(n_818), .A3(n_823), .B(n_827), .Y(n_817) );
AND2x4_ASAP7_75t_L g882 ( .A(n_662), .B(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_662), .B(n_746), .Y(n_904) );
INVx4_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2x1_ASAP7_75t_L g872 ( .A(n_663), .B(n_706), .Y(n_872) );
OR2x2_ASAP7_75t_L g923 ( .A(n_663), .B(n_826), .Y(n_923) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_674), .Y(n_663) );
INVx2_ASAP7_75t_L g730 ( .A(n_664), .Y(n_730) );
INVx2_ASAP7_75t_L g704 ( .A(n_674), .Y(n_704) );
AND2x2_ASAP7_75t_L g729 ( .A(n_674), .B(n_730), .Y(n_729) );
AND2x4_ASAP7_75t_L g749 ( .A(n_674), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g779 ( .A(n_674), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_674), .B(n_752), .Y(n_811) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_681), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_676), .A2(n_682), .B(n_685), .Y(n_681) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g850 ( .A(n_687), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_687), .B(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g703 ( .A(n_688), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g852 ( .A(n_688), .B(n_708), .Y(n_852) );
INVx2_ASAP7_75t_L g775 ( .A(n_689), .Y(n_775) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g719 ( .A(n_690), .Y(n_719) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g752 ( .A(n_691), .Y(n_752) );
INVx1_ASAP7_75t_L g799 ( .A(n_691), .Y(n_799) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g857 ( .A(n_702), .Y(n_857) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_703), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_703), .B(n_775), .Y(n_774) );
AND2x4_ASAP7_75t_SL g801 ( .A(n_704), .B(n_802), .Y(n_801) );
OR2x2_ASAP7_75t_L g815 ( .A(n_704), .B(n_785), .Y(n_815) );
AND2x2_ASAP7_75t_L g894 ( .A(n_704), .B(n_708), .Y(n_894) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g777 ( .A(n_706), .B(n_778), .Y(n_777) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_719), .Y(n_706) );
AND2x2_ASAP7_75t_L g944 ( .A(n_707), .B(n_719), .Y(n_944) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g728 ( .A(n_708), .B(n_719), .Y(n_728) );
BUFx2_ASAP7_75t_L g746 ( .A(n_708), .Y(n_746) );
INVx1_ASAP7_75t_L g750 ( .A(n_708), .Y(n_750) );
INVx2_ASAP7_75t_L g785 ( .A(n_708), .Y(n_785) );
INVx2_ASAP7_75t_L g802 ( .A(n_708), .Y(n_802) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_708), .Y(n_935) );
OR2x6_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_719), .Y(n_861) );
AND2x2_ASAP7_75t_L g926 ( .A(n_720), .B(n_907), .Y(n_926) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx2_ASAP7_75t_L g876 ( .A(n_721), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_721), .B(n_907), .Y(n_937) );
INVx1_ASAP7_75t_L g813 ( .A(n_722), .Y(n_813) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g771 ( .A(n_724), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVxp67_ASAP7_75t_L g927 ( .A(n_728), .Y(n_927) );
AND2x2_ASAP7_75t_L g834 ( .A(n_729), .B(n_810), .Y(n_834) );
INVx2_ASAP7_75t_L g862 ( .A(n_729), .Y(n_862) );
AND2x2_ASAP7_75t_L g751 ( .A(n_730), .B(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g822 ( .A(n_730), .B(n_799), .Y(n_822) );
INVx1_ASAP7_75t_L g838 ( .A(n_730), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_731), .B(n_806), .Y(n_812) );
AND2x2_ASAP7_75t_L g866 ( .A(n_731), .B(n_830), .Y(n_866) );
AOI21xp33_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_743), .B(n_747), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_739), .Y(n_734) );
INVx2_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_738), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_738), .B(n_755), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_739), .A2(n_748), .B1(n_753), .B2(n_757), .Y(n_747) );
OR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g756 ( .A(n_740), .Y(n_756) );
OR2x2_ASAP7_75t_L g888 ( .A(n_740), .B(n_841), .Y(n_888) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g905 ( .A(n_742), .B(n_906), .Y(n_905) );
AND2x2_ASAP7_75t_L g917 ( .A(n_742), .B(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g889 ( .A(n_745), .B(n_862), .Y(n_889) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
AND2x2_ASAP7_75t_L g758 ( .A(n_749), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_749), .B(n_850), .Y(n_849) );
AND2x2_ASAP7_75t_L g877 ( .A(n_749), .B(n_878), .Y(n_877) );
AND2x2_ASAP7_75t_L g897 ( .A(n_749), .B(n_861), .Y(n_897) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_750), .Y(n_899) );
INVx1_ASAP7_75t_L g782 ( .A(n_751), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_751), .B(n_935), .Y(n_934) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_752), .Y(n_759) );
INVx1_ASAP7_75t_L g826 ( .A(n_752), .Y(n_826) );
AND2x2_ASAP7_75t_L g837 ( .A(n_752), .B(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx2_ASAP7_75t_L g805 ( .A(n_754), .Y(n_805) );
AND2x2_ASAP7_75t_L g831 ( .A(n_754), .B(n_832), .Y(n_831) );
BUFx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_755), .Y(n_769) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_792), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_773), .B(n_776), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .Y(n_762) );
OAI22xp33_ASAP7_75t_SL g859 ( .A1(n_763), .A2(n_809), .B1(n_860), .B2(n_863), .Y(n_859) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
AND2x2_ASAP7_75t_L g851 ( .A(n_766), .B(n_790), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g884 ( .A1(n_766), .A2(n_773), .B1(n_882), .B2(n_885), .C(n_886), .Y(n_884) );
OR2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_770), .Y(n_767) );
OR2x2_ASAP7_75t_L g863 ( .A(n_770), .B(n_789), .Y(n_863) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g800 ( .A(n_775), .B(n_801), .Y(n_800) );
OR2x2_ASAP7_75t_L g814 ( .A(n_775), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g883 ( .A(n_775), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_780), .B(n_786), .Y(n_776) );
INVx1_ASAP7_75t_L g797 ( .A(n_778), .Y(n_797) );
AND2x4_ASAP7_75t_SL g855 ( .A(n_778), .B(n_821), .Y(n_855) );
INVx4_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
AOI311xp33_ASAP7_75t_L g890 ( .A1(n_782), .A2(n_891), .A3(n_892), .B(n_895), .C(n_902), .Y(n_890) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
BUFx3_ASAP7_75t_L g810 ( .A(n_785), .Y(n_810) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
OR2x2_ASAP7_75t_L g856 ( .A(n_787), .B(n_789), .Y(n_856) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OR2x2_ASAP7_75t_L g887 ( .A(n_789), .B(n_829), .Y(n_887) );
INVx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g793 ( .A(n_790), .B(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g921 ( .A(n_790), .B(n_829), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_796), .B1(n_800), .B2(n_803), .C(n_808), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_793), .B(n_876), .Y(n_945) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g833 ( .A1(n_795), .A2(n_834), .B(n_835), .C(n_840), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_797), .B(n_825), .Y(n_824) );
BUFx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_801), .B(n_940), .Y(n_939) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g901 ( .A(n_805), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx2_ASAP7_75t_L g820 ( .A(n_810), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_810), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g915 ( .A(n_811), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_812), .A2(n_854), .B1(n_856), .B2(n_857), .Y(n_853) );
INVx2_ASAP7_75t_L g839 ( .A(n_815), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g816 ( .A(n_817), .B(n_833), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g870 ( .A(n_822), .Y(n_870) );
INVx2_ASAP7_75t_SL g878 ( .A(n_822), .Y(n_878) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_822), .Y(n_940) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NAND2x1p5_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_830), .Y(n_930) );
INVx1_ASAP7_75t_L g880 ( .A(n_831), .Y(n_880) );
AND2x4_ASAP7_75t_L g873 ( .A(n_832), .B(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_839), .Y(n_836) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AND4x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_858), .C(n_884), .D(n_890), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_848), .B1(n_851), .B2(n_852), .C(n_853), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
AOI21xp33_ASAP7_75t_L g941 ( .A1(n_849), .A2(n_942), .B(n_945), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_850), .B(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g920 ( .A(n_856), .Y(n_920) );
NOR3xp33_ASAP7_75t_SL g858 ( .A(n_859), .B(n_864), .C(n_879), .Y(n_858) );
OR2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_867), .B(n_871), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B1(n_875), .B2(n_877), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AOI21xp33_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B(n_889), .Y(n_886) );
INVx2_ASAP7_75t_L g891 ( .A(n_888), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_893), .A2(n_910), .B1(n_912), .B2(n_916), .C(n_919), .Y(n_909) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
AOI211xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_898), .B(n_900), .C(n_901), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
AND2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NOR3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_924), .C(n_941), .Y(n_908) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_921), .B(n_922), .Y(n_919) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI21xp33_ASAP7_75t_SL g924 ( .A1(n_925), .A2(n_927), .B(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_933), .B1(n_936), .B2(n_938), .Y(n_928) );
NOR2x1p5_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
BUFx3_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVxp67_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
BUFx6f_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx2_ASAP7_75t_SL g959 ( .A(n_960), .Y(n_959) );
endmodule