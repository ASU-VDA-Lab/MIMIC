module fake_jpeg_4932_n_29 (n_3, n_2, n_1, n_0, n_4, n_5, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_3),
.Y(n_6)
);

BUFx5_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

HB1xp67_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_0),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

OAI32xp33_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_18),
.B1(n_7),
.B2(n_9),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_1),
.B(n_2),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_17),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_4),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_5),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_15),
.B(n_14),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_9),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_20),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_11),
.C(n_12),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_20),
.C(n_21),
.Y(n_27)
);

OAI22x1_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_26),
.B1(n_8),
.B2(n_27),
.Y(n_29)
);


endmodule