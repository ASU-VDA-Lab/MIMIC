module fake_jpeg_7016_n_272 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_239;
wire n_72;
wire n_107;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_40),
.B(n_42),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_41),
.B(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_43),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_50),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_18),
.B1(n_36),
.B2(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_58),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_1),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_22),
.B(n_3),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_79),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_17),
.B(n_19),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_8),
.B(n_9),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_18),
.B1(n_39),
.B2(n_23),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_75),
.B(n_11),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_82),
.B1(n_89),
.B2(n_16),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_37),
.C(n_32),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_20),
.C(n_8),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_37),
.B1(n_26),
.B2(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_90),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_40),
.A2(n_29),
.B1(n_38),
.B2(n_24),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_97),
.B1(n_68),
.B2(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_38),
.B1(n_24),
.B2(n_28),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_38),
.B1(n_28),
.B2(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_28),
.B1(n_20),
.B2(n_6),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_58),
.B1(n_64),
.B2(n_48),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_47),
.A2(n_20),
.B1(n_4),
.B2(n_7),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_109),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_112),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_8),
.B(n_10),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_116),
.C(n_118),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_10),
.C(n_11),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_10),
.C(n_11),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_85),
.B1(n_81),
.B2(n_96),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_15),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_126),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_15),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_16),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_134),
.Y(n_149)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_128),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_93),
.B1(n_69),
.B2(n_92),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_130),
.B1(n_116),
.B2(n_132),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_72),
.B(n_86),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_101),
.B1(n_105),
.B2(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_145),
.B(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_155),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_80),
.Y(n_148)
);

OAI21x1_ASAP7_75t_SL g192 ( 
.A1(n_148),
.A2(n_139),
.B(n_143),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_90),
.B1(n_71),
.B2(n_70),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_157),
.B1(n_161),
.B2(n_106),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_98),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_162),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_127),
.B(n_78),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_96),
.B1(n_79),
.B2(n_71),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_117),
.B1(n_126),
.B2(n_129),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_70),
.B1(n_83),
.B2(n_78),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_160),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_95),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_109),
.B(n_110),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_113),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_171),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_175),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_179),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_180),
.B(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_182),
.Y(n_210)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_194),
.C(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_118),
.Y(n_186)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_108),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_142),
.B(n_112),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_191),
.B(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_112),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_166),
.B(n_149),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_141),
.B1(n_143),
.B2(n_156),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_206),
.B1(n_214),
.B2(n_186),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_207),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_188),
.B1(n_194),
.B2(n_174),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_169),
.B1(n_171),
.B2(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_161),
.B1(n_140),
.B2(n_154),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_157),
.B(n_147),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_140),
.B(n_154),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_154),
.B(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_170),
.Y(n_219)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_145),
.C(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_165),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_185),
.B(n_173),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_217),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_190),
.C(n_189),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_220),
.C(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_167),
.C(n_158),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_183),
.B1(n_176),
.B2(n_184),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_225),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_226),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_167),
.C(n_183),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_172),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_181),
.C(n_178),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_230),
.C(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_172),
.A3(n_146),
.B1(n_155),
.B2(n_159),
.C1(n_165),
.C2(n_144),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_223),
.B(n_201),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_205),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_212),
.B1(n_197),
.B2(n_203),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_221),
.B1(n_215),
.B2(n_214),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.C(n_224),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_212),
.B1(n_195),
.B2(n_205),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_204),
.B(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_247),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_250),
.B(n_207),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_246),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_248),
.B(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_217),
.B1(n_233),
.B2(n_238),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_238),
.B1(n_229),
.B2(n_231),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_255),
.C(n_239),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_245),
.A3(n_250),
.B1(n_231),
.B2(n_247),
.C1(n_220),
.C2(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_262),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_258),
.B(n_261),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_128),
.C(n_123),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_123),
.C(n_107),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_265),
.B(n_267),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_252),
.B1(n_256),
.B2(n_123),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_266),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_268),
.B(n_107),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_121),
.Y(n_272)
);


endmodule