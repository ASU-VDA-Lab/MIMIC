module fake_jpeg_1719_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_SL g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_48),
.B1(n_47),
.B2(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_77),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_57),
.B1(n_45),
.B2(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_49),
.B1(n_50),
.B2(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_61),
.B1(n_47),
.B2(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_57),
.B1(n_69),
.B2(n_64),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_90),
.B1(n_97),
.B2(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_69),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_44),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_74),
.B1(n_50),
.B2(n_44),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_105),
.B1(n_8),
.B2(n_9),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_50),
.B1(n_44),
.B2(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_114),
.B1(n_5),
.B2(n_7),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_1),
.B(n_2),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_10),
.B(n_12),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_20),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_23),
.C(n_40),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_111),
.C(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_4),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_95),
.B(n_7),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_16),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_129),
.B1(n_24),
.B2(n_26),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_8),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_100),
.B(n_109),
.C(n_104),
.D(n_103),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_131),
.B(n_36),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_29),
.C(n_39),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_134),
.C(n_22),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_14),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_27),
.C(n_38),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_15),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_32),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_42),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_17),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_18),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_152),
.C(n_134),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_151),
.B(n_153),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_150),
.B(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_34),
.C(n_35),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_152),
.C(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_124),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_153),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_139),
.B1(n_142),
.B2(n_145),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_169),
.B(n_163),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_167),
.B(n_159),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_157),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_146),
.Y(n_177)
);


endmodule