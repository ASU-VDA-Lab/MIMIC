module fake_netlist_6_60_n_1828 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1828);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1828;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_84),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_49),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_150),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_114),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_31),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_59),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_63),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_42),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_30),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_44),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_93),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_148),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_57),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_79),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_102),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_133),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_71),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_47),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_94),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_113),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_123),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_31),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_144),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_80),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_82),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_30),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_12),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_115),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_141),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_3),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_77),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_55),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_96),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_152),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_35),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_23),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_154),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_34),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_165),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_101),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_76),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_147),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_21),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_118),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_15),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_126),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_15),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_109),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_170),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_128),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_121),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_51),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_140),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_52),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_39),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_95),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_43),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_52),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_85),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_108),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_70),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_180),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_72),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_63),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_125),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_10),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_32),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_56),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_181),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_8),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_10),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_122),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_4),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_103),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_183),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_53),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_25),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_11),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_25),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_41),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_104),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_81),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_42),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_62),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_3),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_143),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_14),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_45),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_74),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_159),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_117),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_99),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_158),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_169),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_22),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_129),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_2),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_33),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_164),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_75),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_78),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_66),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_40),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_139),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_135),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_33),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_69),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_12),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_21),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_46),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_89),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_137),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_151),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_179),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_156),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_6),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_111),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_43),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_0),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_132),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_26),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_47),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_14),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_145),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_58),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_178),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_39),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_32),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_105),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_119),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_65),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_168),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_266),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_266),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_240),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_184),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_266),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_266),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_307),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_187),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_282),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_266),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_239),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_193),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_239),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_200),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_294),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_188),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_190),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_196),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_307),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_197),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_294),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_202),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_289),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_326),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_207),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_359),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_211),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_240),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_189),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_210),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_206),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_199),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_300),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_212),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_206),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_217),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_218),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_199),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_201),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_201),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_203),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_220),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_203),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_230),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_250),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_230),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_226),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_191),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_243),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_243),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_231),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_233),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_258),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_234),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_258),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_264),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_264),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_270),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_210),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_235),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_283),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_271),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_283),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_185),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_270),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_277),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_238),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_277),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_244),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_245),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_246),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_286),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_252),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_286),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_291),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_210),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_291),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_215),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_297),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_254),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_259),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_185),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_297),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_195),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_298),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_298),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_261),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_271),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_371),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_375),
.B(n_219),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_383),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_369),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_369),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_384),
.B(n_219),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_373),
.Y(n_481)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_379),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_422),
.B(n_315),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_373),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_377),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_376),
.A2(n_251),
.B1(n_311),
.B2(n_255),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_387),
.B(n_315),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_457),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_404),
.B(n_237),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_391),
.Y(n_495)
);

AND2x2_ASAP7_75t_SL g496 ( 
.A(n_397),
.B(n_186),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_378),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_411),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_380),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_396),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_439),
.B(n_323),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_412),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_398),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_381),
.A2(n_232),
.B1(n_299),
.B2(n_303),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_416),
.B(n_271),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_407),
.B(n_409),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_380),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_415),
.B(n_421),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_425),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_392),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_406),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_426),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_400),
.A2(n_302),
.B1(n_366),
.B2(n_301),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_388),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_370),
.A2(n_321),
.B1(n_253),
.B2(n_242),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_416),
.B(n_284),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_428),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_419),
.A2(n_299),
.B1(n_303),
.B2(n_312),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_437),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_389),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_389),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_410),
.Y(n_539)
);

OA21x2_ASAP7_75t_L g540 ( 
.A1(n_390),
.A2(n_198),
.B(n_194),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_374),
.B(n_323),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_386),
.B(n_358),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

AO21x2_ASAP7_75t_L g544 ( 
.A1(n_470),
.A2(n_198),
.B(n_194),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_467),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_490),
.B(n_541),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_493),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_493),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_479),
.B(n_435),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_541),
.B(n_442),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_445),
.Y(n_552)
);

AND3x2_ASAP7_75t_L g553 ( 
.A(n_484),
.B(n_337),
.C(n_186),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_446),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_481),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_448),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_533),
.B(n_397),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_468),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_511),
.B(n_358),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_474),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_208),
.C(n_205),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_529),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_503),
.A2(n_256),
.B1(n_237),
.B2(n_408),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_481),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_481),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_475),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_503),
.B(n_455),
.Y(n_571)
);

AOI21x1_ASAP7_75t_L g572 ( 
.A1(n_475),
.A2(n_208),
.B(n_205),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_216),
.C(n_214),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_494),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_504),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_494),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_494),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_523),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_503),
.B(n_542),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_476),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_496),
.B(n_419),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_456),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_467),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_542),
.A2(n_256),
.B1(n_438),
.B2(n_436),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_523),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_523),
.Y(n_589)
);

INVx6_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_216),
.C(n_214),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_523),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_496),
.A2(n_335),
.B1(n_312),
.B2(n_355),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_531),
.A2(n_213),
.B1(n_305),
.B2(n_306),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_477),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_477),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_526),
.A2(n_463),
.B1(n_405),
.B2(n_430),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_496),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_486),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_508),
.A2(n_463),
.B1(n_434),
.B2(n_437),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_485),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_540),
.A2(n_335),
.B1(n_355),
.B2(n_328),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_523),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_523),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_513),
.B(n_429),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_531),
.A2(n_330),
.B1(n_328),
.B2(n_316),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_539),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_535),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_486),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_488),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_535),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_486),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_499),
.Y(n_615)
);

INVx8_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_489),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_469),
.B(n_395),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_486),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_495),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_499),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_469),
.B(n_192),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_506),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_483),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_489),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_489),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_508),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_487),
.B(n_444),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_535),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_464),
.B(n_480),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_500),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_535),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_505),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_505),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_489),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_519),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_480),
.B(n_462),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_510),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_469),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_492),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_510),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_486),
.Y(n_647)
);

AO22x2_ASAP7_75t_L g648 ( 
.A1(n_509),
.A2(n_330),
.B1(n_222),
.B2(n_280),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_520),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_486),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_464),
.B(n_403),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_516),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_502),
.B(n_215),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_517),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_517),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_524),
.A2(n_222),
.B1(n_296),
.B2(n_324),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_537),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_469),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_514),
.B(n_284),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_489),
.B(n_227),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_521),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_526),
.A2(n_317),
.B1(n_336),
.B2(n_285),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_464),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_518),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_522),
.Y(n_669)
);

AO22x2_ASAP7_75t_L g670 ( 
.A1(n_527),
.A2(n_280),
.B1(n_224),
.B2(n_228),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_522),
.B(n_224),
.C(n_221),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_464),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_528),
.B(n_530),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_530),
.B(n_221),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_534),
.Y(n_677)
);

BUFx6f_ASAP7_75t_SL g678 ( 
.A(n_480),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_537),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_534),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_536),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_536),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_466),
.B(n_260),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_466),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_466),
.B(n_274),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_538),
.B(n_229),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_497),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_471),
.B(n_308),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_497),
.B(n_390),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_497),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_480),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_498),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_498),
.B(n_451),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_546),
.B(n_471),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_636),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_617),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_580),
.B(n_548),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_556),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_548),
.B(n_471),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_550),
.B(n_487),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_549),
.B(n_498),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_617),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_673),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_636),
.Y(n_705)
);

INVx8_ASAP7_75t_L g706 ( 
.A(n_616),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_598),
.A2(n_337),
.B1(n_367),
.B2(n_361),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_549),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_571),
.B(n_332),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_598),
.B(n_501),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_658),
.A2(n_585),
.B(n_551),
.C(n_554),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_552),
.B(n_215),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_584),
.A2(n_287),
.B1(n_263),
.B2(n_365),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_640),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_617),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_640),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_681),
.B(n_615),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_673),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_692),
.B(n_215),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_681),
.B(n_473),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_694),
.B(n_420),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_692),
.B(n_597),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_658),
.B(n_215),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_645),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_645),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_681),
.B(n_473),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_615),
.B(n_473),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_627),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_621),
.B(n_478),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_627),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_593),
.A2(n_361),
.B1(n_367),
.B2(n_364),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_690),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_690),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_621),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_676),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_628),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_606),
.B(n_204),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_R g738 ( 
.A(n_664),
.B(n_267),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_628),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_634),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_634),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_672),
.B(n_272),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_575),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_637),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_637),
.B(n_478),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_575),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_638),
.B(n_478),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_607),
.A2(n_318),
.B(n_313),
.C(n_249),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_576),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_638),
.B(n_247),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_624),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_643),
.B(n_247),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_662),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_643),
.B(n_248),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_676),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_577),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_599),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_603),
.A2(n_288),
.B1(n_364),
.B2(n_257),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_646),
.B(n_248),
.Y(n_759)
);

INVxp33_ASAP7_75t_L g760 ( 
.A(n_558),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_646),
.B(n_257),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_565),
.B(n_423),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_650),
.B(n_269),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_650),
.A2(n_288),
.B(n_273),
.C(n_278),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_653),
.B(n_656),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_631),
.A2(n_340),
.B1(n_295),
.B2(n_292),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_661),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_672),
.B(n_241),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_653),
.B(n_269),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_660),
.B(n_668),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_656),
.B(n_273),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_657),
.B(n_278),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_657),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_659),
.B(n_296),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_659),
.B(n_324),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_577),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_676),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_667),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_544),
.A2(n_341),
.B1(n_325),
.B2(n_327),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_667),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_562),
.A2(n_334),
.B1(n_275),
.B2(n_276),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_676),
.B(n_325),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_669),
.B(n_501),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_669),
.B(n_327),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_652),
.B(n_209),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_675),
.B(n_329),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_660),
.B(n_241),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_668),
.B(n_241),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_578),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_675),
.B(n_329),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_677),
.B(n_341),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_633),
.B(n_223),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_677),
.B(n_348),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_666),
.B(n_664),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_680),
.B(n_348),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_674),
.B(n_241),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_680),
.B(n_682),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_682),
.A2(n_427),
.B(n_431),
.C(n_432),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_627),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_689),
.B(n_491),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_689),
.B(n_543),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_578),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_674),
.B(n_241),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_544),
.A2(n_333),
.B1(n_284),
.B2(n_515),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_543),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_557),
.B(n_491),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_557),
.B(n_491),
.Y(n_807)
);

INVxp33_ASAP7_75t_L g808 ( 
.A(n_631),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_641),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_559),
.B(n_491),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_649),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_639),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_642),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_559),
.B(n_501),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_562),
.A2(n_345),
.B1(n_293),
.B2(n_304),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_686),
.B(n_512),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_560),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_661),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_562),
.B(n_225),
.Y(n_819)
);

AOI221xp5_ASAP7_75t_L g820 ( 
.A1(n_630),
.A2(n_262),
.B1(n_236),
.B2(n_265),
.C(n_268),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_560),
.B(n_512),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_561),
.B(n_512),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_679),
.B(n_333),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_561),
.B(n_515),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_679),
.B(n_333),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_562),
.B(n_279),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_671),
.A2(n_443),
.B(n_423),
.C(n_424),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_661),
.B(n_564),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_686),
.B(n_515),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_599),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_687),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_687),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_563),
.B(n_525),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_563),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_587),
.B(n_362),
.C(n_309),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_671),
.A2(n_686),
.B(n_573),
.C(n_591),
.Y(n_836)
);

INVx8_ASAP7_75t_L g837 ( 
.A(n_616),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_570),
.B(n_581),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_544),
.A2(n_333),
.B1(n_532),
.B2(n_525),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_564),
.B(n_333),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_686),
.B(n_525),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_562),
.A2(n_339),
.B1(n_290),
.B2(n_314),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_570),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_670),
.A2(n_532),
.B1(n_281),
.B2(n_363),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_581),
.B(n_532),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_583),
.B(n_319),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_566),
.B(n_424),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_666),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_573),
.B(n_322),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_639),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_663),
.B(n_310),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_583),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_665),
.B(n_331),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_691),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_595),
.A2(n_461),
.B(n_460),
.C(n_458),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_595),
.B(n_346),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_596),
.B(n_347),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_670),
.A2(n_354),
.B1(n_351),
.B2(n_349),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_596),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_591),
.B(n_623),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_601),
.B(n_482),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_601),
.B(n_602),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_648),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_SL g865 ( 
.A1(n_828),
.A2(n_618),
.B(n_644),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_816),
.Y(n_866)
);

BUFx8_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_698),
.B(n_602),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_749),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_701),
.A2(n_670),
.B1(n_648),
.B2(n_594),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_728),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_737),
.A2(n_678),
.B1(n_670),
.B2(n_648),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_711),
.B(n_620),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_853),
.A2(n_648),
.B1(n_616),
.B2(n_678),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_695),
.A2(n_626),
.B(n_684),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_610),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_702),
.B(n_610),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_703),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_721),
.B(n_813),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_816),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_829),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_735),
.B(n_620),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_735),
.B(n_620),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_709),
.A2(n_755),
.B1(n_777),
.B2(n_722),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_703),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_702),
.B(n_612),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_841),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_706),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_710),
.B(n_612),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_841),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_797),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_SL g893 ( 
.A1(n_808),
.A2(n_600),
.B1(n_625),
.B2(n_649),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_755),
.A2(n_678),
.B1(n_688),
.B2(n_685),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_710),
.B(n_683),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_731),
.A2(n_594),
.B1(n_693),
.B2(n_665),
.Y(n_896)
);

NOR2x2_ASAP7_75t_L g897 ( 
.A(n_766),
.B(n_641),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_797),
.B(n_654),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_704),
.B(n_639),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_696),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_708),
.B(n_626),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_848),
.B(n_616),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_732),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_718),
.B(n_655),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_708),
.B(n_582),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_777),
.A2(n_655),
.B1(n_616),
.B2(n_620),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_732),
.B(n_582),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_733),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_864),
.A2(n_693),
.B1(n_569),
.B2(n_568),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_733),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_734),
.B(n_553),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_847),
.B(n_608),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_783),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_758),
.A2(n_555),
.B1(n_568),
.B2(n_569),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_706),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_809),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_SL g917 ( 
.A(n_792),
.B(n_344),
.C(n_350),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_736),
.B(n_739),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_767),
.B(n_579),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_738),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_783),
.Y(n_921)
);

BUFx8_ASAP7_75t_L g922 ( 
.A(n_847),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_722),
.A2(n_605),
.B1(n_592),
.B2(n_635),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_760),
.B(n_545),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_751),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_760),
.B(n_427),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_779),
.A2(n_555),
.B1(n_338),
.B2(n_360),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_740),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_696),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_SL g930 ( 
.A1(n_808),
.A2(n_352),
.B1(n_353),
.B2(n_357),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_706),
.B(n_431),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_741),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_705),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_744),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_773),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_723),
.A2(n_356),
.B1(n_443),
.B2(n_458),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_811),
.B(n_432),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_782),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_851),
.A2(n_579),
.B1(n_588),
.B2(n_635),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_778),
.B(n_582),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_780),
.B(n_582),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_728),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_848),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_717),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_706),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_767),
.B(n_588),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_714),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_794),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_861),
.A2(n_647),
.B(n_589),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_753),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_805),
.B(n_586),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_817),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_728),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_834),
.B(n_433),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_837),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_785),
.B(n_433),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_843),
.B(n_586),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_837),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_715),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_715),
.B(n_611),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_SL g961 ( 
.A1(n_723),
.A2(n_613),
.B(n_609),
.C(n_605),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_852),
.B(n_586),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_837),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_782),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_846),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_742),
.B(n_572),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_860),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_714),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_767),
.B(n_589),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_765),
.B(n_586),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_801),
.B(n_545),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_700),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_818),
.B(n_592),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_730),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_818),
.B(n_604),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_820),
.B(n_440),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_716),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_818),
.B(n_604),
.Y(n_978)
);

AO22x1_ASAP7_75t_L g979 ( 
.A1(n_819),
.A2(n_449),
.B1(n_447),
.B2(n_441),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_838),
.B(n_609),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_730),
.B(n_440),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_727),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_863),
.B(n_836),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_712),
.A2(n_613),
.B1(n_632),
.B2(n_629),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_856),
.B(n_545),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_713),
.B(n_572),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_840),
.A2(n_441),
.B1(n_460),
.B2(n_454),
.Y(n_987)
);

OAI22xp33_ASAP7_75t_L g988 ( 
.A1(n_750),
.A2(n_461),
.B1(n_454),
.B2(n_452),
.Y(n_988)
);

BUFx2_ASAP7_75t_SL g989 ( 
.A(n_812),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_752),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_452),
.C(n_450),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_857),
.B(n_547),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_754),
.B(n_759),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_728),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_812),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_836),
.B(n_622),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_729),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_850),
.B(n_697),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_761),
.B(n_547),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_850),
.B(n_447),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_712),
.A2(n_719),
.B1(n_849),
.B2(n_861),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_763),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_769),
.B(n_771),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_697),
.B(n_449),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_799),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_716),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_697),
.B(n_450),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_745),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_724),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_799),
.B(n_647),
.Y(n_1010)
);

INVx6_ASAP7_75t_L g1011 ( 
.A(n_799),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_747),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_772),
.B(n_547),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_840),
.A2(n_622),
.B1(n_632),
.B2(n_629),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_799),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_774),
.B(n_567),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_831),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_775),
.B(n_567),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_707),
.A2(n_402),
.B1(n_399),
.B2(n_393),
.Y(n_1019)
);

AND2x6_ASAP7_75t_L g1020 ( 
.A(n_831),
.B(n_567),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_835),
.B(n_402),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_804),
.A2(n_393),
.B1(n_399),
.B2(n_574),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_784),
.B(n_786),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_790),
.B(n_574),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_724),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_770),
.A2(n_574),
.B(n_611),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_814),
.B(n_651),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_791),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_793),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_832),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_795),
.B(n_611),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_828),
.A2(n_611),
.B(n_614),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_844),
.B(n_0),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_757),
.B(n_651),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_821),
.B(n_651),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_832),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_798),
.B(n_651),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_748),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_822),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_719),
.B(n_614),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_854),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_824),
.B(n_651),
.Y(n_1042)
);

OR2x2_ASAP7_75t_SL g1043 ( 
.A(n_748),
.B(n_1),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_833),
.B(n_845),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_854),
.B(n_614),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_858),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_858),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_725),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_725),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_849),
.A2(n_614),
.B1(n_599),
.B2(n_482),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_781),
.B(n_599),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_855),
.A2(n_614),
.B(n_599),
.C(n_9),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_768),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_815),
.B(n_153),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_942),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_879),
.B(n_842),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_SL g1058 ( 
.A(n_893),
.B(n_859),
.C(n_827),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_983),
.A2(n_726),
.B(n_720),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_983),
.A2(n_830),
.B(n_770),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_904),
.B(n_965),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_917),
.A2(n_768),
.B(n_827),
.C(n_764),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1047),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_956),
.B(n_944),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_917),
.A2(n_876),
.B(n_1002),
.C(n_1033),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_944),
.B(n_743),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1054),
.A2(n_800),
.B1(n_806),
.B2(n_807),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1054),
.A2(n_810),
.B1(n_746),
.B2(n_756),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_885),
.A2(n_839),
.B1(n_789),
.B2(n_746),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_870),
.B(n_925),
.C(n_976),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_916),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_912),
.B(n_743),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1031),
.A2(n_862),
.B(n_756),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_869),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_993),
.A2(n_776),
.B(n_789),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_904),
.B(n_776),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_871),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_889),
.B(n_802),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1003),
.A2(n_802),
.B(n_619),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1028),
.B(n_825),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_900),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_SL g1082 ( 
.A(n_920),
.B(n_825),
.C(n_823),
.Y(n_1082)
);

OAI22x1_ASAP7_75t_L g1083 ( 
.A1(n_872),
.A2(n_823),
.B1(n_803),
.B2(n_796),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_929),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_933),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_950),
.B(n_788),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1002),
.B(n_787),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_892),
.B(n_787),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_870),
.A2(n_590),
.B1(n_619),
.B2(n_482),
.Y(n_1089)
);

OR2x6_ASAP7_75t_SL g1090 ( 
.A(n_948),
.B(n_5),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1023),
.A2(n_619),
.B(n_482),
.Y(n_1091)
);

NAND2x2_ASAP7_75t_L g1092 ( 
.A(n_943),
.B(n_7),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_871),
.Y(n_1093)
);

INVx11_ASAP7_75t_L g1094 ( 
.A(n_922),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_928),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_889),
.B(n_958),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_926),
.B(n_7),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_867),
.Y(n_1098)
);

NAND2x1_ASAP7_75t_L g1099 ( 
.A(n_915),
.B(n_590),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_990),
.B(n_9),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1001),
.A2(n_619),
.B(n_482),
.C(n_18),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_868),
.B(n_11),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_932),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_937),
.B(n_16),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_895),
.A2(n_482),
.B(n_619),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_913),
.A2(n_590),
.B1(n_619),
.B2(n_177),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_873),
.A2(n_590),
.B1(n_175),
.B2(n_173),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_896),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1029),
.B(n_19),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_972),
.B(n_20),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_934),
.B(n_22),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_981),
.B(n_23),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_898),
.A2(n_163),
.B(n_162),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_866),
.B(n_24),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_921),
.A2(n_160),
.B1(n_157),
.B2(n_131),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_985),
.A2(n_98),
.B(n_86),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_947),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_880),
.B(n_24),
.Y(n_1118)
);

INVx6_ASAP7_75t_L g1119 ( 
.A(n_922),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_896),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_992),
.A2(n_83),
.B(n_73),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1038),
.A2(n_882),
.B1(n_891),
.B2(n_888),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_996),
.A2(n_67),
.B(n_130),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_SL g1124 ( 
.A1(n_1040),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_881),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_968),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_996),
.A2(n_36),
.B(n_37),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_877),
.B(n_36),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_887),
.A2(n_38),
.B1(n_41),
.B2(n_44),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_1040),
.A2(n_38),
.B(n_48),
.C(n_49),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_977),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_988),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.C(n_55),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_935),
.B(n_50),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_890),
.B(n_58),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_952),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1021),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1044),
.A2(n_60),
.B(n_61),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_867),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_982),
.B(n_60),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1044),
.A2(n_61),
.B(n_62),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_865),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_997),
.B(n_1008),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_918),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_902),
.B(n_938),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_874),
.A2(n_908),
.B1(n_910),
.B2(n_903),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1012),
.B(n_1039),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_964),
.A2(n_874),
.B1(n_936),
.B2(n_1039),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_909),
.A2(n_1053),
.B1(n_989),
.B2(n_995),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1006),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_954),
.B(n_924),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1009),
.Y(n_1151)
);

NOR3xp33_ASAP7_75t_SL g1152 ( 
.A(n_930),
.B(n_991),
.C(n_884),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_954),
.B(n_924),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1025),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_981),
.B(n_1000),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_875),
.A2(n_970),
.B(n_971),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1017),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1032),
.A2(n_1018),
.B(n_1024),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_909),
.A2(n_995),
.B1(n_878),
.B2(n_959),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_902),
.B(n_906),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1000),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_999),
.A2(n_1016),
.B(n_1013),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_911),
.B(n_979),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_986),
.A2(n_936),
.B(n_873),
.C(n_894),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_974),
.B(n_911),
.Y(n_1165)
);

AO32x2_ASAP7_75t_L g1166 ( 
.A1(n_1036),
.A2(n_1005),
.A3(n_1015),
.B1(n_1052),
.B2(n_961),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1004),
.B(n_1007),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1004),
.B(n_1007),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_923),
.A2(n_980),
.B(n_907),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_998),
.B(n_899),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_871),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_883),
.A2(n_884),
.B1(n_899),
.B2(n_1051),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_R g1173 ( 
.A(n_878),
.B(n_886),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_L g1174 ( 
.A(n_974),
.B(n_883),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_901),
.B(n_959),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1027),
.A2(n_1035),
.B(n_1042),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_871),
.Y(n_1177)
);

OAI22x1_ASAP7_75t_L g1178 ( 
.A1(n_1051),
.A2(n_897),
.B1(n_1043),
.B2(n_886),
.Y(n_1178)
);

NOR3xp33_ASAP7_75t_L g1179 ( 
.A(n_988),
.B(n_1052),
.C(n_1019),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_980),
.A2(n_961),
.B(n_951),
.C(n_957),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_998),
.B(n_942),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1034),
.A2(n_945),
.B(n_955),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_953),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1030),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1048),
.B(n_1049),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1014),
.A2(n_975),
.B(n_978),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_905),
.B(n_1036),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_SL g1188 ( 
.A(n_919),
.B(n_978),
.C(n_969),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_919),
.A2(n_946),
.B(n_973),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_966),
.A2(n_927),
.B(n_962),
.C(n_941),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_953),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_946),
.A2(n_969),
.B(n_973),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_953),
.B(n_994),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_975),
.A2(n_1010),
.B(n_960),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1041),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_940),
.A2(n_1045),
.B(n_1050),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1046),
.B(n_1011),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_960),
.A2(n_1050),
.B1(n_1011),
.B2(n_963),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_987),
.B(n_927),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_L g1200 ( 
.A1(n_1045),
.A2(n_949),
.B(n_1010),
.C(n_1015),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1022),
.B(n_994),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1022),
.B(n_994),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_939),
.A2(n_1014),
.B(n_1037),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_914),
.A2(n_984),
.B(n_1026),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_953),
.B(n_994),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1005),
.B(n_915),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1011),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1019),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_963),
.Y(n_1209)
);

OAI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_931),
.A2(n_1037),
.B1(n_987),
.B2(n_914),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_931),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1037),
.A2(n_701),
.B(n_853),
.C(n_722),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1071),
.Y(n_1213)
);

OAI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1104),
.A2(n_1020),
.B(n_1064),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1098),
.Y(n_1215)
);

AOI221x1_ASAP7_75t_L g1216 ( 
.A1(n_1179),
.A2(n_1020),
.B1(n_1145),
.B2(n_1141),
.C(n_1164),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1212),
.B(n_1136),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1143),
.B(n_1142),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1065),
.A2(n_1210),
.B(n_1199),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1095),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1191),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1146),
.B(n_1072),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_SL g1223 ( 
.A1(n_1108),
.A2(n_1120),
.B(n_1101),
.C(n_1130),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_SL g1224 ( 
.A(n_1132),
.B(n_1152),
.C(n_1058),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1150),
.B(n_1153),
.Y(n_1225)
);

AO21x2_ASAP7_75t_L g1226 ( 
.A1(n_1204),
.A2(n_1156),
.B(n_1158),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1119),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1062),
.A2(n_1203),
.B(n_1102),
.C(n_1068),
.Y(n_1228)
);

NAND2x1_ASAP7_75t_L g1229 ( 
.A(n_1055),
.B(n_1171),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1103),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1208),
.B(n_1056),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1097),
.B(n_1066),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1135),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1119),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1162),
.A2(n_1158),
.B(n_1190),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1169),
.A2(n_1196),
.B(n_1059),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_SL g1237 ( 
.A1(n_1139),
.A2(n_1110),
.B(n_1134),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1127),
.A2(n_1172),
.B(n_1188),
.C(n_1123),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1155),
.B(n_1122),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1060),
.A2(n_1073),
.B(n_1075),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1159),
.A2(n_1079),
.A3(n_1187),
.B(n_1123),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_SL g1242 ( 
.A(n_1211),
.B(n_1055),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1109),
.A2(n_1086),
.B(n_1128),
.C(n_1107),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1061),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1180),
.A2(n_1194),
.B(n_1182),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1087),
.B(n_1076),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1200),
.A2(n_1186),
.B(n_1182),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1167),
.B(n_1168),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1198),
.A2(n_1067),
.B(n_1202),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1074),
.B(n_1170),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1105),
.A2(n_1099),
.B(n_1091),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1161),
.B(n_1165),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1105),
.A2(n_1185),
.B(n_1113),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1113),
.A2(n_1201),
.B(n_1121),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1119),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1080),
.A2(n_1077),
.B(n_1181),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1193),
.A2(n_1174),
.B(n_1175),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1147),
.B(n_1163),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1077),
.A2(n_1160),
.B(n_1148),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1100),
.B(n_1111),
.Y(n_1260)
);

NOR4xp25_ASAP7_75t_L g1261 ( 
.A(n_1132),
.B(n_1129),
.C(n_1125),
.D(n_1133),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1077),
.A2(n_1206),
.B(n_1205),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1137),
.A2(n_1140),
.A3(n_1106),
.B(n_1121),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1114),
.B(n_1118),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_1116),
.B(n_1112),
.C(n_1124),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1209),
.B(n_1211),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1096),
.A2(n_1093),
.B(n_1089),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1195),
.B(n_1178),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1144),
.A2(n_1082),
.B1(n_1197),
.B2(n_1138),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1207),
.B(n_1085),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1116),
.A2(n_1088),
.B(n_1184),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1078),
.A2(n_1157),
.B(n_1171),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1081),
.A2(n_1117),
.B(n_1154),
.C(n_1151),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1084),
.B(n_1126),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1131),
.B(n_1149),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1078),
.A2(n_1096),
.B(n_1063),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1057),
.B(n_1173),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1115),
.A2(n_1077),
.B(n_1183),
.C(n_1177),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1177),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1183),
.A2(n_1166),
.B(n_1092),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1090),
.B(n_1094),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1189),
.A2(n_949),
.B(n_1192),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1156),
.A2(n_1162),
.B(n_1158),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1164),
.A2(n_915),
.B(n_889),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1064),
.B(n_879),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1212),
.A2(n_701),
.B(n_853),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1212),
.B(n_699),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1204),
.A2(n_1164),
.B(n_1176),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1071),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1212),
.A2(n_701),
.B(n_853),
.Y(n_1290)
);

NOR4xp25_ASAP7_75t_L g1291 ( 
.A(n_1212),
.B(n_1120),
.C(n_1108),
.D(n_1132),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1083),
.A2(n_1164),
.A3(n_1145),
.B(n_1101),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1095),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1064),
.B(n_879),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1212),
.B(n_699),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_873),
.B(n_1204),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1142),
.B(n_1143),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1212),
.B(n_699),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1071),
.Y(n_1299)
);

OAI22x1_ASAP7_75t_L g1300 ( 
.A1(n_1070),
.A2(n_701),
.B1(n_872),
.B2(n_853),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1083),
.A2(n_1164),
.A3(n_1145),
.B(n_1101),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1072),
.B(n_608),
.Y(n_1302)
);

BUFx2_ASAP7_75t_R g1303 ( 
.A(n_1071),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1077),
.B(n_889),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1072),
.B(n_608),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1064),
.B(n_879),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_L g1307 ( 
.A(n_1212),
.B(n_737),
.C(n_701),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1095),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1095),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1072),
.B(n_608),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1095),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1072),
.B(n_608),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1164),
.A2(n_873),
.B(n_1204),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1071),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1064),
.B(n_879),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1064),
.B(n_879),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1071),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1212),
.A2(n_701),
.B(n_737),
.C(n_1065),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1064),
.B(n_879),
.Y(n_1319)
);

AOI211x1_ASAP7_75t_L g1320 ( 
.A1(n_1070),
.A2(n_722),
.B(n_1033),
.C(n_1127),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1064),
.B(n_879),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1064),
.B(n_879),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1212),
.B(n_699),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1083),
.A2(n_1164),
.A3(n_1145),
.B(n_1101),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1055),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1097),
.B(n_912),
.Y(n_1326)
);

AO32x2_ASAP7_75t_L g1327 ( 
.A1(n_1145),
.A2(n_864),
.A3(n_1129),
.B1(n_1069),
.B2(n_707),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1097),
.B(n_912),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1212),
.B(n_699),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1095),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1159),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1071),
.Y(n_1332)
);

AOI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1212),
.A2(n_737),
.B(n_701),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1056),
.A2(n_701),
.B1(n_853),
.B2(n_737),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1212),
.A2(n_701),
.B(n_737),
.C(n_1065),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1071),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1203),
.A2(n_1059),
.B(n_1162),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1141),
.A2(n_1164),
.B(n_1212),
.C(n_1120),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1195),
.Y(n_1339)
);

AOI31xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1132),
.A2(n_701),
.A3(n_853),
.B(n_699),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1064),
.B(n_879),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1095),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1070),
.A2(n_870),
.B1(n_1212),
.B2(n_1142),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1156),
.A2(n_1162),
.B(n_1158),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1072),
.B(n_608),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1212),
.A2(n_701),
.B(n_737),
.C(n_1065),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1071),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_1074),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1224),
.A2(n_1334),
.B1(n_1307),
.B2(n_1333),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1235),
.A2(n_1216),
.A3(n_1228),
.B(n_1344),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1260),
.A2(n_1218),
.B1(n_1297),
.B2(n_1231),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1297),
.B(n_1285),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1325),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1230),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1255),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1343),
.A2(n_1340),
.B1(n_1258),
.B2(n_1326),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1233),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1293),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1247),
.A2(n_1253),
.B(n_1240),
.Y(n_1359)
);

INVx6_ASAP7_75t_L g1360 ( 
.A(n_1221),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1308),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1248),
.B(n_1239),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1309),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1311),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1318),
.A2(n_1335),
.A3(n_1346),
.B(n_1238),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1328),
.B(n_1270),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1330),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1261),
.A2(n_1243),
.B(n_1264),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1280),
.A2(n_1257),
.B(n_1259),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1342),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1244),
.Y(n_1371)
);

AOI21xp33_ASAP7_75t_L g1372 ( 
.A1(n_1287),
.A2(n_1329),
.B(n_1295),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1217),
.B(n_1298),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1219),
.A2(n_1343),
.B(n_1337),
.C(n_1249),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1269),
.A2(n_1268),
.B1(n_1294),
.B2(n_1341),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1213),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_SL g1377 ( 
.A1(n_1256),
.A2(n_1271),
.B(n_1262),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1339),
.B(n_1266),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1219),
.A2(n_1271),
.B(n_1226),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1323),
.A2(n_1265),
.B1(n_1214),
.B2(n_1225),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1265),
.A2(n_1331),
.B(n_1278),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1246),
.A2(n_1232),
.B(n_1222),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1325),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1272),
.A2(n_1273),
.B(n_1276),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1237),
.A2(n_1288),
.B(n_1284),
.Y(n_1385)
);

AOI222xp33_ASAP7_75t_L g1386 ( 
.A1(n_1306),
.A2(n_1319),
.B1(n_1316),
.B2(n_1321),
.C1(n_1315),
.C2(n_1322),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1288),
.A2(n_1267),
.B(n_1304),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1325),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1338),
.A2(n_1236),
.B(n_1296),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1304),
.A2(n_1229),
.B(n_1275),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1347),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1215),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1279),
.A2(n_1277),
.B(n_1274),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1310),
.B(n_1345),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1250),
.A2(n_1252),
.B1(n_1312),
.B2(n_1313),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1320),
.B(n_1289),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1292),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1292),
.A2(n_1324),
.B(n_1301),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1325),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1340),
.A2(n_1291),
.B(n_1223),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1289),
.B(n_1261),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1291),
.A2(n_1242),
.B(n_1317),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1266),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1242),
.A2(n_1241),
.B(n_1324),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_SL g1406 ( 
.A(n_1299),
.B(n_1314),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1336),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1348),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_SL g1409 ( 
.A1(n_1327),
.A2(n_1263),
.B(n_1301),
.C(n_1324),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1332),
.A2(n_1281),
.B(n_1227),
.C(n_1234),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1241),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1348),
.A2(n_1290),
.B(n_1286),
.C(n_1340),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1334),
.A2(n_701),
.B1(n_1290),
.B2(n_1286),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1224),
.A2(n_701),
.B1(n_1334),
.B2(n_1307),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1336),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1220),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1220),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1218),
.B(n_1297),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1307),
.B(n_1212),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1220),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1220),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_SL g1422 ( 
.A(n_1303),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1286),
.A2(n_1212),
.B(n_1290),
.C(n_1334),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1224),
.A2(n_701),
.B1(n_1334),
.B2(n_1307),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1220),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1220),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1225),
.B(n_1300),
.Y(n_1427)
);

NAND2x1p5_ASAP7_75t_L g1428 ( 
.A(n_1325),
.B(n_1077),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1220),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1336),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1220),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1347),
.Y(n_1432)
);

BUFx12f_ASAP7_75t_L g1433 ( 
.A(n_1213),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1286),
.A2(n_1290),
.B(n_1340),
.C(n_1333),
.Y(n_1434)
);

INVx3_ASAP7_75t_SL g1435 ( 
.A(n_1213),
.Y(n_1435)
);

AND2x2_ASAP7_75t_SL g1436 ( 
.A(n_1291),
.B(n_1261),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1220),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1220),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1220),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1235),
.A2(n_1216),
.A3(n_1228),
.B(n_1283),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1286),
.A2(n_1290),
.B(n_1340),
.C(n_1333),
.Y(n_1441)
);

AO21x2_ASAP7_75t_L g1442 ( 
.A1(n_1240),
.A2(n_1235),
.B(n_1245),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1307),
.A2(n_1334),
.B(n_1333),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1240),
.A2(n_1235),
.B(n_1283),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1251),
.A2(n_1245),
.B(n_1282),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1334),
.B(n_701),
.C(n_737),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1235),
.A2(n_1216),
.A3(n_1228),
.B(n_1283),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1224),
.A2(n_701),
.B1(n_1334),
.B2(n_1307),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1251),
.A2(n_1245),
.B(n_1282),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1251),
.A2(n_1245),
.B(n_1282),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1218),
.B(n_1297),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1224),
.A2(n_701),
.B1(n_1334),
.B2(n_1307),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1220),
.Y(n_1455)
);

OAI21xp33_ASAP7_75t_L g1456 ( 
.A1(n_1334),
.A2(n_701),
.B(n_737),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1362),
.B(n_1386),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1362),
.B(n_1436),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1414),
.A2(n_1424),
.B1(n_1450),
.B2(n_1454),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1389),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1366),
.B(n_1427),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1456),
.A2(n_1448),
.B(n_1423),
.Y(n_1462)
);

INVxp67_ASAP7_75t_SL g1463 ( 
.A(n_1407),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1427),
.B(n_1356),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1402),
.B(n_1395),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1397),
.B(n_1375),
.Y(n_1466)
);

AOI21x1_ASAP7_75t_SL g1467 ( 
.A1(n_1418),
.A2(n_1453),
.B(n_1352),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1436),
.B(n_1368),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1423),
.A2(n_1443),
.B(n_1410),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1430),
.B(n_1389),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1351),
.B(n_1444),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1444),
.B(n_1446),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1442),
.A2(n_1445),
.B(n_1374),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1349),
.A2(n_1413),
.B1(n_1374),
.B2(n_1422),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1380),
.A2(n_1434),
.B1(n_1441),
.B2(n_1396),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1382),
.B(n_1373),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1419),
.A2(n_1412),
.B(n_1372),
.C(n_1373),
.Y(n_1477)
);

NOR2xp67_ASAP7_75t_L g1478 ( 
.A(n_1408),
.B(n_1415),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1428),
.A2(n_1353),
.B(n_1381),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1408),
.B(n_1433),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1354),
.A2(n_1361),
.B1(n_1439),
.B2(n_1438),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1401),
.A2(n_1403),
.B(n_1377),
.C(n_1369),
.Y(n_1482)
);

CKINVDCx8_ASAP7_75t_R g1483 ( 
.A(n_1376),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1390),
.A2(n_1405),
.B(n_1359),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1435),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1357),
.A2(n_1455),
.B1(n_1420),
.B2(n_1421),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1417),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1409),
.A2(n_1358),
.B(n_1367),
.C(n_1437),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1381),
.B(n_1365),
.Y(n_1489)
);

BUFx8_ASAP7_75t_L g1490 ( 
.A(n_1392),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1363),
.A2(n_1426),
.B1(n_1370),
.B2(n_1416),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1428),
.A2(n_1353),
.B(n_1381),
.Y(n_1492)
);

INVx3_ASAP7_75t_SL g1493 ( 
.A(n_1435),
.Y(n_1493)
);

AOI221x1_ASAP7_75t_SL g1494 ( 
.A1(n_1364),
.A2(n_1429),
.B1(n_1425),
.B2(n_1378),
.C(n_1431),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1371),
.B(n_1406),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1394),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1394),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1371),
.A2(n_1398),
.B1(n_1360),
.B2(n_1432),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1353),
.A2(n_1445),
.B(n_1404),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1387),
.B(n_1385),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1393),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1360),
.A2(n_1355),
.B1(n_1399),
.B2(n_1411),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1383),
.A2(n_1400),
.B1(n_1388),
.B2(n_1365),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1350),
.B(n_1449),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1350),
.A2(n_1449),
.B1(n_1440),
.B2(n_1384),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1393),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1350),
.A2(n_1449),
.B1(n_1440),
.B2(n_1384),
.Y(n_1507)
);

CKINVDCx6p67_ASAP7_75t_R g1508 ( 
.A(n_1391),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1440),
.B(n_1449),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1391),
.B(n_1379),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1452),
.B(n_1447),
.Y(n_1511)
);

AOI221x1_ASAP7_75t_SL g1512 ( 
.A1(n_1451),
.A2(n_701),
.B1(n_853),
.B2(n_1368),
.C(n_1456),
.Y(n_1512)
);

AND2x6_ASAP7_75t_L g1513 ( 
.A(n_1451),
.B(n_1353),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1456),
.A2(n_1212),
.B(n_1318),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1402),
.B(n_1395),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1366),
.B(n_1427),
.Y(n_1516)
);

A2O1A1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1456),
.A2(n_1290),
.B(n_1286),
.C(n_1448),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1456),
.A2(n_1448),
.B1(n_701),
.B2(n_1333),
.C(n_1334),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1362),
.B(n_1351),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1408),
.B(n_1302),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1390),
.A2(n_1405),
.B(n_1254),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1402),
.B(n_1395),
.Y(n_1522)
);

AOI221x1_ASAP7_75t_SL g1523 ( 
.A1(n_1368),
.A2(n_701),
.B1(n_853),
.B2(n_1456),
.C(n_1448),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1392),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1362),
.B(n_1386),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1355),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1456),
.A2(n_1212),
.B(n_1318),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1407),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1496),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1500),
.B(n_1510),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1509),
.B(n_1504),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1459),
.A2(n_1474),
.B1(n_1518),
.B2(n_1457),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1488),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1500),
.B(n_1513),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1500),
.B(n_1513),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1459),
.A2(n_1474),
.B1(n_1457),
.B2(n_1525),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1473),
.B(n_1499),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1526),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1470),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_L g1541 ( 
.A(n_1462),
.B(n_1517),
.C(n_1525),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1505),
.B(n_1507),
.Y(n_1542)
);

INVx3_ASAP7_75t_SL g1543 ( 
.A(n_1508),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1479),
.B(n_1492),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1458),
.B(n_1519),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1489),
.B(n_1521),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1521),
.B(n_1505),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1458),
.B(n_1466),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1513),
.Y(n_1549)
);

OR2x6_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1527),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1471),
.B(n_1487),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1502),
.B(n_1484),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1513),
.B(n_1511),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1461),
.B(n_1516),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1502),
.B(n_1468),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1471),
.A2(n_1476),
.B(n_1475),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1481),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1486),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1475),
.A2(n_1472),
.B1(n_1464),
.B2(n_1460),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1494),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1503),
.A2(n_1482),
.B(n_1469),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1491),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1528),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1465),
.B(n_1522),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1515),
.B(n_1463),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1498),
.B(n_1477),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1498),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1512),
.Y(n_1568)
);

NAND4xp25_ASAP7_75t_L g1569 ( 
.A(n_1533),
.B(n_1523),
.C(n_1520),
.D(n_1495),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1552),
.B(n_1524),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1529),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1529),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1530),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1549),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1530),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1533),
.A2(n_1483),
.B1(n_1478),
.B2(n_1506),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1556),
.B(n_1467),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1535),
.B(n_1480),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1560),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1532),
.B(n_1553),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1485),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1541),
.A2(n_1537),
.B1(n_1550),
.B2(n_1559),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1493),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1553),
.B(n_1506),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_SL g1588 ( 
.A(n_1561),
.B(n_1506),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1501),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1571),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1585),
.B(n_1541),
.C(n_1537),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1571),
.Y(n_1593)
);

AOI33xp33_ASAP7_75t_L g1594 ( 
.A1(n_1585),
.A2(n_1559),
.A3(n_1568),
.B1(n_1540),
.B2(n_1566),
.B3(n_1555),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1583),
.B(n_1573),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1572),
.Y(n_1596)
);

AOI211xp5_ASAP7_75t_L g1597 ( 
.A1(n_1569),
.A2(n_1566),
.B(n_1568),
.C(n_1534),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1571),
.Y(n_1598)
);

AO21x1_ASAP7_75t_SL g1599 ( 
.A1(n_1580),
.A2(n_1560),
.B(n_1552),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1585),
.A2(n_1550),
.B1(n_1566),
.B2(n_1534),
.C(n_1538),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1576),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1582),
.B(n_1540),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1584),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1579),
.A2(n_1550),
.B1(n_1567),
.B2(n_1545),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1574),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1570),
.B(n_1542),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1573),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1579),
.A2(n_1550),
.B1(n_1567),
.B2(n_1545),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1583),
.B(n_1531),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1583),
.B(n_1531),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1590),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1564),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1569),
.A2(n_1548),
.B1(n_1564),
.B2(n_1555),
.C(n_1563),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1542),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.B(n_1542),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1576),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1578),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_1531),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1579),
.A2(n_1550),
.B1(n_1556),
.B2(n_1561),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1589),
.B(n_1539),
.Y(n_1621)
);

OAI33xp33_ASAP7_75t_L g1622 ( 
.A1(n_1582),
.A2(n_1548),
.A3(n_1565),
.B1(n_1551),
.B2(n_1557),
.B3(n_1558),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1582),
.A2(n_1567),
.B1(n_1556),
.B2(n_1555),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1531),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1590),
.B(n_1536),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1575),
.B(n_1562),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1591),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1596),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1625),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1596),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1626),
.B(n_1575),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1613),
.B(n_1589),
.Y(n_1634)
);

INVx4_ASAP7_75t_SL g1635 ( 
.A(n_1612),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1612),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1593),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1601),
.Y(n_1638)
);

OR2x6_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1538),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1617),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1592),
.B(n_1556),
.C(n_1580),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1618),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1625),
.B(n_1538),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1592),
.B(n_1597),
.C(n_1614),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1605),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1611),
.Y(n_1648)
);

OR2x6_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1538),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1647),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1647),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1633),
.B(n_1626),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1643),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1629),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1634),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1646),
.B(n_1602),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1646),
.A2(n_1597),
.B(n_1594),
.C(n_1600),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1629),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1643),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1610),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1603),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1635),
.B(n_1610),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1633),
.B(n_1640),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1641),
.B(n_1556),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1641),
.B(n_1640),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1636),
.B(n_1589),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1638),
.B(n_1554),
.Y(n_1670)
);

BUFx12f_ASAP7_75t_L g1671 ( 
.A(n_1636),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1627),
.Y(n_1672)
);

NAND4xp25_ASAP7_75t_L g1673 ( 
.A(n_1644),
.B(n_1620),
.C(n_1604),
.D(n_1608),
.Y(n_1673)
);

NAND4xp25_ASAP7_75t_L g1674 ( 
.A(n_1644),
.B(n_1608),
.C(n_1604),
.D(n_1623),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1589),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1635),
.B(n_1595),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1627),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1624),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1628),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1628),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1636),
.B(n_1588),
.C(n_1623),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1632),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1632),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1635),
.B(n_1624),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_SL g1685 ( 
.A1(n_1636),
.A2(n_1539),
.B1(n_1544),
.B2(n_1581),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1637),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1637),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1638),
.B(n_1616),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1642),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1639),
.B(n_1611),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1639),
.A2(n_1561),
.B1(n_1621),
.B2(n_1588),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1672),
.Y(n_1692)
);

INVxp67_ASAP7_75t_SL g1693 ( 
.A(n_1668),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1586),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1663),
.B(n_1639),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1666),
.B(n_1586),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1671),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1657),
.A2(n_1674),
.B(n_1673),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1656),
.B(n_1622),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1658),
.B(n_1644),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1654),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_SL g1703 ( 
.A(n_1656),
.B(n_1577),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1654),
.B(n_1644),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_1606),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.B(n_1606),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1660),
.B(n_1670),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1662),
.B(n_1615),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1672),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1666),
.B(n_1586),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1660),
.B(n_1615),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1688),
.B(n_1616),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1677),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1671),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1677),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_1665),
.B(n_1580),
.C(n_1551),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1667),
.B(n_1586),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1667),
.B(n_1639),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1655),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1688),
.B(n_1607),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1669),
.B(n_1587),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1679),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1651),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1679),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1675),
.B(n_1587),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1680),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1676),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1711),
.B(n_1653),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1701),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1728),
.B(n_1678),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1728),
.B(n_1678),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1703),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1695),
.B(n_1684),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1694),
.Y(n_1736)
);

INVxp67_ASAP7_75t_L g1737 ( 
.A(n_1694),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1704),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1702),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1714),
.B(n_1684),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1719),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1692),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1709),
.Y(n_1743)
);

INVxp33_ASAP7_75t_L g1744 ( 
.A(n_1700),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1713),
.Y(n_1745)
);

NOR2x1_ASAP7_75t_L g1746 ( 
.A(n_1700),
.B(n_1652),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1696),
.B(n_1676),
.Y(n_1747)
);

CKINVDCx16_ASAP7_75t_R g1748 ( 
.A(n_1698),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1697),
.B(n_1650),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1693),
.A2(n_1691),
.B1(n_1681),
.B2(n_1685),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1707),
.B(n_1652),
.Y(n_1751)
);

NOR2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1693),
.B(n_1577),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1719),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1705),
.Y(n_1754)
);

XNOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1746),
.B(n_1750),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1744),
.A2(n_1699),
.B1(n_1718),
.B2(n_1696),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1730),
.A2(n_1716),
.B(n_1723),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_L g1758 ( 
.A(n_1730),
.B(n_1723),
.C(n_1722),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1747),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

AOI222xp33_ASAP7_75t_L g1761 ( 
.A1(n_1746),
.A2(n_1750),
.B1(n_1738),
.B2(n_1734),
.C1(n_1737),
.C2(n_1739),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1736),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1737),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1747),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1739),
.B(n_1696),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1739),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1738),
.B(n_1721),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1721),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1741),
.Y(n_1769)
);

NAND2x1_ASAP7_75t_SL g1770 ( 
.A(n_1747),
.B(n_1718),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1726),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1733),
.A2(n_1706),
.B1(n_1712),
.B2(n_1708),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1741),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1740),
.A2(n_1726),
.B1(n_1727),
.B2(n_1715),
.C(n_1725),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1767),
.B(n_1754),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1759),
.B(n_1754),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1764),
.B(n_1754),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_1768),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1765),
.B(n_1747),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1755),
.Y(n_1781)
);

OAI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1757),
.A2(n_1733),
.B1(n_1729),
.B2(n_1751),
.Y(n_1782)
);

NAND2x1_ASAP7_75t_SL g1783 ( 
.A(n_1760),
.B(n_1731),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1761),
.B(n_1749),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1756),
.A2(n_1732),
.B(n_1731),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1771),
.B(n_1751),
.Y(n_1786)
);

AO22x1_ASAP7_75t_L g1787 ( 
.A1(n_1781),
.A2(n_1762),
.B1(n_1766),
.B2(n_1763),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1784),
.A2(n_1785),
.B(n_1783),
.Y(n_1788)
);

OA22x2_ASAP7_75t_L g1789 ( 
.A1(n_1785),
.A2(n_1765),
.B1(n_1732),
.B2(n_1769),
.Y(n_1789)
);

NAND4xp25_ASAP7_75t_L g1790 ( 
.A(n_1786),
.B(n_1758),
.C(n_1774),
.D(n_1773),
.Y(n_1790)
);

AOI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1782),
.A2(n_1758),
.B(n_1772),
.C(n_1742),
.Y(n_1791)
);

OAI32xp33_ASAP7_75t_L g1792 ( 
.A1(n_1778),
.A2(n_1775),
.A3(n_1776),
.B1(n_1777),
.B2(n_1780),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1779),
.A2(n_1765),
.B(n_1743),
.Y(n_1793)
);

OAI222xp33_ASAP7_75t_L g1794 ( 
.A1(n_1781),
.A2(n_1729),
.B1(n_1735),
.B2(n_1749),
.C1(n_1742),
.C2(n_1745),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1784),
.B(n_1741),
.C(n_1753),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1781),
.A2(n_1752),
.B1(n_1735),
.B2(n_1718),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1787),
.B(n_1752),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_SL g1798 ( 
.A1(n_1793),
.A2(n_1753),
.B(n_1745),
.Y(n_1798)
);

O2A1O1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1788),
.A2(n_1743),
.B(n_1753),
.C(n_1720),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1791),
.A2(n_1717),
.B(n_1710),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1790),
.A2(n_1724),
.B1(n_1648),
.B2(n_1645),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1800),
.B(n_1796),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_SL g1803 ( 
.A(n_1798),
.B(n_1794),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1799),
.Y(n_1804)
);

NOR4xp75_ASAP7_75t_L g1805 ( 
.A(n_1797),
.B(n_1789),
.C(n_1792),
.D(n_1795),
.Y(n_1805)
);

NOR2xp67_ASAP7_75t_L g1806 ( 
.A(n_1801),
.B(n_1680),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1799),
.Y(n_1807)
);

OAI221xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1804),
.A2(n_1587),
.B1(n_1639),
.B2(n_1649),
.C(n_1645),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_1803),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1804),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1807),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_SL g1812 ( 
.A(n_1802),
.B(n_1599),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1809),
.B(n_1806),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1811),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_SL g1815 ( 
.A(n_1810),
.B(n_1805),
.C(n_1812),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1815),
.B(n_1812),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1814),
.B1(n_1813),
.B2(n_1808),
.C(n_1686),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1817),
.A2(n_1655),
.B1(n_1659),
.B2(n_1687),
.Y(n_1818)
);

XNOR2xp5_ASAP7_75t_L g1819 ( 
.A(n_1817),
.B(n_1490),
.Y(n_1819)
);

XNOR2xp5_ASAP7_75t_L g1820 ( 
.A(n_1819),
.B(n_1490),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1818),
.A2(n_1659),
.B1(n_1689),
.B2(n_1682),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1820),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1822),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1821),
.B(n_1683),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1683),
.B(n_1682),
.Y(n_1825)
);

AOI322xp5_ASAP7_75t_L g1826 ( 
.A1(n_1825),
.A2(n_1689),
.A3(n_1687),
.B1(n_1686),
.B2(n_1690),
.C1(n_1648),
.C2(n_1661),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1648),
.B1(n_1631),
.B2(n_1629),
.Y(n_1827)
);

AOI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1827),
.A2(n_1543),
.B(n_1690),
.C(n_1661),
.Y(n_1828)
);


endmodule