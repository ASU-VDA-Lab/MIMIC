module fake_jpeg_6112_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_1),
.Y(n_12)
);

INVx4_ASAP7_75t_SL g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_18),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_5),
.B1(n_14),
.B2(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_8),
.B1(n_12),
.B2(n_9),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_32),
.B1(n_25),
.B2(n_24),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_34),
.C(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_36),
.C(n_41),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_33),
.C(n_45),
.Y(n_48)
);


endmodule