module real_jpeg_31981_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_1),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_2),
.A2(n_14),
.B(n_470),
.Y(n_13)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_2),
.Y(n_472)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_61),
.B1(n_78),
.B2(n_83),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_3),
.B(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_R g138 ( 
.A(n_4),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_55),
.B1(n_138),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_4),
.A2(n_138),
.B1(n_256),
.B2(n_259),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_4),
.B(n_113),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_4),
.B(n_67),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_4),
.B(n_399),
.C(n_402),
.Y(n_398)
);

NAND2xp67_ASAP7_75t_L g414 ( 
.A(n_4),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_4),
.B(n_25),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_5),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_5),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_7),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_7),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_12),
.A2(n_105),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_12),
.A2(n_105),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_12),
.A2(n_105),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_178),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_177),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2x1_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_160),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_18),
.B(n_160),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_147),
.C(n_148),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_21),
.B(n_146),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_109),
.B2(n_146),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_65),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_24),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_24),
.A2(n_150),
.B1(n_159),
.B2(n_454),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_41),
.B(n_59),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_25),
.A2(n_237),
.B(n_245),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_25),
.A2(n_41),
.B1(n_59),
.B2(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_25),
.B(n_237),
.Y(n_280)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_27),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_27)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_28),
.Y(n_211)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_28),
.Y(n_234)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_30),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_30),
.Y(n_209)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_30),
.Y(n_220)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_34),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_36),
.Y(n_222)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g245 ( 
.A(n_42),
.B(n_246),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_43),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_52),
.B2(n_55),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_51),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_51),
.Y(n_359)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_58),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_61),
.A2(n_216),
.B(n_221),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_65),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_77),
.B1(n_87),
.B2(n_99),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_66),
.A2(n_77),
.B(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_88),
.B1(n_100),
.B2(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2x1p5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_89),
.Y(n_88)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_68),
.A2(n_88),
.B(n_151),
.Y(n_188)
);

OAI22x1_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_71),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_71),
.Y(n_368)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_81),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_104),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_150),
.C(n_158),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_110),
.B(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_110),
.A2(n_146),
.B1(n_226),
.B2(n_456),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2x1p5_ASAP7_75t_L g249 ( 
.A(n_111),
.B(n_250),
.Y(n_249)
);

AOI22x1_ASAP7_75t_L g281 ( 
.A1(n_111),
.A2(n_247),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_111),
.B(n_192),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

AO22x2_ASAP7_75t_L g187 ( 
.A1(n_112),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_124),
.B(n_137),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_116),
.Y(n_301)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

NAND2x1_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_135),
.Y(n_308)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_142),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_152),
.B(n_156),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_142),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_158),
.C(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_146),
.A2(n_147),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_149),
.B(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_150),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_155),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_156),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_175),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_168),
.B2(n_174),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_445),
.B(n_465),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_432),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_345),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_319),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_284),
.Y(n_182)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_183),
.Y(n_434)
);

NAND2x1p5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_267),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_184),
.B(n_267),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_225),
.C(n_248),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_186),
.B(n_225),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B1(n_223),
.B2(n_224),
.Y(n_186)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_187),
.B(n_253),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_187),
.A2(n_223),
.B1(n_292),
.B2(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_188),
.B(n_190),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_188),
.B(n_192),
.Y(n_329)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_190),
.Y(n_283)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_191),
.A2(n_249),
.B(n_264),
.Y(n_276)
);

NAND2x1p5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_192),
.B(n_254),
.Y(n_253)
);

XOR2x2_ASAP7_75t_SL g290 ( 
.A(n_192),
.B(n_197),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_192),
.A2(n_254),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_192),
.B(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_192),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_192),
.A2(n_293),
.B1(n_294),
.B2(n_325),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_192),
.A2(n_325),
.B1(n_393),
.B2(n_394),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_194),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_205),
.B1(n_212),
.B2(n_214),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_198),
.A2(n_205),
.B1(n_255),
.B2(n_260),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx4f_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2x1_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_235),
.B1(n_236),
.B2(n_247),
.Y(n_225)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OR2x6_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_255),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_233),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_252),
.B(n_264),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_266),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_272),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AND3x1_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_329),
.C(n_330),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_275),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_269),
.B(n_277),
.C(n_464),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_270),
.B(n_293),
.C(n_343),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_SL g348 ( 
.A1(n_270),
.A2(n_349),
.B(n_351),
.C(n_375),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_270),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_273),
.B(n_450),
.C(n_455),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_273),
.A2(n_274),
.B1(n_451),
.B2(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_276),
.Y(n_464)
);

XOR2x1_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_278),
.Y(n_456)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_284),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_285),
.B(n_287),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_290),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_296),
.Y(n_340)
);

NAND2x1p5_ASAP7_75t_L g379 ( 
.A(n_293),
.B(n_352),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_293),
.A2(n_294),
.B1(n_343),
.B2(n_344),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_293),
.B(n_380),
.C(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_293),
.B(n_422),
.Y(n_421)
);

CKINVDCx11_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_294),
.B(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_294),
.B(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_294),
.B(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_304),
.B(n_309),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx4f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_313),
.B(n_318),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_333),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_320),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_331),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_321),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.C(n_327),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_324),
.A2(n_327),
.B1(n_328),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_334),
.B(n_337),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.C(n_341),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_338),
.B(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_339),
.B(n_351),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_340),
.B(n_342),
.Y(n_430)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI21x1_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_427),
.B(n_431),
.Y(n_345)
);

AOI21x1_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_385),
.B(n_426),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_376),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_376),
.Y(n_426)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_350),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_350),
.B(n_379),
.C(n_381),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_356),
.B(n_364),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_369),
.B(n_373),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

OAI21x1_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_390),
.B(n_425),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_388),
.Y(n_425)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_391),
.A2(n_410),
.B(n_423),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_406),
.Y(n_391)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_392),
.Y(n_424)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_421),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_419),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_429),
.Y(n_431)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_436),
.B(n_442),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_443),
.B(n_444),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_459),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_467),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_457),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_457),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_451),
.Y(n_462)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_463),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);


endmodule