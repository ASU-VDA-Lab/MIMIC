module fake_jpeg_22316_n_80 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_1),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_3),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_56),
.B1(n_44),
.B2(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_62),
.C(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_57),
.Y(n_67)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_68),
.CI(n_57),
.CON(n_69),
.SN(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_63),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_70),
.CI(n_45),
.CON(n_72),
.SN(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_37),
.C(n_30),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_36),
.B(n_43),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_72),
.B(n_42),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_42),
.A3(n_38),
.B1(n_25),
.B2(n_70),
.C1(n_20),
.C2(n_23),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_9),
.B(n_38),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_60),
.B(n_58),
.Y(n_76)
);

OA21x2_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_28),
.B(n_39),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_55),
.C(n_48),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_78),
.C(n_4),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_28),
.Y(n_80)
);


endmodule