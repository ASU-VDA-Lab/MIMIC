module real_jpeg_28108_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_335, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_335;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_0),
.A2(n_31),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_0),
.A2(n_55),
.B1(n_64),
.B2(n_67),
.Y(n_119)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_1),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_2),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_130),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_64),
.B1(n_67),
.B2(n_130),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_130),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_135),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_135),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_3),
.A2(n_64),
.B1(n_67),
.B2(n_135),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_5),
.B(n_30),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_33),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_5),
.A2(n_33),
.B(n_175),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_133),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_5),
.A2(n_64),
.B(n_68),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_5),
.B(n_91),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_5),
.A2(n_112),
.B1(n_225),
.B2(n_226),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_7),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_128),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_128),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_7),
.A2(n_64),
.B1(n_67),
.B2(n_128),
.Y(n_217)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_9),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_9),
.A2(n_35),
.B1(n_64),
.B2(n_67),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_52),
.B1(n_64),
.B2(n_67),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_12),
.A2(n_37),
.B1(n_64),
.B2(n_67),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_12),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_258)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_15),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_98),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_96),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_77),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_20),
.A2(n_21),
.B1(n_73),
.B2(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_72),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_23),
.A2(n_38),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_23),
.A2(n_38),
.B1(n_141),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_23),
.A2(n_265),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_24),
.B(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_24),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_24),
.A2(n_30),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_24),
.A2(n_88),
.B(n_285),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_25),
.B(n_33),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_27),
.B(n_133),
.CON(n_132),
.SN(n_132)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_29),
.A2(n_31),
.B1(n_132),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_30),
.B(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_33),
.B1(n_46),
.B2(n_58),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_31),
.A2(n_47),
.A3(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_38),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_59),
.B2(n_71),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_59),
.C(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_43),
.A2(n_79),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_44),
.A2(n_56),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_44),
.A2(n_56),
.B1(n_127),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_44),
.A2(n_56),
.B1(n_158),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_44),
.A2(n_56),
.B1(n_81),
.B2(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_48),
.B(n_58),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_48),
.A2(n_62),
.B(n_133),
.C(n_203),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_53),
.A2(n_91),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_58),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_59),
.A2(n_71),
.B1(n_78),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_69),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_60),
.A2(n_69),
.B(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_60),
.A2(n_63),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_60),
.A2(n_183),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_60),
.A2(n_63),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_60),
.A2(n_63),
.B1(n_182),
.B2(n_201),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_60),
.A2(n_63),
.B1(n_107),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_60),
.A2(n_123),
.B(n_258),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_63),
.B(n_133),
.Y(n_223)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_67),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_70),
.B(n_124),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_73),
.C(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_73),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_73),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_77),
.B(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_78),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_82),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_79),
.A2(n_82),
.B(n_92),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI321xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_314),
.A3(n_326),
.B1(n_332),
.B2(n_333),
.C(n_335),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_296),
.B(n_313),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_271),
.B(n_295),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_164),
.B(n_249),
.C(n_270),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_150),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_103),
.B(n_150),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_136),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_120),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_105),
.B(n_120),
.C(n_136),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_106),
.B(n_111),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_108),
.B(n_193),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B(n_117),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_112),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_112),
.A2(n_217),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_112),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_113),
.A2(n_118),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_113),
.A2(n_114),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_114),
.B(n_172),
.Y(n_212)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_114),
.Y(n_290)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_149),
.B(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_131),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_133),
.B(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_138),
.B(n_143),
.C(n_145),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_151),
.A2(n_152),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_162),
.B(n_212),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_248),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_241),
.B(n_247),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_194),
.B(n_240),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_184),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_168),
.B(n_184),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.C(n_180),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_169),
.A2(n_170),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_173),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_172),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_191),
.C(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_234),
.B(n_239),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_213),
.B(n_233),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_221),
.B(n_232),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_219),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_231),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_250),
.B(n_251),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_268),
.B2(n_269),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_259),
.B2(n_260),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_260),
.C(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_263),
.C(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_273),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_294),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_286),
.B2(n_287),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_287),
.C(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_281),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_289),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_292),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_307),
.B(n_310),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_311),
.B2(n_312),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_306),
.C(n_312),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_316),
.C(n_322),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_316),
.B1(n_317),
.B2(n_331),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_305),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_323),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule