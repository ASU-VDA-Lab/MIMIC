module fake_jpeg_10949_n_84 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_24),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_30),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_32),
.B(n_33),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_54),
.B(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_34),
.Y(n_57)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_39),
.B(n_35),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_41),
.C(n_27),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_38),
.B(n_37),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_63),
.B1(n_40),
.B2(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_44),
.B1(n_40),
.B2(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_65),
.B1(n_46),
.B2(n_15),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_61),
.B1(n_65),
.B2(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_72),
.B1(n_2),
.B2(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_76),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_58),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_70),
.C(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_67),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_72),
.B1(n_66),
.B2(n_77),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_74),
.B(n_5),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_23),
.B(n_8),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_7),
.B1(n_12),
.B2(n_16),
.C(n_17),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_18),
.Y(n_84)
);


endmodule