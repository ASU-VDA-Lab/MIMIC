module fake_jpeg_28452_n_456 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_456);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_456;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_45),
.Y(n_142)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_68),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_87),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_16),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_16),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_90),
.Y(n_118)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_37),
.B(n_15),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_103),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_58),
.B(n_41),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_116),
.C(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_59),
.B(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_30),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_30),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_69),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_70),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_45),
.B(n_20),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_159),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_32),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_157),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_152),
.Y(n_204)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_107),
.A2(n_35),
.B1(n_55),
.B2(n_71),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_26),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_47),
.B1(n_53),
.B2(n_56),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_179),
.B1(n_186),
.B2(n_101),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_113),
.A2(n_79),
.B1(n_80),
.B2(n_65),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_182),
.B1(n_73),
.B2(n_96),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_26),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_35),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_35),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_171),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_135),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_99),
.B(n_33),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_62),
.B1(n_57),
.B2(n_32),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_183),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_99),
.A2(n_20),
.B1(n_86),
.B2(n_83),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_33),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_182),
.Y(n_200)
);

BUFx24_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_101),
.C(n_115),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_197),
.B1(n_208),
.B2(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_150),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_105),
.B1(n_95),
.B2(n_102),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_144),
.B1(n_95),
.B2(n_102),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_144),
.B1(n_105),
.B2(n_112),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_158),
.B1(n_175),
.B2(n_180),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_198),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_151),
.B1(n_157),
.B2(n_156),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_220),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_188),
.A2(n_158),
.B1(n_175),
.B2(n_183),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_168),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_160),
.B1(n_167),
.B2(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_223),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_153),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_238),
.B(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_148),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_194),
.B(n_192),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_184),
.B(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_227),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_230),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_205),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_236),
.Y(n_264)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_149),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_195),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_239),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_190),
.A2(n_206),
.B1(n_202),
.B2(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_198),
.A2(n_163),
.B(n_178),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_225),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_204),
.B(n_209),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_254),
.B(n_244),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_202),
.C(n_196),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_233),
.C(n_115),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_197),
.B1(n_208),
.B2(n_206),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_217),
.A2(n_209),
.B(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_262),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_214),
.B1(n_210),
.B2(n_180),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_193),
.B1(n_112),
.B2(n_174),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_193),
.B1(n_154),
.B2(n_147),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_229),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_221),
.B1(n_218),
.B2(n_222),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_232),
.B1(n_220),
.B2(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_275),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_278),
.B(n_284),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_274),
.A2(n_249),
.B1(n_254),
.B2(n_245),
.Y(n_312)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_166),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_281),
.C(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_239),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_285),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_237),
.B(n_186),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_243),
.A2(n_186),
.B(n_212),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_288),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_244),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_162),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_262),
.B(n_236),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_203),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_230),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_249),
.C(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_251),
.B1(n_256),
.B2(n_278),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_304),
.A2(n_309),
.B1(n_317),
.B2(n_242),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_250),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_251),
.B1(n_265),
.B2(n_259),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_265),
.B1(n_252),
.B2(n_247),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_310),
.A2(n_312),
.B1(n_321),
.B2(n_281),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_283),
.B(n_245),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_319),
.C(n_277),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_266),
.B1(n_267),
.B2(n_257),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_263),
.C(n_203),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_269),
.A2(n_270),
.B1(n_282),
.B2(n_275),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_285),
.A2(n_266),
.B(n_212),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_227),
.B(n_234),
.Y(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_297),
.A2(n_286),
.B(n_289),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_326),
.A2(n_338),
.B(n_340),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_311),
.A2(n_272),
.B1(n_234),
.B2(n_227),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_327),
.A2(n_336),
.B1(n_348),
.B2(n_313),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_332),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_231),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_337),
.C(n_343),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_324),
.B(n_11),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_335),
.B(n_344),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_165),
.C(n_173),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_186),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_342),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_312),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_211),
.C(n_131),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_310),
.A2(n_215),
.B1(n_176),
.B2(n_147),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_152),
.C(n_140),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_305),
.C(n_315),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_24),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_304),
.A2(n_176),
.B1(n_172),
.B2(n_104),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_298),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_359),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_298),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_355),
.A2(n_344),
.B1(n_348),
.B2(n_172),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_302),
.B1(n_323),
.B2(n_299),
.Y(n_356)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_367),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_307),
.Y(n_359)
);

AOI21xp33_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_307),
.B(n_300),
.Y(n_360)
);

OA21x2_ASAP7_75t_SL g374 ( 
.A1(n_360),
.A2(n_340),
.B(n_334),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_302),
.B1(n_323),
.B2(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_362),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_317),
.C(n_318),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_363),
.B(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_320),
.C(n_308),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_331),
.A2(n_315),
.B1(n_301),
.B2(n_309),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_322),
.C(n_301),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_187),
.C(n_140),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_370),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_128),
.Y(n_370)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_374),
.A2(n_386),
.B1(n_391),
.B2(n_369),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_352),
.A2(n_329),
.B(n_346),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_376),
.A2(n_14),
.B(n_13),
.Y(n_402)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_358),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_10),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_381),
.A2(n_383),
.B1(n_390),
.B2(n_166),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_357),
.A2(n_172),
.B1(n_104),
.B2(n_137),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_365),
.Y(n_384)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_370),
.A2(n_137),
.B1(n_135),
.B2(n_96),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_367),
.A2(n_119),
.B1(n_134),
.B2(n_138),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_350),
.A2(n_119),
.B1(n_134),
.B2(n_11),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_404),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_359),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_393),
.B(n_400),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_353),
.C(n_363),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_387),
.C(n_372),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_395),
.A2(n_381),
.B1(n_382),
.B2(n_390),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_396),
.A2(n_386),
.B1(n_391),
.B2(n_379),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_377),
.A2(n_353),
.B(n_364),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_398),
.A2(n_401),
.B(n_403),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_372),
.B(n_364),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_375),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_10),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_380),
.B(n_375),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_90),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_384),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_405),
.A2(n_166),
.B1(n_125),
.B2(n_33),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_407),
.B(n_413),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_411),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_397),
.A2(n_398),
.B(n_394),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_410),
.A2(n_3),
.B(n_4),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_414),
.A2(n_416),
.B1(n_402),
.B2(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_376),
.C(n_383),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_419),
.C(n_0),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_378),
.B1(n_12),
.B2(n_66),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_125),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_415),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_423),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_424),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_427),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_125),
.Y(n_424)
);

AOI31xp67_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_425),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_436)
);

AO21x1_ASAP7_75t_L g426 ( 
.A1(n_413),
.A2(n_1),
.B(n_3),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_426),
.B(n_6),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_33),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_412),
.C(n_416),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_4),
.B(n_5),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_5),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_432),
.Y(n_446)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_433),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_414),
.Y(n_435)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_435),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_436),
.A2(n_439),
.B(n_426),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_411),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_437),
.A2(n_420),
.B(n_429),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_443),
.Y(n_448)
);

AOI321xp33_ASAP7_75t_SL g445 ( 
.A1(n_440),
.A2(n_429),
.A3(n_8),
.B1(n_9),
.B2(n_6),
.C(n_24),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_445),
.A2(n_433),
.B(n_434),
.C(n_8),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_438),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_450),
.C(n_441),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_446),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_449),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_448),
.C(n_9),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_451),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_9),
.C(n_24),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_455),
.A2(n_24),
.B(n_431),
.Y(n_456)
);


endmodule