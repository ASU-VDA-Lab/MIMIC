module fake_jpeg_24261_n_88 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2x1_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_5),
.B(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_4),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_48),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_7),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_17),
.B(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_58),
.C(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_24),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_41),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_61),
.B1(n_39),
.B2(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_33),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_49),
.B(n_60),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_61),
.C(n_56),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.C(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_71),
.B1(n_70),
.B2(n_69),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_38),
.B(n_36),
.Y(n_74)
);

XNOR2x1_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_38),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_80),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_54),
.B(n_27),
.C(n_64),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_81),
.C(n_63),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_87),
.B(n_24),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_82),
.C(n_62),
.Y(n_87)
);


endmodule