module fake_jpeg_3858_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_32),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_19),
.B1(n_27),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_64),
.Y(n_87)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_21),
.B1(n_27),
.B2(n_17),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_60),
.B(n_65),
.Y(n_95)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_19),
.B1(n_44),
.B2(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_21),
.B1(n_27),
.B2(n_19),
.Y(n_66)
);

NAND2x1p5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_30),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_43),
.B(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_96),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_74),
.B1(n_84),
.B2(n_95),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_67),
.B1(n_91),
.B2(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_121),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_47),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_47),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_53),
.C(n_72),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_123),
.C(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_112),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_120),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_55),
.B1(n_65),
.B2(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_93),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_44),
.B1(n_51),
.B2(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_51),
.B1(n_57),
.B2(n_67),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_70),
.B(n_62),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_62),
.C(n_49),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_130),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_131),
.B1(n_140),
.B2(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_78),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_67),
.B1(n_63),
.B2(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_136),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_78),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_41),
.B1(n_54),
.B2(n_48),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_80),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_24),
.Y(n_179)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_149),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_52),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_107),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_80),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_128),
.B1(n_148),
.B2(n_145),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_157),
.B1(n_164),
.B2(n_165),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_103),
.B1(n_114),
.B2(n_121),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_150),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_163),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_103),
.B1(n_112),
.B2(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_172),
.B1(n_143),
.B2(n_138),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_126),
.B(n_109),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_167),
.B(n_26),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_109),
.B1(n_93),
.B2(n_46),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_154),
.B1(n_133),
.B2(n_140),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_41),
.B1(n_42),
.B2(n_99),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_169),
.B1(n_179),
.B2(n_26),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_42),
.B(n_120),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_102),
.B1(n_119),
.B2(n_110),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_33),
.B1(n_16),
.B2(n_119),
.Y(n_172)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_34),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_34),
.C(n_86),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_157),
.C(n_159),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_182),
.B1(n_61),
.B2(n_90),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_190),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_160),
.C(n_175),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_207),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_171),
.B1(n_156),
.B2(n_155),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_191),
.B1(n_202),
.B2(n_34),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_147),
.B1(n_146),
.B2(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_193),
.B(n_195),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_194),
.A2(n_30),
.B(n_33),
.Y(n_232)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_115),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_201),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_141),
.B1(n_119),
.B2(n_104),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_166),
.C(n_181),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_86),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_24),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_86),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_212),
.C(n_218),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_206),
.C(n_188),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_202),
.B(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_29),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_61),
.C(n_174),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_205),
.B1(n_116),
.B2(n_134),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_180),
.C(n_139),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_225),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_40),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_40),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_228),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_40),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_184),
.B1(n_201),
.B2(n_194),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_137),
.B(n_16),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_230),
.A2(n_232),
.B(n_29),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_68),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_68),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_249),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_183),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_258),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_221),
.B1(n_230),
.B2(n_234),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_134),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_245),
.A2(n_250),
.B(n_9),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_255),
.C(n_217),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_116),
.B1(n_134),
.B2(n_22),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_22),
.B(n_24),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_31),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_31),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_223),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_28),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_213),
.A2(n_28),
.B1(n_1),
.B2(n_3),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_28),
.B1(n_1),
.B2(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_15),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_28),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_232),
.A3(n_233),
.B1(n_219),
.B2(n_218),
.C1(n_225),
.C2(n_210),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_SL g290 ( 
.A(n_259),
.B(n_13),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_264),
.C(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_221),
.C(n_227),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_216),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_8),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_236),
.C(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_237),
.C(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_273),
.C(n_250),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_248),
.B1(n_256),
.B2(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_14),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_215),
.C(n_28),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_238),
.B(n_8),
.Y(n_275)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_260),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_248),
.B1(n_244),
.B2(n_254),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_244),
.B1(n_258),
.B2(n_251),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_291),
.C(n_292),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_287),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_288),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_14),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_263),
.B1(n_265),
.B2(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_261),
.B(n_266),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_0),
.C(n_1),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_13),
.B(n_12),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_302),
.B(n_303),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_3),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_282),
.B(n_291),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_262),
.B1(n_9),
.B2(n_10),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_262),
.B1(n_13),
.B2(n_12),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_4),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_12),
.B(n_11),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_11),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_304),
.A2(n_307),
.B(n_7),
.Y(n_318)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_0),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_293),
.B(n_11),
.Y(n_307)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_311),
.B(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_3),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_4),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_4),
.C(n_5),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_318),
.B(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_300),
.B(n_4),
.Y(n_317)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_303),
.B(n_295),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_322),
.B(n_324),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_321),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_304),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_327),
.A2(n_330),
.B(n_331),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_312),
.B(n_316),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_5),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_6),
.B1(n_7),
.B2(n_322),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

NAND2x1p5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_329),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_332),
.B(n_334),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_6),
.Y(n_338)
);


endmodule