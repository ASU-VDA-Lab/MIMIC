module fake_jpeg_11978_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_23),
.C(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_72),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_0),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_56),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_77),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_80),
.B1(n_58),
.B2(n_61),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_58),
.B1(n_79),
.B2(n_71),
.Y(n_119)
);

NAND2xp67_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_54),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_67),
.B1(n_78),
.B2(n_73),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_79),
.B1(n_70),
.B2(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_104),
.Y(n_108)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_76),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_114),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_97),
.B(n_84),
.C(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_62),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_55),
.B1(n_62),
.B2(n_80),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_57),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_126),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_75),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_59),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_74),
.B(n_66),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_137),
.B(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_25),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_117),
.B1(n_123),
.B2(n_121),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_143),
.B1(n_43),
.B2(n_15),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_11),
.Y(n_165)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_55),
.B1(n_60),
.B2(n_4),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_149),
.B1(n_7),
.B2(n_8),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_24),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_146),
.B(n_144),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_156),
.C(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_5),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_51),
.C(n_30),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_6),
.B(n_7),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_161),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_168),
.B1(n_133),
.B2(n_140),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_8),
.B(n_10),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_177),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_13),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_180),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_150),
.B1(n_171),
.B2(n_172),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_170),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_189),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_166),
.B1(n_169),
.B2(n_181),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_167),
.C(n_20),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_192),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_182),
.B(n_173),
.CI(n_176),
.CON(n_192),
.SN(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_190),
.Y(n_197)
);

OA21x2_ASAP7_75t_SL g198 ( 
.A1(n_197),
.A2(n_192),
.B(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_188),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_199),
.A2(n_187),
.B1(n_194),
.B2(n_186),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_189),
.B(n_21),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_19),
.C(n_35),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_36),
.B(n_38),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_41),
.Y(n_204)
);


endmodule