module fake_jpeg_1320_n_356 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_64),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_25),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_68),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_6),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_75),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_77),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_37),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_40),
.B1(n_39),
.B2(n_15),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_95),
.B1(n_105),
.B2(n_110),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_23),
.B1(n_34),
.B2(n_33),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_49),
.B1(n_73),
.B2(n_62),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_104),
.A2(n_84),
.B(n_113),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_121),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_15),
.B1(n_39),
.B2(n_30),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_15),
.B1(n_39),
.B2(n_30),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_30),
.B1(n_28),
.B2(n_36),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_47),
.A2(n_32),
.B1(n_38),
.B2(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_38),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_125),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_47),
.A2(n_32),
.B1(n_27),
.B2(n_37),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_27),
.B1(n_21),
.B2(n_41),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_18),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_41),
.C(n_21),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_69),
.A2(n_18),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_42),
.A2(n_45),
.B1(n_61),
.B2(n_54),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_43),
.B(n_5),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_3),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_50),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_52),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_130),
.B(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_114),
.B1(n_81),
.B2(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_132),
.A2(n_140),
.B1(n_169),
.B2(n_168),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_137),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_72),
.B(n_70),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_138),
.B(n_164),
.C(n_152),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_166),
.B1(n_128),
.B2(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_10),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_103),
.B1(n_127),
.B2(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_149),
.A2(n_171),
.B1(n_135),
.B2(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_153),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_2),
.B(n_3),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_171),
.B(n_132),
.C(n_165),
.Y(n_193)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_4),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_160),
.Y(n_181)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_85),
.B(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_162),
.Y(n_201)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_87),
.B(n_107),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_107),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_127),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_99),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_167),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_101),
.B1(n_104),
.B2(n_87),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_169),
.Y(n_210)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_86),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_172),
.Y(n_190)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_182),
.B1(n_188),
.B2(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_102),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_191),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_129),
.B1(n_161),
.B2(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_138),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_193),
.A2(n_208),
.B(n_202),
.C(n_190),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_137),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_199),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_137),
.B(n_148),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_207),
.B1(n_176),
.B2(n_211),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_167),
.B1(n_156),
.B2(n_158),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_196),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_191),
.A2(n_146),
.B1(n_173),
.B2(n_200),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_213),
.A2(n_214),
.B(n_238),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_197),
.B(n_185),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_199),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_201),
.B1(n_212),
.B2(n_194),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_218),
.A2(n_220),
.B1(n_241),
.B2(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_175),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_212),
.A2(n_181),
.B1(n_187),
.B2(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_175),
.B(n_177),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_225),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_179),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_186),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_231),
.Y(n_266)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_229),
.Y(n_250)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_176),
.A2(n_190),
.B1(n_208),
.B2(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_237),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_189),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_198),
.B(n_202),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_238),
.B(n_214),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_184),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_174),
.B(n_198),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_204),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_197),
.B1(n_191),
.B2(n_200),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_252),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_257),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_260),
.C(n_263),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_224),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_218),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_268),
.A2(n_236),
.B(n_223),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_217),
.C(n_213),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_260),
.C(n_249),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_216),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_282),
.C(n_265),
.Y(n_308)
);

BUFx12_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_233),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_279),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_238),
.B(n_226),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_280),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_237),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_246),
.C(n_245),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_238),
.B1(n_222),
.B2(n_231),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_229),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_285),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_238),
.B1(n_230),
.B2(n_223),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_269),
.B1(n_250),
.B2(n_265),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_247),
.B(n_258),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_292),
.B(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_270),
.B(n_248),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_251),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_294),
.Y(n_313)
);

XOR2x2_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_271),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_272),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_252),
.B1(n_254),
.B2(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_302),
.B1(n_309),
.B2(n_277),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_254),
.B1(n_264),
.B2(n_267),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_261),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_307),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_250),
.B(n_261),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_308),
.B(n_281),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_269),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_273),
.B1(n_277),
.B2(n_286),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_317),
.Y(n_334)
);

BUFx12f_ASAP7_75t_SL g311 ( 
.A(n_297),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_311),
.A2(n_298),
.B(n_302),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_323),
.B1(n_276),
.B2(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

AOI221xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_273),
.B1(n_292),
.B2(n_276),
.C(n_291),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_316),
.B(n_321),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_307),
.C(n_295),
.Y(n_326)
);

BUFx12_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_320),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_303),
.C(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_329),
.Y(n_336)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_301),
.C(n_306),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_304),
.C(n_293),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_332),
.B(n_315),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_313),
.B(n_315),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_339),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_338),
.Y(n_344)
);

BUFx4f_ASAP7_75t_SL g340 ( 
.A(n_330),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_326),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_329),
.C(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_331),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_347),
.B(n_339),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_350),
.C(n_347),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_351),
.A2(n_352),
.A3(n_311),
.B1(n_340),
.B2(n_336),
.C1(n_333),
.C2(n_320),
.Y(n_353)
);

OAI31xp33_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_343),
.A3(n_345),
.B(n_335),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

AOI221xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_332),
.B1(n_324),
.B2(n_342),
.C(n_283),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_324),
.Y(n_356)
);


endmodule