module fake_jpeg_24014_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_2),
.B(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_51),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_24),
.B1(n_27),
.B2(n_21),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_53),
.B1(n_18),
.B2(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_24),
.B1(n_17),
.B2(n_12),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_21),
.B(n_13),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_5),
.B(n_7),
.Y(n_74)
);

NOR4xp25_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_58),
.B(n_62),
.C(n_54),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_27),
.B1(n_13),
.B2(n_15),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_15),
.C(n_22),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_72),
.B1(n_77),
.B2(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_23),
.B1(n_18),
.B2(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_4),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_80),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_78),
.B(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_5),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_83),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_5),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_46),
.B(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_6),
.B1(n_49),
.B2(n_44),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_64),
.B(n_60),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_95),
.B1(n_96),
.B2(n_73),
.Y(n_104)
);

CKINVDCx10_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_94),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_69),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_74),
.B1(n_68),
.B2(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_105),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_107),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_90),
.B(n_86),
.Y(n_111)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_71),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_91),
.B(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_83),
.B1(n_88),
.B2(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_104),
.B1(n_102),
.B2(n_97),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_95),
.B(n_90),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_111),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_100),
.Y(n_118)
);

OAI322xp33_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_97),
.A3(n_76),
.B1(n_75),
.B2(n_70),
.C1(n_69),
.C2(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_99),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_118),
.C(n_120),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_114),
.B1(n_112),
.B2(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_103),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_110),
.C(n_109),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.C(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_121),
.B(n_106),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_129),
.B(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_89),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_130),
.A2(n_131),
.B(n_105),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_81),
.B(n_50),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_82),
.Y(n_134)
);


endmodule