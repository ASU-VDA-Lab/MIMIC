module fake_jpeg_5474_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_12),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_56),
.B1(n_53),
.B2(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_63),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_54),
.B(n_57),
.C(n_50),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_49),
.B(n_51),
.C(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_58),
.B1(n_41),
.B2(n_46),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_69),
.B1(n_47),
.B2(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_15),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_68),
.B1(n_9),
.B2(n_11),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_83),
.B1(n_17),
.B2(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_84),
.C(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_86),
.Y(n_92)
);

NAND4xp25_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_21),
.C(n_22),
.D(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_25),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_36),
.C(n_37),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_38),
.Y(n_99)
);


endmodule