module fake_netlist_1_10641_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
NOR2xp33_ASAP7_75t_L g7 ( .A(n_6), .B(n_4), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_2), .B(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx5_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_14), .B(n_13), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
NOR3xp33_ASAP7_75t_L g17 ( .A(n_16), .B(n_8), .C(n_11), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_17), .B(n_7), .C(n_12), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_18), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
endmodule