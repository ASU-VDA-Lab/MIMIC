module fake_jpeg_2303_n_394 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_394);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_394;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_53),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_67),
.Y(n_88)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_8),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_68),
.Y(n_98)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_65),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_29),
.B(n_10),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_75),
.Y(n_100)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_0),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_23),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_29),
.B(n_13),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_81),
.Y(n_108)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_80),
.Y(n_131)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_82),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_11),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_84),
.Y(n_110)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_37),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_78),
.B1(n_66),
.B2(n_46),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_87),
.A2(n_5),
.B1(n_12),
.B2(n_120),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_20),
.B1(n_18),
.B2(n_37),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_103),
.B1(n_129),
.B2(n_69),
.Y(n_138)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_42),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_36),
.B1(n_28),
.B2(n_16),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_15),
.CON(n_107),
.SN(n_107)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_36),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_26),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_26),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_20),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_52),
.B(n_23),
.C(n_18),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_82),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_15),
.B1(n_40),
.B2(n_35),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_48),
.A2(n_15),
.B1(n_40),
.B2(n_35),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_65),
.B1(n_74),
.B2(n_4),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_138),
.A2(n_149),
.B1(n_159),
.B2(n_163),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_65),
.B1(n_79),
.B2(n_58),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_144),
.B(n_90),
.C(n_93),
.Y(n_182)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_74),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_175),
.B1(n_135),
.B2(n_117),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_12),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_99),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_110),
.B1(n_96),
.B2(n_127),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_169),
.Y(n_196)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_134),
.B1(n_98),
.B2(n_87),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_167),
.A2(n_171),
.B1(n_93),
.B2(n_122),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_88),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_168),
.B(n_173),
.Y(n_211)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_99),
.A2(n_106),
.B1(n_132),
.B2(n_107),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_100),
.A2(n_86),
.B1(n_126),
.B2(n_88),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_116),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_150),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_182),
.A2(n_139),
.B(n_170),
.C(n_146),
.Y(n_228)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_118),
.A3(n_99),
.B1(n_121),
.B2(n_95),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_153),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_86),
.B1(n_126),
.B2(n_114),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_201),
.B1(n_197),
.B2(n_173),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_136),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_199),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_95),
.B1(n_117),
.B2(n_135),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_186),
.B1(n_209),
.B2(n_189),
.Y(n_224)
);

NAND2x1_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_122),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_214),
.B(n_180),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_139),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_170),
.B(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_148),
.B(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_151),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_170),
.B(n_144),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_161),
.B(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_183),
.B1(n_203),
.B2(n_181),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_223),
.B(n_247),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_228),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_226),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_248),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_230),
.A2(n_237),
.B(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_164),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_186),
.B(n_155),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_240),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_157),
.C(n_169),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_204),
.C(n_207),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_139),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_179),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_244),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_209),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_211),
.B(n_189),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_183),
.A2(n_191),
.B(n_204),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_190),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_200),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_188),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_192),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_206),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_268),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_257),
.B1(n_272),
.B2(n_238),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_200),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_261),
.C(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_229),
.A2(n_182),
.B1(n_201),
.B2(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_202),
.C(n_195),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_202),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

OAI22x1_ASAP7_75t_SL g272 ( 
.A1(n_228),
.A2(n_212),
.B1(n_210),
.B2(n_207),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_223),
.B(n_188),
.CI(n_212),
.CON(n_273),
.SN(n_273)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_274),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_278),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_234),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_229),
.B(n_250),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_289),
.B1(n_299),
.B2(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_224),
.B1(n_236),
.B2(n_221),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_275),
.A2(n_252),
.B1(n_241),
.B2(n_230),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_264),
.B1(n_266),
.B2(n_268),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_236),
.B(n_249),
.Y(n_292)
);

BUFx4f_ASAP7_75t_SL g325 ( 
.A(n_292),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_258),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_293),
.B(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_302),
.C(n_225),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_304),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_240),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_248),
.B(n_228),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_308),
.B(n_301),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_309),
.A2(n_316),
.B1(n_317),
.B2(n_284),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_278),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_310),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_266),
.B1(n_276),
.B2(n_280),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_311),
.A2(n_313),
.B1(n_315),
.B2(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_265),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_320),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_272),
.B1(n_253),
.B2(n_255),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_265),
.B1(n_261),
.B2(n_273),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_232),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_277),
.C(n_226),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_273),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_306),
.A2(n_304),
.B(n_295),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_320),
.B1(n_307),
.B2(n_310),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_286),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_332),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_286),
.C(n_291),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_344),
.C(n_319),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_333),
.A2(n_312),
.B1(n_326),
.B2(n_321),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_303),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_335),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_323),
.B(n_244),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_342),
.C(n_318),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_227),
.Y(n_340)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_322),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_305),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_208),
.Y(n_343)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_235),
.C(n_288),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_345),
.A2(n_349),
.B1(n_339),
.B2(n_338),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_334),
.Y(n_359)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_270),
.C(n_326),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_351),
.B(n_208),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_355),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g355 ( 
.A(n_331),
.B(n_294),
.CI(n_282),
.CON(n_355),
.SN(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_321),
.C(n_247),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_210),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_366),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_363),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_355),
.A2(n_327),
.B(n_332),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_362),
.A2(n_364),
.B(n_365),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_347),
.A2(n_335),
.B1(n_337),
.B2(n_222),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_353),
.A2(n_344),
.B(n_259),
.Y(n_364)
);

OAI221xp5_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_233),
.B1(n_245),
.B2(n_220),
.C(n_231),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_259),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_210),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_347),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_357),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_369),
.B(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_361),
.B(n_352),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_374),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_377),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_360),
.B(n_351),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_350),
.C(n_243),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_366),
.C(n_363),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_379),
.B(n_373),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_375),
.A2(n_367),
.B(n_243),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_380),
.A2(n_243),
.B(n_384),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_372),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_386),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_378),
.C(n_376),
.Y(n_387)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_387),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_389),
.B(n_382),
.C(n_381),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_SL g393 ( 
.A(n_392),
.B(n_390),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_388),
.Y(n_394)
);


endmodule