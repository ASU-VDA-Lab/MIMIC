module fake_jpeg_2841_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

AND2x6_ASAP7_75t_L g5 ( 
.A(n_3),
.B(n_0),
.Y(n_5)
);

AND2x2_ASAP7_75t_L g6 ( 
.A(n_0),
.B(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_2),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

O2A1O1Ixp33_ASAP7_75t_SL g11 ( 
.A1(n_9),
.A2(n_10),
.B(n_8),
.C(n_1),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_6),
.C(n_8),
.Y(n_10)
);


endmodule