module fake_jpeg_5939_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_42),
.Y(n_56)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx2_ASAP7_75t_SL g65 ( 
.A(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_33),
.B1(n_26),
.B2(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_47),
.B1(n_31),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_33),
.B1(n_20),
.B2(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_55),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_42),
.C(n_17),
.Y(n_84)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_67),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_57),
.B1(n_27),
.B2(n_19),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_78),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_34),
.B(n_42),
.C(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_45),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_32),
.B(n_62),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_69),
.B(n_76),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_24),
.B(n_18),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_29),
.B(n_23),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_43),
.B1(n_60),
.B2(n_49),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_105),
.B1(n_109),
.B2(n_74),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_18),
.B1(n_19),
.B2(n_27),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_36),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_113),
.C(n_80),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_43),
.B1(n_36),
.B2(n_67),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_43),
.B1(n_36),
.B2(n_54),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_82),
.B(n_68),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_52),
.B1(n_64),
.B2(n_59),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_52),
.B1(n_64),
.B2(n_59),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_50),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_37),
.C(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_118),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_137),
.B(n_94),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_73),
.B1(n_75),
.B2(n_88),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_123),
.B1(n_125),
.B2(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_134),
.C(n_99),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_130),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g126 ( 
.A(n_108),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_69),
.B1(n_75),
.B2(n_68),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_106),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_76),
.B1(n_77),
.B2(n_70),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_77),
.C(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_82),
.B(n_28),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_81),
.B1(n_55),
.B2(n_38),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_144),
.C(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_143),
.Y(n_178)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_98),
.C(n_101),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_148),
.B(n_153),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_97),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_100),
.C(n_96),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_131),
.C(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_152),
.C(n_162),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_100),
.C(n_96),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_111),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_163),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_97),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_93),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_50),
.A3(n_25),
.B1(n_89),
.B2(n_28),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_114),
.B1(n_130),
.B2(n_117),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_187),
.B1(n_22),
.B2(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_185),
.C(n_148),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_114),
.B1(n_124),
.B2(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_173),
.B1(n_176),
.B2(n_179),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_129),
.B1(n_128),
.B2(n_25),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_129),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_145),
.B(n_159),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_25),
.B1(n_28),
.B2(n_37),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_150),
.B1(n_155),
.B2(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_181),
.A2(n_189),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_28),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_165),
.B(n_22),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_162),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_191),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_149),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_178),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_180),
.B(n_182),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_200),
.C(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_148),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_180),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_143),
.B1(n_158),
.B2(n_141),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_203),
.B1(n_187),
.B2(n_168),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_141),
.C(n_22),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_22),
.C(n_1),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_0),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_208),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_15),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_210),
.C(n_170),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_179),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_173),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_15),
.C(n_6),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_189),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_183),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_223),
.B(n_227),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_225),
.C(n_191),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_176),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_176),
.B1(n_210),
.B2(n_192),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_201),
.B(n_194),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_237),
.C(n_214),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_224),
.CI(n_216),
.CON(n_241),
.SN(n_241)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_205),
.B1(n_200),
.B2(n_190),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_240),
.B1(n_9),
.B2(n_10),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_202),
.C(n_207),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_239),
.B(n_236),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_220),
.B(n_4),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_250),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_216),
.B(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_219),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_246),
.C(n_251),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_7),
.C(n_9),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

AOI21x1_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_10),
.B(n_11),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_12),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_10),
.C(n_11),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_11),
.C(n_12),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_236),
.B1(n_234),
.B2(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_234),
.B1(n_231),
.B2(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_256),
.B(n_249),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_232),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_262),
.B(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_245),
.C(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_241),
.B(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_252),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_252),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_258),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_256),
.B(n_257),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_270),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_259),
.B(n_272),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_277),
.B(n_243),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_279),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_14),
.Y(n_281)
);


endmodule