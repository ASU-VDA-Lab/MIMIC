module real_aes_15520_n_361 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_1957, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_361);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_1957;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_361;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1632;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1638;
wire n_495;
wire n_1078;
wire n_1072;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_1942;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_0), .A2(n_284), .B1(n_1139), .B2(n_1501), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_0), .A2(n_247), .B1(n_483), .B2(n_1519), .Y(n_1518) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_1), .A2(n_114), .B1(n_507), .B2(n_511), .Y(n_1349) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_1), .A2(n_189), .B1(n_432), .B2(n_435), .Y(n_1384) );
AND2x2_ASAP7_75t_L g464 ( .A(n_2), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g478 ( .A(n_2), .B(n_255), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_2), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g547 ( .A(n_2), .Y(n_547) );
INVx1_ASAP7_75t_L g1119 ( .A(n_3), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_3), .A2(n_77), .B1(n_385), .B2(n_1133), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_4), .A2(n_274), .B1(n_633), .B2(n_637), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_4), .A2(n_274), .B1(n_670), .B2(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g940 ( .A(n_5), .Y(n_940) );
INVx1_ASAP7_75t_L g1108 ( .A(n_6), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g1687 ( .A1(n_7), .A2(n_206), .B1(n_1674), .B2(n_1688), .Y(n_1687) );
INVxp67_ASAP7_75t_SL g924 ( .A(n_8), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_8), .A2(n_121), .B1(n_875), .B2(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g922 ( .A(n_9), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_9), .A2(n_168), .B1(n_440), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g1503 ( .A1(n_10), .A2(n_211), .B1(n_704), .B2(n_713), .Y(n_1503) );
AOI221xp5_ASAP7_75t_L g1516 ( .A1(n_10), .A2(n_118), .B1(n_985), .B2(n_1329), .C(n_1517), .Y(n_1516) );
AOI22xp33_ASAP7_75t_L g1708 ( .A1(n_11), .A2(n_89), .B1(n_1674), .B2(n_1678), .Y(n_1708) );
AOI22xp33_ASAP7_75t_L g1771 ( .A1(n_12), .A2(n_345), .B1(n_1681), .B2(n_1684), .Y(n_1771) );
INVx1_ASAP7_75t_L g625 ( .A(n_13), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g1155 ( .A1(n_14), .A2(n_352), .B1(n_385), .B2(n_390), .C(n_396), .Y(n_1155) );
OAI21xp33_ASAP7_75t_SL g1185 ( .A1(n_14), .A2(n_501), .B(n_753), .Y(n_1185) );
INVx2_ASAP7_75t_L g381 ( .A(n_15), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_16), .A2(n_168), .B1(n_483), .B2(n_936), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_16), .A2(n_320), .B1(n_964), .B2(n_966), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g1278 ( .A(n_17), .Y(n_1278) );
INVx1_ASAP7_75t_L g565 ( .A(n_18), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_19), .A2(n_297), .B1(n_432), .B2(n_435), .Y(n_1168) );
INVx1_ASAP7_75t_L g1184 ( .A(n_19), .Y(n_1184) );
INVx1_ASAP7_75t_L g824 ( .A(n_20), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_21), .A2(n_617), .B(n_618), .C(n_624), .Y(n_616) );
INVx1_ASAP7_75t_L g668 ( .A(n_21), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_22), .A2(n_351), .B1(n_418), .B2(n_1462), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_22), .A2(n_166), .B1(n_734), .B2(n_835), .Y(n_1476) );
XOR2x1_ASAP7_75t_L g1397 ( .A(n_23), .B(n_1398), .Y(n_1397) );
AOI22xp5_ASAP7_75t_L g1680 ( .A1(n_23), .A2(n_217), .B1(n_1681), .B2(n_1684), .Y(n_1680) );
INVx1_ASAP7_75t_L g1225 ( .A(n_24), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g1241 ( .A1(n_24), .A2(n_151), .B1(n_441), .B2(n_1242), .C(n_1245), .Y(n_1241) );
INVx1_ASAP7_75t_L g1075 ( .A(n_25), .Y(n_1075) );
AOI221x1_ASAP7_75t_SL g1080 ( .A1(n_25), .A2(n_201), .B1(n_483), .B2(n_1002), .C(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g581 ( .A(n_26), .Y(n_581) );
OA22x2_ASAP7_75t_L g1529 ( .A1(n_27), .A2(n_1530), .B1(n_1593), .B2(n_1594), .Y(n_1529) );
INVxp67_ASAP7_75t_L g1594 ( .A(n_27), .Y(n_1594) );
HB1xp67_ASAP7_75t_L g1661 ( .A(n_28), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_28), .B(n_1659), .Y(n_1675) );
AOI22xp33_ASAP7_75t_L g1769 ( .A1(n_29), .A2(n_190), .B1(n_1674), .B2(n_1770), .Y(n_1769) );
AOI22xp33_ASAP7_75t_L g1722 ( .A1(n_30), .A2(n_203), .B1(n_1674), .B2(n_1678), .Y(n_1722) );
INVx1_ASAP7_75t_L g1071 ( .A(n_31), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_31), .A2(n_181), .B1(n_622), .B2(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1552 ( .A(n_32), .Y(n_1552) );
INVx1_ASAP7_75t_L g692 ( .A(n_33), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_33), .A2(n_58), .B1(n_755), .B2(n_756), .Y(n_754) );
OAI211xp5_ASAP7_75t_SL g820 ( .A1(n_34), .A2(n_821), .B(n_823), .C(n_828), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_34), .A2(n_282), .B1(n_901), .B2(n_903), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_35), .A2(n_262), .B1(n_402), .B2(n_409), .Y(n_1404) );
INVxp33_ASAP7_75t_L g1447 ( .A(n_35), .Y(n_1447) );
INVx1_ASAP7_75t_L g1231 ( .A(n_36), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_36), .A2(n_48), .B1(n_385), .B2(n_390), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_37), .A2(n_247), .B1(n_1139), .B2(n_1501), .Y(n_1500) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_37), .A2(n_284), .B1(n_727), .B2(n_802), .C(n_1004), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_38), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_38), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_39), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_40), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_40), .A2(n_88), .B1(n_875), .B2(n_962), .Y(n_967) );
INVx1_ASAP7_75t_L g782 ( .A(n_41), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_42), .A2(n_409), .B1(n_1265), .B2(n_1268), .Y(n_1264) );
INVx1_ASAP7_75t_L g1283 ( .A(n_42), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1495 ( .A(n_43), .Y(n_1495) );
INVx1_ASAP7_75t_L g779 ( .A(n_44), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g806 ( .A1(n_44), .A2(n_271), .B1(n_802), .B2(n_807), .C(n_808), .Y(n_806) );
OAI221xp5_ASAP7_75t_L g838 ( .A1(n_45), .A2(n_120), .B1(n_839), .B2(n_843), .C(n_847), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_45), .A2(n_120), .B1(n_887), .B2(n_889), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_46), .A2(n_194), .B1(n_483), .B2(n_937), .Y(n_1005) );
INVx1_ASAP7_75t_L g1035 ( .A(n_46), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1354 ( .A1(n_47), .A2(n_63), .B1(n_609), .B2(n_1355), .C(n_1357), .Y(n_1354) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_47), .A2(n_141), .B1(n_875), .B2(n_1376), .C(n_1382), .Y(n_1381) );
OAI221xp5_ASAP7_75t_L g1227 ( .A1(n_48), .A2(n_312), .B1(n_501), .B2(n_756), .C(n_1093), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_49), .A2(n_259), .B1(n_855), .B2(n_856), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_49), .A2(n_354), .B1(n_862), .B2(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g1466 ( .A1(n_50), .A2(n_131), .B1(n_907), .B2(n_1467), .Y(n_1466) );
INVxp67_ASAP7_75t_SL g1486 ( .A(n_50), .Y(n_1486) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_51), .A2(n_167), .B1(n_1674), .B2(n_1678), .Y(n_1695) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_52), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_53), .A2(n_337), .B1(n_414), .B2(n_712), .C(n_714), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_53), .A2(n_174), .B1(n_721), .B2(n_725), .Y(n_720) );
INVx1_ASAP7_75t_L g1507 ( .A(n_54), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_55), .A2(n_202), .B1(n_402), .B2(n_409), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_55), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g1220 ( .A(n_56), .Y(n_1220) );
INVx1_ASAP7_75t_L g1271 ( .A(n_57), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_57), .A2(n_60), .B1(n_932), .B2(n_937), .Y(n_1292) );
INVx1_ASAP7_75t_L g717 ( .A(n_58), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_59), .A2(n_222), .B1(n_936), .B2(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1029 ( .A(n_59), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1259 ( .A1(n_60), .A2(n_344), .B1(n_964), .B2(n_1244), .C(n_1260), .Y(n_1259) );
OAI222xp33_ASAP7_75t_L g1901 ( .A1(n_61), .A2(n_78), .B1(n_1638), .B2(n_1902), .C1(n_1903), .C2(n_1908), .Y(n_1901) );
INVx1_ASAP7_75t_L g1927 ( .A(n_61), .Y(n_1927) );
INVxp67_ASAP7_75t_SL g1229 ( .A(n_62), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_62), .A2(n_409), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
INVx1_ASAP7_75t_L g1378 ( .A(n_63), .Y(n_1378) );
AOI22xp33_ASAP7_75t_SL g1318 ( .A1(n_64), .A2(n_175), .B1(n_1309), .B2(n_1319), .Y(n_1318) );
AOI221xp5_ASAP7_75t_L g1336 ( .A1(n_64), .A2(n_128), .B1(n_830), .B2(n_1337), .C(n_1339), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_65), .A2(n_294), .B1(n_402), .B2(n_409), .Y(n_783) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_65), .Y(n_786) );
INVx1_ASAP7_75t_L g1323 ( .A(n_66), .Y(n_1323) );
AOI21xp33_ASAP7_75t_L g1169 ( .A1(n_67), .A2(n_1170), .B(n_1173), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_67), .A2(n_109), .B1(n_1197), .B2(n_1198), .C(n_1199), .Y(n_1196) );
INVx1_ASAP7_75t_L g693 ( .A(n_68), .Y(n_693) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_68), .A2(n_501), .B(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1944 ( .A1(n_69), .A2(n_1899), .B1(n_1945), .B2(n_1946), .Y(n_1944) );
CKINVDCx5p33_ASAP7_75t_R g1946 ( .A(n_69), .Y(n_1946) );
INVx1_ASAP7_75t_L g1233 ( .A(n_70), .Y(n_1233) );
OAI222xp33_ASAP7_75t_L g1236 ( .A1(n_70), .A2(n_301), .B1(n_312), .B2(n_406), .C1(n_423), .C2(n_1237), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1369 ( .A(n_71), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_71), .A2(n_110), .B1(n_402), .B2(n_409), .Y(n_1373) );
INVx1_ASAP7_75t_L g1325 ( .A(n_72), .Y(n_1325) );
INVx1_ASAP7_75t_L g1457 ( .A(n_73), .Y(n_1457) );
AOI21xp33_ASAP7_75t_L g850 ( .A1(n_74), .A2(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g866 ( .A(n_74), .Y(n_866) );
XOR2x2_ASAP7_75t_L g1150 ( .A(n_75), .B(n_1151), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1620 ( .A1(n_76), .A2(n_327), .B1(n_768), .B2(n_1621), .Y(n_1620) );
AOI221xp5_ASAP7_75t_L g1632 ( .A1(n_76), .A2(n_341), .B1(n_851), .B2(n_1329), .C(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1113 ( .A(n_77), .Y(n_1113) );
INVx1_ASAP7_75t_L g1928 ( .A(n_78), .Y(n_1928) );
OAI22xp33_ASAP7_75t_L g1545 ( .A1(n_79), .A2(n_191), .B1(n_1546), .B2(n_1547), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g1586 ( .A1(n_79), .A2(n_191), .B1(n_1587), .B2(n_1589), .Y(n_1586) );
XNOR2xp5_ASAP7_75t_L g1449 ( .A(n_80), .B(n_1450), .Y(n_1449) );
NAND2xp33_ASAP7_75t_SL g1353 ( .A(n_81), .B(n_604), .Y(n_1353) );
INVx1_ASAP7_75t_L g1383 ( .A(n_81), .Y(n_1383) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_82), .A2(n_129), .B1(n_521), .B2(n_982), .C(n_983), .Y(n_981) );
INVx1_ASAP7_75t_L g1014 ( .A(n_82), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_83), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_84), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g1417 ( .A1(n_85), .A2(n_204), .B1(n_432), .B2(n_435), .Y(n_1417) );
INVxp67_ASAP7_75t_SL g1431 ( .A(n_85), .Y(n_1431) );
XOR2xp5_ASAP7_75t_L g1491 ( .A(n_86), .B(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1567 ( .A(n_87), .Y(n_1567) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_88), .A2(n_121), .B1(n_798), .B2(n_833), .C(n_851), .Y(n_934) );
INVx1_ASAP7_75t_L g986 ( .A(n_90), .Y(n_986) );
OAI221xp5_ASAP7_75t_SL g1019 ( .A1(n_90), .A2(n_125), .B1(n_388), .B2(n_443), .C(n_892), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_91), .A2(n_332), .B1(n_438), .B2(n_441), .C(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g553 ( .A(n_91), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_92), .A2(n_215), .B1(n_402), .B2(n_409), .Y(n_1156) );
INVxp67_ASAP7_75t_SL g1195 ( .A(n_92), .Y(n_1195) );
INVx1_ASAP7_75t_L g1298 ( .A(n_93), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_94), .B(n_1314), .Y(n_1416) );
AOI221xp5_ASAP7_75t_L g1445 ( .A1(n_94), .A2(n_226), .B1(n_609), .B2(n_734), .C(n_835), .Y(n_1445) );
AOI22xp5_ASAP7_75t_L g1699 ( .A1(n_95), .A2(n_216), .B1(n_1681), .B2(n_1684), .Y(n_1699) );
INVx1_ASAP7_75t_L g1522 ( .A(n_96), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_97), .A2(n_324), .B1(n_713), .B2(n_1314), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_97), .A2(n_147), .B1(n_730), .B2(n_1332), .Y(n_1335) );
AOI222xp33_ASAP7_75t_L g1174 ( .A1(n_98), .A2(n_159), .B1(n_340), .B2(n_411), .C1(n_418), .C2(n_699), .Y(n_1174) );
INVx1_ASAP7_75t_L g1200 ( .A(n_98), .Y(n_1200) );
CKINVDCx5p33_ASAP7_75t_R g1221 ( .A(n_99), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_100), .B(n_1412), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_100), .A2(n_178), .B1(n_807), .B2(n_1198), .Y(n_1444) );
INVx1_ASAP7_75t_L g774 ( .A(n_101), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_101), .A2(n_198), .B1(n_798), .B2(n_800), .C(n_803), .Y(n_797) );
INVx1_ASAP7_75t_L g1304 ( .A(n_102), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1460 ( .A1(n_103), .A2(n_199), .B1(n_768), .B2(n_882), .Y(n_1460) );
INVxp67_ASAP7_75t_SL g1485 ( .A(n_103), .Y(n_1485) );
OAI22xp33_ASAP7_75t_L g1279 ( .A1(n_104), .A2(n_155), .B1(n_385), .B2(n_390), .Y(n_1279) );
OAI22xp5_ASAP7_75t_L g1293 ( .A1(n_104), .A2(n_300), .B1(n_756), .B2(n_1093), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g1909 ( .A(n_105), .Y(n_1909) );
AOI22xp33_ASAP7_75t_SL g1933 ( .A1(n_105), .A2(n_288), .B1(n_875), .B2(n_1467), .Y(n_1933) );
INVx1_ASAP7_75t_L g1568 ( .A(n_106), .Y(n_1568) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_107), .Y(n_1226) );
OAI221xp5_ASAP7_75t_L g1603 ( .A1(n_108), .A2(n_236), .B1(n_969), .B2(n_1604), .C(n_1605), .Y(n_1603) );
OAI211xp5_ASAP7_75t_L g1628 ( .A1(n_108), .A2(n_1483), .B(n_1629), .C(n_1634), .Y(n_1628) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_109), .A2(n_229), .B1(n_1159), .B2(n_1161), .C(n_1163), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1389 ( .A(n_110), .Y(n_1389) );
INVx1_ASAP7_75t_L g1659 ( .A(n_111), .Y(n_1659) );
INVx1_ASAP7_75t_L g1267 ( .A(n_112), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_112), .A2(n_344), .B1(n_483), .B2(n_937), .Y(n_1289) );
INVx1_ASAP7_75t_L g1230 ( .A(n_113), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_114), .A2(n_139), .B1(n_385), .B2(n_390), .C(n_396), .Y(n_1372) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_115), .A2(n_160), .B1(n_833), .B2(n_1002), .C(n_1003), .Y(n_1006) );
INVx1_ASAP7_75t_L g1024 ( .A(n_115), .Y(n_1024) );
INVx1_ASAP7_75t_L g1154 ( .A(n_116), .Y(n_1154) );
OAI21xp33_ASAP7_75t_L g1181 ( .A1(n_116), .A2(n_1098), .B(n_1182), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1626 ( .A1(n_117), .A2(n_268), .B1(n_903), .B2(n_1343), .Y(n_1626) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_118), .A2(n_254), .B1(n_1310), .B2(n_1499), .Y(n_1498) );
INVx1_ASAP7_75t_L g573 ( .A(n_119), .Y(n_573) );
XOR2x2_ASAP7_75t_L g366 ( .A(n_122), .B(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g1308 ( .A1(n_123), .A2(n_128), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_123), .A2(n_311), .B1(n_985), .B2(n_1198), .C(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1361 ( .A(n_124), .Y(n_1361) );
INVx1_ASAP7_75t_L g997 ( .A(n_125), .Y(n_997) );
INVx1_ASAP7_75t_L g1048 ( .A(n_126), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_126), .A2(n_251), .B1(n_756), .B2(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1920 ( .A(n_127), .Y(n_1920) );
INVx1_ASAP7_75t_L g1011 ( .A(n_129), .Y(n_1011) );
INVx1_ASAP7_75t_L g430 ( .A(n_130), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_131), .A2(n_199), .B1(n_1329), .B2(n_1337), .C(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g446 ( .A(n_132), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g1342 ( .A1(n_133), .A2(n_1343), .B(n_1344), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_134), .A2(n_240), .B1(n_835), .B2(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g870 ( .A(n_134), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g1704 ( .A1(n_135), .A2(n_323), .B1(n_1681), .B2(n_1684), .Y(n_1704) );
INVx1_ASAP7_75t_L g444 ( .A(n_136), .Y(n_444) );
INVx1_ASAP7_75t_L g992 ( .A(n_137), .Y(n_992) );
OAI21xp33_ASAP7_75t_L g1017 ( .A1(n_137), .A2(n_896), .B(n_1018), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g1262 ( .A(n_138), .Y(n_1262) );
INVxp67_ASAP7_75t_SL g1368 ( .A(n_139), .Y(n_1368) );
OAI221xp5_ASAP7_75t_L g1403 ( .A1(n_140), .A2(n_321), .B1(n_385), .B2(n_390), .C(n_396), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1435 ( .A(n_140), .B(n_488), .Y(n_1435) );
AOI221xp5_ASAP7_75t_L g1362 ( .A1(n_141), .A2(n_149), .B1(n_1357), .B2(n_1363), .C(n_1365), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_142), .A2(n_205), .B1(n_432), .B2(n_435), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_142), .A2(n_290), .B1(n_507), .B2(n_511), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g1117 ( .A1(n_143), .A2(n_260), .B1(n_836), .B2(n_936), .Y(n_1117) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_143), .A2(n_339), .B1(n_414), .B2(n_714), .C(n_875), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1673 ( .A1(n_144), .A2(n_219), .B1(n_1674), .B2(n_1678), .Y(n_1673) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_145), .A2(n_328), .B1(n_641), .B2(n_645), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_145), .A2(n_328), .B1(n_653), .B2(n_654), .Y(n_652) );
OAI211xp5_ASAP7_75t_SL g929 ( .A1(n_146), .A2(n_930), .B(n_933), .C(n_938), .Y(n_929) );
INVx1_ASAP7_75t_L g957 ( .A(n_146), .Y(n_957) );
AOI221xp5_ASAP7_75t_L g1315 ( .A1(n_147), .A2(n_311), .B1(n_768), .B2(n_1310), .C(n_1316), .Y(n_1315) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_148), .A2(n_224), .B1(n_402), .B2(n_409), .Y(n_401) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_148), .Y(n_493) );
INVx1_ASAP7_75t_L g1380 ( .A(n_149), .Y(n_1380) );
OAI222xp33_ASAP7_75t_L g919 ( .A1(n_150), .A2(n_276), .B1(n_839), .B2(n_843), .C1(n_920), .C2(n_923), .Y(n_919) );
INVx1_ASAP7_75t_L g952 ( .A(n_150), .Y(n_952) );
INVx1_ASAP7_75t_L g1213 ( .A(n_151), .Y(n_1213) );
INVx1_ASAP7_75t_L g1613 ( .A(n_152), .Y(n_1613) );
INVx1_ASAP7_75t_L g1905 ( .A(n_153), .Y(n_1905) );
AOI22xp33_ASAP7_75t_L g1934 ( .A1(n_153), .A2(n_210), .B1(n_1139), .B2(n_1314), .Y(n_1934) );
XNOR2x1_ASAP7_75t_L g915 ( .A(n_154), .B(n_916), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g1689 ( .A1(n_154), .A2(n_230), .B1(n_1681), .B2(n_1684), .Y(n_1689) );
INVx1_ASAP7_75t_L g1284 ( .A(n_155), .Y(n_1284) );
AOI221xp5_ASAP7_75t_SL g1001 ( .A1(n_156), .A2(n_319), .B1(n_1002), .B2(n_1003), .C(n_1004), .Y(n_1001) );
INVx1_ASAP7_75t_L g1032 ( .A(n_156), .Y(n_1032) );
OAI222xp33_ASAP7_75t_L g1468 ( .A1(n_157), .A2(n_249), .B1(n_256), .B2(n_895), .C1(n_903), .C2(n_1343), .Y(n_1468) );
OAI211xp5_ASAP7_75t_L g1470 ( .A1(n_157), .A2(n_930), .B(n_1471), .C(n_1477), .Y(n_1470) );
CKINVDCx5p33_ASAP7_75t_R g999 ( .A(n_158), .Y(n_999) );
INVx1_ASAP7_75t_L g1192 ( .A(n_159), .Y(n_1192) );
INVx1_ASAP7_75t_L g1036 ( .A(n_160), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_161), .A2(n_354), .B1(n_830), .B2(n_831), .C(n_833), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_161), .A2(n_259), .B1(n_875), .B2(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g701 ( .A(n_162), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_162), .A2(n_169), .B1(n_730), .B2(n_732), .Y(n_729) );
INVxp67_ASAP7_75t_SL g1608 ( .A(n_163), .Y(n_1608) );
AOI221xp5_ASAP7_75t_L g1643 ( .A1(n_163), .A2(n_257), .B1(n_802), .B2(n_1004), .C(n_1633), .Y(n_1643) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_164), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g775 ( .A1(n_165), .A2(n_198), .B1(n_441), .B2(n_776), .C(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g812 ( .A(n_165), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_166), .A2(n_349), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g710 ( .A(n_169), .Y(n_710) );
INVx1_ASAP7_75t_L g1494 ( .A(n_170), .Y(n_1494) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_171), .A2(n_290), .B1(n_385), .B2(n_390), .C(n_396), .Y(n_384) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_171), .Y(n_491) );
INVx1_ASAP7_75t_L g1273 ( .A(n_172), .Y(n_1273) );
INVx1_ASAP7_75t_L g1625 ( .A(n_173), .Y(n_1625) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_174), .A2(n_309), .B1(n_438), .B2(n_703), .C(n_705), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g1330 ( .A1(n_175), .A2(n_324), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
INVx1_ASAP7_75t_L g1454 ( .A(n_176), .Y(n_1454) );
OAI221xp5_ASAP7_75t_SL g1482 ( .A1(n_176), .A2(n_182), .B1(n_843), .B2(n_1483), .C(n_1484), .Y(n_1482) );
INVx1_ASAP7_75t_L g628 ( .A(n_177), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_177), .A2(n_589), .B(n_658), .C(n_660), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g1418 ( .A1(n_178), .A2(n_209), .B1(n_1419), .B2(n_1422), .C(n_1423), .Y(n_1418) );
INVx1_ASAP7_75t_L g939 ( .A(n_179), .Y(n_939) );
INVx1_ASAP7_75t_L g1402 ( .A(n_180), .Y(n_1402) );
INVx1_ASAP7_75t_L g1063 ( .A(n_181), .Y(n_1063) );
INVx1_ASAP7_75t_L g1455 ( .A(n_182), .Y(n_1455) );
INVx2_ASAP7_75t_L g1677 ( .A(n_183), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_183), .B(n_305), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_183), .B(n_1683), .Y(n_1685) );
AOI21xp5_ASAP7_75t_L g1414 ( .A1(n_184), .A2(n_875), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1442 ( .A(n_184), .Y(n_1442) );
AOI22xp5_ASAP7_75t_L g1694 ( .A1(n_185), .A2(n_281), .B1(n_1681), .B2(n_1684), .Y(n_1694) );
INVxp67_ASAP7_75t_SL g1912 ( .A(n_186), .Y(n_1912) );
AOI22xp33_ASAP7_75t_SL g1937 ( .A1(n_186), .A2(n_326), .B1(n_1052), .B2(n_1938), .Y(n_1937) );
XNOR2xp5_ASAP7_75t_L g817 ( .A(n_187), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g1509 ( .A(n_188), .Y(n_1509) );
OAI211xp5_ASAP7_75t_L g1347 ( .A1(n_189), .A2(n_457), .B(n_1348), .C(n_1366), .Y(n_1347) );
OAI21xp33_ASAP7_75t_L g1110 ( .A1(n_192), .A2(n_1096), .B(n_1111), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_192), .A2(n_292), .B1(n_879), .B2(n_1144), .C(n_1145), .Y(n_1143) );
AOI22xp5_ASAP7_75t_L g1705 ( .A1(n_193), .A2(n_314), .B1(n_1674), .B2(n_1688), .Y(n_1705) );
INVx1_ASAP7_75t_L g1023 ( .A(n_194), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_195), .A2(n_286), .B1(n_385), .B2(n_390), .C(n_396), .Y(n_784) );
INVx1_ASAP7_75t_L g816 ( .A(n_195), .Y(n_816) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_196), .A2(n_457), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g716 ( .A(n_196), .Y(n_716) );
INVx1_ASAP7_75t_L g569 ( .A(n_197), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_200), .Y(n_1057) );
INVx1_ASAP7_75t_L g1066 ( .A(n_201), .Y(n_1066) );
INVx1_ASAP7_75t_L g746 ( .A(n_202), .Y(n_746) );
INVx1_ASAP7_75t_L g1399 ( .A(n_204), .Y(n_1399) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_205), .A2(n_457), .B(n_471), .C(n_492), .Y(n_456) );
INVx1_ASAP7_75t_L g1391 ( .A(n_207), .Y(n_1391) );
AOI22xp33_ASAP7_75t_SL g1116 ( .A1(n_208), .A2(n_329), .B1(n_723), .B2(n_807), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_208), .A2(n_237), .B1(n_414), .B2(n_705), .C(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1443 ( .A(n_209), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1916 ( .A1(n_210), .A2(n_356), .B1(n_1091), .B2(n_1917), .Y(n_1916) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_211), .A2(n_254), .B1(n_836), .B2(n_936), .Y(n_1514) );
INVx2_ASAP7_75t_L g383 ( .A(n_212), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_212), .B(n_381), .Y(n_405) );
INVx1_ASAP7_75t_L g449 ( .A(n_212), .Y(n_449) );
INVx1_ASAP7_75t_L g899 ( .A(n_213), .Y(n_899) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_214), .A2(n_396), .B(n_690), .C(n_691), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_214), .Y(n_751) );
INVxp67_ASAP7_75t_SL g1177 ( .A(n_215), .Y(n_1177) );
XOR2xp5_ASAP7_75t_L g1038 ( .A(n_216), .B(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1206 ( .A(n_218), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_220), .A2(n_318), .B1(n_445), .B2(n_772), .Y(n_1049) );
INVx1_ASAP7_75t_L g1101 ( .A(n_220), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1707 ( .A1(n_221), .A2(n_317), .B1(n_1681), .B2(n_1684), .Y(n_1707) );
INVx1_ASAP7_75t_L g1033 ( .A(n_222), .Y(n_1033) );
INVx1_ASAP7_75t_L g1559 ( .A(n_223), .Y(n_1559) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_224), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_225), .A2(n_338), .B1(n_936), .B2(n_1123), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_225), .A2(n_260), .B1(n_875), .B2(n_964), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_226), .A2(n_277), .B1(n_440), .B2(n_964), .Y(n_1424) );
INVx1_ASAP7_75t_L g1904 ( .A(n_227), .Y(n_1904) );
AOI22xp33_ASAP7_75t_SL g1935 ( .A1(n_227), .A2(n_356), .B1(n_1314), .B2(n_1936), .Y(n_1935) );
BUFx3_ASAP7_75t_L g375 ( .A(n_228), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_229), .B(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1165 ( .A(n_231), .Y(n_1165) );
INVx1_ASAP7_75t_L g1112 ( .A(n_232), .Y(n_1112) );
OAI221xp5_ASAP7_75t_L g1274 ( .A1(n_233), .A2(n_300), .B1(n_1275), .B2(n_1276), .C(n_1277), .Y(n_1274) );
OAI211xp5_ASAP7_75t_L g1281 ( .A1(n_233), .A2(n_788), .B(n_1282), .C(n_1285), .Y(n_1281) );
OAI21xp5_ASAP7_75t_SL g1921 ( .A1(n_234), .A2(n_1343), .B(n_1922), .Y(n_1921) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_235), .Y(n_1261) );
OAI221xp5_ASAP7_75t_SL g1635 ( .A1(n_236), .A2(n_334), .B1(n_1636), .B2(n_1638), .C(n_1639), .Y(n_1635) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_237), .A2(n_339), .B1(n_721), .B2(n_1126), .Y(n_1125) );
OAI21xp5_ASAP7_75t_L g942 ( .A1(n_238), .A2(n_901), .B(n_943), .Y(n_942) );
OAI211xp5_ASAP7_75t_SL g1538 ( .A1(n_239), .A2(n_658), .B(n_1539), .C(n_1541), .Y(n_1538) );
INVx1_ASAP7_75t_L g1583 ( .A(n_239), .Y(n_1583) );
INVx1_ASAP7_75t_L g880 ( .A(n_240), .Y(n_880) );
INVx1_ASAP7_75t_L g425 ( .A(n_241), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g1700 ( .A1(n_242), .A2(n_266), .B1(n_1674), .B2(n_1678), .Y(n_1700) );
INVx1_ASAP7_75t_L g1544 ( .A(n_243), .Y(n_1544) );
OAI211xp5_ASAP7_75t_SL g1579 ( .A1(n_243), .A2(n_618), .B(n_1580), .C(n_1581), .Y(n_1579) );
CKINVDCx5p33_ASAP7_75t_R g1218 ( .A(n_244), .Y(n_1218) );
INVx1_ASAP7_75t_L g1367 ( .A(n_245), .Y(n_1367) );
INVx1_ASAP7_75t_L g1408 ( .A(n_246), .Y(n_1408) );
INVx1_ASAP7_75t_L g1919 ( .A(n_248), .Y(n_1919) );
INVx1_ASAP7_75t_L g370 ( .A(n_250), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g1053 ( .A1(n_251), .A2(n_273), .B1(n_388), .B2(n_570), .C(n_892), .Y(n_1053) );
INVx1_ASAP7_75t_L g826 ( .A(n_252), .Y(n_826) );
INVx1_ASAP7_75t_L g1302 ( .A(n_253), .Y(n_1302) );
INVx1_ASAP7_75t_L g465 ( .A(n_255), .Y(n_465) );
BUFx3_ASAP7_75t_L g519 ( .A(n_255), .Y(n_519) );
INVx1_ASAP7_75t_L g1616 ( .A(n_257), .Y(n_1616) );
OAI211xp5_ASAP7_75t_L g1913 ( .A1(n_258), .A2(n_930), .B(n_1914), .C(n_1918), .Y(n_1913) );
INVx1_ASAP7_75t_L g1930 ( .A(n_258), .Y(n_1930) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_261), .Y(n_1073) );
INVxp67_ASAP7_75t_SL g1426 ( .A(n_262), .Y(n_1426) );
OAI322xp33_ASAP7_75t_SL g1606 ( .A1(n_263), .A2(n_582), .A3(n_1570), .B1(n_1607), .B2(n_1612), .C1(n_1615), .C2(n_1622), .Y(n_1606) );
OAI22xp33_ASAP7_75t_SL g1644 ( .A1(n_263), .A2(n_268), .B1(n_930), .B2(n_1645), .Y(n_1644) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_264), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_265), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g1299 ( .A(n_267), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g1270 ( .A(n_269), .Y(n_1270) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_270), .A2(n_336), .B1(n_441), .B2(n_768), .C(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g804 ( .A(n_270), .Y(n_804) );
INVx1_ASAP7_75t_L g771 ( .A(n_271), .Y(n_771) );
INVx1_ASAP7_75t_L g1619 ( .A(n_272), .Y(n_1619) );
OA222x2_ASAP7_75t_L g1095 ( .A1(n_273), .A2(n_289), .B1(n_342), .B2(n_753), .C1(n_1096), .C2(n_1098), .Y(n_1095) );
INVx1_ASAP7_75t_L g588 ( .A(n_275), .Y(n_588) );
INVx1_ASAP7_75t_L g955 ( .A(n_276), .Y(n_955) );
AOI32xp33_ASAP7_75t_L g1433 ( .A1(n_277), .A2(n_985), .A3(n_1434), .B1(n_1436), .B2(n_1957), .Y(n_1433) );
XOR2xp5_ASAP7_75t_L g762 ( .A(n_278), .B(n_763), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g1525 ( .A1(n_279), .A2(n_1343), .B(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1167 ( .A(n_280), .Y(n_1167) );
XOR2x2_ASAP7_75t_L g1898 ( .A(n_281), .B(n_1899), .Y(n_1898) );
AOI22xp33_ASAP7_75t_L g1942 ( .A1(n_281), .A2(n_1943), .B1(n_1947), .B2(n_1950), .Y(n_1942) );
OAI22xp5_ASAP7_75t_SL g1596 ( .A1(n_283), .A2(n_1597), .B1(n_1598), .B2(n_1646), .Y(n_1596) );
INVx1_ASAP7_75t_L g1646 ( .A(n_283), .Y(n_1646) );
AOI22xp5_ASAP7_75t_L g1648 ( .A1(n_283), .A2(n_1597), .B1(n_1598), .B2(n_1646), .Y(n_1648) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_285), .A2(n_414), .B(n_416), .C(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g541 ( .A(n_285), .Y(n_541) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_286), .Y(n_792) );
INVx1_ASAP7_75t_L g378 ( .A(n_287), .Y(n_378) );
INVx1_ASAP7_75t_L g395 ( .A(n_287), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g1915 ( .A1(n_288), .A2(n_326), .B1(n_833), .B2(n_985), .C(n_1002), .Y(n_1915) );
INVx1_ASAP7_75t_L g1051 ( .A(n_289), .Y(n_1051) );
INVx1_ASAP7_75t_L g1120 ( .A(n_291), .Y(n_1120) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_292), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g1216 ( .A(n_293), .Y(n_1216) );
INVx1_ASAP7_75t_L g796 ( .A(n_294), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_295), .A2(n_330), .B1(n_432), .B2(n_435), .Y(n_766) );
INVx1_ASAP7_75t_L g794 ( .A(n_295), .Y(n_794) );
INVx1_ASAP7_75t_L g1561 ( .A(n_296), .Y(n_1561) );
INVxp67_ASAP7_75t_SL g1180 ( .A(n_297), .Y(n_1180) );
INVx1_ASAP7_75t_L g578 ( .A(n_298), .Y(n_578) );
INVx1_ASAP7_75t_L g1564 ( .A(n_299), .Y(n_1564) );
INVx1_ASAP7_75t_L g1252 ( .A(n_301), .Y(n_1252) );
INVx1_ASAP7_75t_L g1555 ( .A(n_302), .Y(n_1555) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_303), .Y(n_848) );
INVx1_ASAP7_75t_L g1458 ( .A(n_304), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_305), .B(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1683 ( .A(n_305), .Y(n_1683) );
CKINVDCx5p33_ASAP7_75t_R g1924 ( .A(n_306), .Y(n_1924) );
XNOR2xp5_ASAP7_75t_L g1295 ( .A(n_307), .B(n_1296), .Y(n_1295) );
OAI22xp33_ASAP7_75t_L g1534 ( .A1(n_308), .A2(n_359), .B1(n_1535), .B2(n_1537), .Y(n_1534) );
OAI22xp33_ASAP7_75t_L g1591 ( .A1(n_308), .A2(n_359), .B1(n_643), .B2(n_1592), .Y(n_1591) );
AOI221xp5_ASAP7_75t_SL g736 ( .A1(n_309), .A2(n_310), .B1(n_725), .B2(n_737), .C(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g709 ( .A(n_310), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_313), .A2(n_684), .B1(n_685), .B2(n_757), .Y(n_683) );
INVx1_ASAP7_75t_L g757 ( .A(n_313), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1723 ( .A1(n_313), .A2(n_346), .B1(n_1681), .B2(n_1684), .Y(n_1723) );
INVx1_ASAP7_75t_L g1360 ( .A(n_315), .Y(n_1360) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_315), .A2(n_360), .B1(n_708), .B2(n_1376), .C(n_1377), .Y(n_1375) );
INVx1_ASAP7_75t_L g574 ( .A(n_316), .Y(n_574) );
INVx1_ASAP7_75t_L g1100 ( .A(n_318), .Y(n_1100) );
INVx1_ASAP7_75t_L g1026 ( .A(n_319), .Y(n_1026) );
INVx1_ASAP7_75t_L g921 ( .A(n_320), .Y(n_921) );
INVxp67_ASAP7_75t_SL g1430 ( .A(n_321), .Y(n_1430) );
INVx1_ASAP7_75t_L g419 ( .A(n_322), .Y(n_419) );
INVx1_ASAP7_75t_L g1521 ( .A(n_325), .Y(n_1521) );
INVxp67_ASAP7_75t_SL g1642 ( .A(n_327), .Y(n_1642) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_329), .A2(n_338), .B1(n_964), .B2(n_966), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_330), .Y(n_814) );
INVx1_ASAP7_75t_L g1543 ( .A(n_331), .Y(n_1543) );
INVx1_ASAP7_75t_L g526 ( .A(n_332), .Y(n_526) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_333), .Y(n_468) );
INVxp67_ASAP7_75t_SL g1600 ( .A(n_334), .Y(n_1600) );
CKINVDCx5p33_ASAP7_75t_R g1266 ( .A(n_335), .Y(n_1266) );
INVx1_ASAP7_75t_L g809 ( .A(n_336), .Y(n_809) );
INVx1_ASAP7_75t_L g740 ( .A(n_337), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g1194 ( .A1(n_340), .A2(n_516), .B(n_985), .Y(n_1194) );
INVx1_ASAP7_75t_L g1614 ( .A(n_341), .Y(n_1614) );
INVx1_ASAP7_75t_L g1046 ( .A(n_342), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_343), .Y(n_1214) );
INVx2_ASAP7_75t_L g455 ( .A(n_347), .Y(n_455) );
INVx1_ASAP7_75t_L g462 ( .A(n_347), .Y(n_462) );
INVx1_ASAP7_75t_L g475 ( .A(n_347), .Y(n_475) );
XOR2x2_ASAP7_75t_L g557 ( .A(n_348), .B(n_558), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g1487 ( .A1(n_349), .A2(n_351), .B1(n_852), .B2(n_985), .C(n_1188), .Y(n_1487) );
INVx1_ASAP7_75t_L g780 ( .A(n_350), .Y(n_780) );
INVx1_ASAP7_75t_L g1183 ( .A(n_352), .Y(n_1183) );
INVx1_ASAP7_75t_L g1255 ( .A(n_353), .Y(n_1255) );
INVx1_ASAP7_75t_L g590 ( .A(n_355), .Y(n_590) );
INVx1_ASAP7_75t_L g1611 ( .A(n_357), .Y(n_1611) );
INVx1_ASAP7_75t_L g1557 ( .A(n_358), .Y(n_1557) );
INVx1_ASAP7_75t_L g1352 ( .A(n_360), .Y(n_1352) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_1653), .B(n_1665), .Y(n_361) );
XNOR2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_910), .Y(n_362) );
XOR2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_759), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_554), .B2(n_555), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI211x1_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_450), .B(n_456), .C(n_499), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_412), .Y(n_368) );
AOI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_384), .C(n_401), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g471 ( .A1(n_370), .A2(n_472), .B1(n_479), .B2(n_480), .C1(n_487), .C2(n_491), .Y(n_471) );
INVx2_ASAP7_75t_L g690 ( .A(n_371), .Y(n_690) );
AOI211xp5_ASAP7_75t_SL g781 ( .A1(n_371), .A2(n_782), .B(n_783), .C(n_784), .Y(n_781) );
AOI211xp5_ASAP7_75t_SL g1153 ( .A1(n_371), .A2(n_1154), .B(n_1155), .C(n_1156), .Y(n_1153) );
AOI221xp5_ASAP7_75t_L g1235 ( .A1(n_371), .A2(n_1043), .B1(n_1230), .B2(n_1236), .C(n_1239), .Y(n_1235) );
AOI221xp5_ASAP7_75t_L g1272 ( .A1(n_371), .A2(n_1043), .B1(n_1273), .B2(n_1274), .C(n_1279), .Y(n_1272) );
AOI211xp5_ASAP7_75t_SL g1371 ( .A1(n_371), .A2(n_1367), .B(n_1372), .C(n_1373), .Y(n_1371) );
AOI211xp5_ASAP7_75t_SL g1401 ( .A1(n_371), .A2(n_1402), .B(n_1403), .C(n_1404), .Y(n_1401) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x6_ASAP7_75t_L g903 ( .A(n_372), .B(n_904), .Y(n_903) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_373), .B(n_379), .Y(n_372) );
AND2x2_ASAP7_75t_L g433 ( .A(n_373), .B(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g713 ( .A(n_373), .Y(n_713) );
INVx8_ASAP7_75t_L g769 ( .A(n_373), .Y(n_769) );
BUFx3_ASAP7_75t_L g1244 ( .A(n_373), .Y(n_1244) );
HB1xp67_ASAP7_75t_L g1499 ( .A(n_373), .Y(n_1499) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
AND2x4_ASAP7_75t_L g407 ( .A(n_374), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_375), .Y(n_389) );
AND2x4_ASAP7_75t_L g415 ( .A(n_375), .B(n_394), .Y(n_415) );
OR2x2_ASAP7_75t_L g424 ( .A(n_375), .B(n_377), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_375), .B(n_395), .Y(n_429) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g408 ( .A(n_378), .Y(n_408) );
AND2x6_ASAP7_75t_L g386 ( .A(n_379), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g391 ( .A(n_379), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g400 ( .A(n_379), .Y(n_400) );
AND2x4_ASAP7_75t_L g863 ( .A(n_379), .B(n_474), .Y(n_863) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_380), .B(n_449), .Y(n_448) );
NAND3x1_ASAP7_75t_L g585 ( .A(n_380), .B(n_449), .C(n_586), .Y(n_585) );
OR2x4_ASAP7_75t_L g653 ( .A(n_380), .B(n_424), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_380), .Y(n_656) );
AND2x4_ASAP7_75t_L g659 ( .A(n_380), .B(n_415), .Y(n_659) );
OR2x6_ASAP7_75t_L g674 ( .A(n_380), .B(n_675), .Y(n_674) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
NAND2xp33_ASAP7_75t_SL g563 ( .A(n_381), .B(n_383), .Y(n_563) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_383), .Y(n_679) );
AND3x4_ASAP7_75t_L g960 ( .A(n_383), .B(n_421), .C(n_859), .Y(n_960) );
INVx4_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_386), .A2(n_391), .B1(n_692), .B2(n_693), .Y(n_691) );
AND2x4_ASAP7_75t_SL g888 ( .A(n_387), .B(n_863), .Y(n_888) );
NAND2x1_ASAP7_75t_L g954 ( .A(n_387), .B(n_863), .Y(n_954) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_387), .B(n_863), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_387), .B(n_863), .Y(n_1508) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_389), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g411 ( .A(n_389), .B(n_393), .Y(n_411) );
BUFx2_ASAP7_75t_L g664 ( .A(n_389), .Y(n_664) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g1134 ( .A(n_391), .Y(n_1134) );
INVx1_ASAP7_75t_L g892 ( .A(n_392), .Y(n_892) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g399 ( .A(n_395), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g1135 ( .A(n_396), .Y(n_1135) );
OR2x6_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g1172 ( .A(n_397), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g1265 ( .A1(n_397), .A2(n_447), .B1(n_568), .B2(n_1266), .C(n_1267), .Y(n_1265) );
INVx1_ASAP7_75t_L g1422 ( .A(n_397), .Y(n_1422) );
INVx1_ASAP7_75t_L g1540 ( .A(n_397), .Y(n_1540) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_398), .Y(n_571) );
BUFx2_ASAP7_75t_L g667 ( .A(n_399), .Y(n_667) );
INVx1_ASAP7_75t_L g1054 ( .A(n_400), .Y(n_1054) );
OR2x6_ASAP7_75t_SL g402 ( .A(n_403), .B(n_406), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g410 ( .A(n_404), .B(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_404), .Y(n_1044) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g434 ( .A(n_405), .Y(n_434) );
OR2x2_ASAP7_75t_L g897 ( .A(n_405), .B(n_548), .Y(n_897) );
BUFx2_ASAP7_75t_L g577 ( .A(n_406), .Y(n_577) );
INVx3_ASAP7_75t_L g945 ( .A(n_406), .Y(n_945) );
INVx1_ASAP7_75t_L g1610 ( .A(n_406), .Y(n_1610) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx8_ASAP7_75t_L g418 ( .A(n_407), .Y(n_418) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_407), .Y(n_773) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g441 ( .A(n_411), .Y(n_441) );
BUFx12f_ASAP7_75t_L g964 ( .A(n_411), .Y(n_964) );
INVx5_ASAP7_75t_L g1164 ( .A(n_411), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1314 ( .A(n_411), .Y(n_1314) );
BUFx2_ASAP7_75t_L g1376 ( .A(n_411), .Y(n_1376) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_431), .C(n_437), .Y(n_412) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g436 ( .A(n_415), .B(n_434), .Y(n_436) );
BUFx2_ASAP7_75t_L g704 ( .A(n_415), .Y(n_704) );
BUFx2_ASAP7_75t_L g862 ( .A(n_415), .Y(n_862) );
INVx2_ASAP7_75t_L g883 ( .A(n_415), .Y(n_883) );
BUFx2_ASAP7_75t_L g962 ( .A(n_415), .Y(n_962) );
BUFx2_ASAP7_75t_L g1621 ( .A(n_415), .Y(n_1621) );
BUFx2_ASAP7_75t_L g1938 ( .A(n_415), .Y(n_1938) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B(n_420), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g865 ( .A1(n_417), .A2(n_866), .B(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g966 ( .A(n_417), .Y(n_966) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g777 ( .A(n_418), .Y(n_777) );
AND2x4_ASAP7_75t_L g909 ( .A(n_418), .B(n_908), .Y(n_909) );
INVx3_ASAP7_75t_L g1249 ( .A(n_418), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g1936 ( .A(n_418), .Y(n_1936) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_419), .A2(n_521), .B1(n_525), .B2(n_526), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_420), .A2(n_443), .B1(n_771), .B2(n_772), .C(n_774), .Y(n_770) );
OAI221xp5_ASAP7_75t_L g1072 ( .A1(n_420), .A2(n_877), .B1(n_1073), .B2(n_1074), .C(n_1075), .Y(n_1072) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_420), .A2(n_1164), .B1(n_1165), .B2(n_1166), .C(n_1167), .Y(n_1163) );
OAI221xp5_ASAP7_75t_L g1245 ( .A1(n_420), .A2(n_443), .B1(n_1031), .B2(n_1218), .C(n_1220), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_420), .A2(n_571), .B1(n_1261), .B2(n_1262), .C(n_1263), .Y(n_1260) );
OAI221xp5_ASAP7_75t_L g1382 ( .A1(n_420), .A2(n_777), .B1(n_1361), .B2(n_1379), .C(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1415 ( .A(n_420), .Y(n_1415) );
INVx3_ASAP7_75t_L g663 ( .A(n_421), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_426), .B2(n_430), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_423), .A2(n_447), .B1(n_1063), .B2(n_1064), .C(n_1066), .Y(n_1062) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx3_ASAP7_75t_L g445 ( .A(n_424), .Y(n_445) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_424), .Y(n_568) );
OR2x4_ASAP7_75t_L g672 ( .A(n_424), .B(n_656), .Y(n_672) );
INVx2_ASAP7_75t_L g699 ( .A(n_424), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_425), .A2(n_446), .B1(n_528), .B2(n_533), .Y(n_527) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g575 ( .A(n_427), .Y(n_575) );
CKINVDCx8_ASAP7_75t_R g879 ( .A(n_427), .Y(n_879) );
INVx3_ASAP7_75t_L g1250 ( .A(n_427), .Y(n_1250) );
INVx3_ASAP7_75t_L g1574 ( .A(n_427), .Y(n_1574) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g580 ( .A(n_428), .Y(n_580) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g675 ( .A(n_429), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_430), .A2(n_550), .B1(n_552), .B2(n_553), .Y(n_549) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_433), .A2(n_436), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_439), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g655 ( .A(n_440), .B(n_656), .Y(n_655) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_440), .Y(n_708) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_440), .Y(n_878) );
INVx2_ASAP7_75t_L g1144 ( .A(n_440), .Y(n_1144) );
INVx1_ASAP7_75t_L g1160 ( .A(n_440), .Y(n_1160) );
INVx2_ASAP7_75t_L g1263 ( .A(n_440), .Y(n_1263) );
AOI221xp5_ASAP7_75t_SL g1045 ( .A1(n_441), .A2(n_1046), .B1(n_1047), .B2(n_1048), .C(n_1049), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_445), .B2(n_446), .C(n_447), .Y(n_442) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_443), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_443), .A2(n_447), .B1(n_568), .B2(n_779), .C(n_780), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_443), .A2(n_568), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_443), .A2(n_445), .B1(n_447), .B2(n_1214), .C(n_1221), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_444), .A2(n_538), .B1(n_541), .B2(n_542), .Y(n_537) );
INVx1_ASAP7_75t_L g1421 ( .A(n_445), .Y(n_1421) );
INVx3_ASAP7_75t_L g714 ( .A(n_447), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_447), .B(n_1174), .Y(n_1173) );
OAI221xp5_ASAP7_75t_L g1377 ( .A1(n_447), .A2(n_566), .B1(n_1378), .B2(n_1379), .C(n_1380), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_447), .B(n_1424), .Y(n_1423) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_448), .B(n_454), .Y(n_1037) );
OR2x6_ASAP7_75t_L g1505 ( .A(n_448), .B(n_454), .Y(n_1505) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g764 ( .A1(n_451), .A2(n_765), .B(n_781), .C(n_785), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g1234 ( .A1(n_451), .A2(n_1235), .B(n_1240), .C(n_1251), .Y(n_1234) );
AOI21xp5_ASAP7_75t_L g1320 ( .A1(n_451), .A2(n_1321), .B(n_1342), .Y(n_1320) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI31xp33_ASAP7_75t_SL g687 ( .A1(n_452), .A2(n_688), .A3(n_689), .B(n_694), .Y(n_687) );
INVx1_ASAP7_75t_L g941 ( .A(n_452), .Y(n_941) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI21xp5_ASAP7_75t_SL g979 ( .A1(n_453), .A2(n_980), .B(n_1000), .Y(n_979) );
INVx1_ASAP7_75t_L g1077 ( .A(n_453), .Y(n_1077) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g517 ( .A(n_454), .B(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_455), .B(n_478), .Y(n_505) );
INVx2_ASAP7_75t_L g859 ( .A(n_455), .Y(n_859) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_458), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_458), .A2(n_494), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_458), .B(n_1108), .Y(n_1107) );
AOI211xp5_ASAP7_75t_L g1179 ( .A1(n_458), .A2(n_1180), .B(n_1181), .C(n_1185), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_458), .B(n_1233), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_458), .B(n_1278), .Y(n_1280) );
AO211x2_ASAP7_75t_L g1398 ( .A1(n_458), .A2(n_1399), .B(n_1400), .C(n_1427), .Y(n_1398) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .Y(n_458) );
AND2x4_ASAP7_75t_L g494 ( .A(n_459), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g511 ( .A(n_460), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g650 ( .A(n_460), .Y(n_650) );
OR2x2_ASAP7_75t_L g756 ( .A(n_460), .B(n_512), .Y(n_756) );
INVxp67_ASAP7_75t_L g904 ( .A(n_460), .Y(n_904) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g548 ( .A(n_461), .Y(n_548) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_463), .Y(n_825) );
INVx1_ASAP7_75t_L g1479 ( .A(n_463), .Y(n_1479) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_464), .B(n_475), .Y(n_482) );
AND2x2_ASAP7_75t_L g495 ( .A(n_464), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g822 ( .A(n_464), .B(n_483), .Y(n_822) );
AND2x4_ASAP7_75t_L g827 ( .A(n_464), .B(n_496), .Y(n_827) );
AND2x4_ASAP7_75t_SL g842 ( .A(n_464), .B(n_622), .Y(n_842) );
AND2x4_ASAP7_75t_L g931 ( .A(n_464), .B(n_932), .Y(n_931) );
BUFx2_ASAP7_75t_L g987 ( .A(n_464), .Y(n_987) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_465), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_466), .B(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g731 ( .A(n_466), .Y(n_731) );
BUFx6f_ASAP7_75t_L g937 ( .A(n_466), .Y(n_937) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
OR2x2_ASAP7_75t_L g524 ( .A(n_467), .B(n_470), .Y(n_524) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g486 ( .A(n_468), .Y(n_486) );
NAND2x1_ASAP7_75t_L g490 ( .A(n_468), .B(n_470), .Y(n_490) );
AND2x2_ASAP7_75t_L g497 ( .A(n_468), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g514 ( .A(n_468), .Y(n_514) );
OR2x2_ASAP7_75t_L g532 ( .A(n_468), .B(n_470), .Y(n_532) );
AND2x2_ASAP7_75t_L g623 ( .A(n_468), .B(n_470), .Y(n_623) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g485 ( .A(n_470), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g498 ( .A(n_470), .Y(n_498) );
BUFx2_ASAP7_75t_L g510 ( .A(n_470), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_470), .B(n_486), .Y(n_536) );
AOI322xp5_ASAP7_75t_L g719 ( .A1(n_472), .A2(n_720), .A3(n_728), .B1(n_729), .B2(n_735), .C1(n_736), .C2(n_742), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g795 ( .A1(n_472), .A2(n_517), .B1(n_728), .B2(n_796), .C1(n_797), .C2(n_806), .Y(n_795) );
AOI322xp5_ASAP7_75t_L g1186 ( .A1(n_472), .A2(n_728), .A3(n_1187), .B1(n_1189), .B2(n_1194), .C1(n_1195), .C2(n_1196), .Y(n_1186) );
AOI222xp33_ASAP7_75t_L g1228 ( .A1(n_472), .A2(n_480), .B1(n_487), .B2(n_1229), .C1(n_1230), .C2(n_1231), .Y(n_1228) );
AOI222xp33_ASAP7_75t_L g1366 ( .A1(n_472), .A2(n_480), .B1(n_487), .B2(n_1367), .C1(n_1368), .C2(n_1369), .Y(n_1366) );
AOI21xp33_ASAP7_75t_L g1446 ( .A1(n_472), .A2(n_500), .B(n_1447), .Y(n_1446) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
AOI332xp33_ASAP7_75t_L g1282 ( .A1(n_473), .A2(n_476), .A3(n_481), .B1(n_483), .B2(n_487), .B3(n_1273), .C1(n_1283), .C2(n_1284), .Y(n_1282) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g898 ( .A(n_474), .B(n_477), .Y(n_898) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g586 ( .A(n_475), .Y(n_586) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_478), .B(n_513), .Y(n_512) );
AND2x6_ASAP7_75t_L g837 ( .A(n_478), .B(n_622), .Y(n_837) );
INVx1_ASAP7_75t_L g846 ( .A(n_478), .Y(n_846) );
AND2x2_ASAP7_75t_L g995 ( .A(n_478), .B(n_996), .Y(n_995) );
AOI211xp5_ASAP7_75t_L g750 ( .A1(n_480), .A2(n_751), .B(n_752), .C(n_754), .Y(n_750) );
AOI222xp33_ASAP7_75t_L g790 ( .A1(n_480), .A2(n_782), .B1(n_791), .B2(n_792), .C1(n_793), .C2(n_794), .Y(n_790) );
INVx1_ASAP7_75t_L g1098 ( .A(n_480), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_480), .A2(n_487), .B1(n_1112), .B2(n_1113), .Y(n_1111) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g488 ( .A(n_482), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g753 ( .A(n_482), .B(n_489), .Y(n_753) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g856 ( .A(n_484), .Y(n_856) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g734 ( .A(n_485), .Y(n_734) );
BUFx3_ASAP7_75t_L g836 ( .A(n_485), .Y(n_836) );
BUFx6f_ASAP7_75t_L g932 ( .A(n_485), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_487), .A2(n_500), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx3_ASAP7_75t_L g1082 ( .A(n_489), .Y(n_1082) );
INVx2_ASAP7_75t_SL g1563 ( .A(n_489), .Y(n_1563) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g748 ( .A(n_494), .Y(n_748) );
INVx1_ASAP7_75t_L g788 ( .A(n_494), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_494), .B(n_1177), .Y(n_1176) );
NAND2xp33_ASAP7_75t_SL g1251 ( .A(n_494), .B(n_1252), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1390 ( .A(n_494), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_494), .B(n_1426), .Y(n_1425) );
INVx2_ASAP7_75t_L g832 ( .A(n_496), .Y(n_832) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_496), .Y(n_851) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g646 ( .A(n_497), .B(n_636), .Y(n_646) );
INVx2_ASAP7_75t_L g724 ( .A(n_497), .Y(n_724) );
BUFx3_ASAP7_75t_L g802 ( .A(n_497), .Y(n_802) );
OR3x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .C(n_515), .Y(n_499) );
AOI31xp33_ASAP7_75t_L g1115 ( .A1(n_500), .A2(n_517), .A3(n_1116), .B(n_1117), .Y(n_1115) );
NOR3xp33_ASAP7_75t_L g1285 ( .A(n_500), .B(n_1286), .C(n_1293), .Y(n_1285) );
NOR3xp33_ASAP7_75t_L g1348 ( .A(n_500), .B(n_1349), .C(n_1350), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g1083 ( .A1(n_501), .A2(n_1084), .B(n_1085), .Y(n_1083) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_502), .Y(n_525) );
INVx4_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_502), .Y(n_606) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_502), .Y(n_617) );
BUFx4f_ASAP7_75t_L g849 ( .A(n_502), .Y(n_849) );
BUFx4f_ASAP7_75t_L g1288 ( .A(n_502), .Y(n_1288) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2x2_ASAP7_75t_L g507 ( .A(n_504), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_507), .Y(n_755) );
INVx1_ASAP7_75t_L g791 ( .A(n_507), .Y(n_791) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_507), .Y(n_1094) );
INVx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g626 ( .A(n_510), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g845 ( .A(n_510), .Y(n_845) );
BUFx2_ASAP7_75t_L g996 ( .A(n_510), .Y(n_996) );
INVx2_ASAP7_75t_SL g793 ( .A(n_511), .Y(n_793) );
AND2x4_ASAP7_75t_L g901 ( .A(n_511), .B(n_902), .Y(n_901) );
AND2x4_ASAP7_75t_L g1343 ( .A(n_511), .B(n_902), .Y(n_1343) );
INVx1_ASAP7_75t_L g998 ( .A(n_512), .Y(n_998) );
AND2x4_ASAP7_75t_L g631 ( .A(n_513), .B(n_519), .Y(n_631) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI33xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_520), .A3(n_527), .B1(n_537), .B2(n_544), .B3(n_549), .Y(n_515) );
OAI33xp33_ASAP7_75t_L g591 ( .A1(n_516), .A2(n_592), .A3(n_598), .B1(n_602), .B2(n_607), .B3(n_612), .Y(n_591) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g744 ( .A(n_517), .Y(n_744) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_517), .Y(n_1079) );
INVx2_ASAP7_75t_L g1211 ( .A(n_517), .Y(n_1211) );
INVx4_ASAP7_75t_L g1365 ( .A(n_517), .Y(n_1365) );
AND2x4_ASAP7_75t_L g546 ( .A(n_519), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g621 ( .A(n_519), .Y(n_621) );
BUFx2_ASAP7_75t_L g627 ( .A(n_519), .Y(n_627) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g1217 ( .A(n_522), .Y(n_1217) );
INVx2_ASAP7_75t_L g1558 ( .A(n_522), .Y(n_1558) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g540 ( .A(n_524), .Y(n_540) );
BUFx3_ASAP7_75t_L g605 ( .A(n_524), .Y(n_605) );
INVx1_ASAP7_75t_L g1087 ( .A(n_524), .Y(n_1087) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g739 ( .A(n_529), .Y(n_739) );
INVx2_ASAP7_75t_L g925 ( .A(n_529), .Y(n_925) );
INVx2_ASAP7_75t_SL g1566 ( .A(n_529), .Y(n_1566) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g805 ( .A(n_530), .Y(n_805) );
INVx3_ASAP7_75t_L g982 ( .A(n_530), .Y(n_982) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g551 ( .A(n_531), .Y(n_551) );
INVx2_ASAP7_75t_L g635 ( .A(n_531), .Y(n_635) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_533), .A2(n_550), .B1(n_1165), .B2(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g552 ( .A(n_534), .Y(n_552) );
INVx4_ASAP7_75t_L g597 ( .A(n_534), .Y(n_597) );
INVx1_ASAP7_75t_L g928 ( .A(n_534), .Y(n_928) );
BUFx6f_ASAP7_75t_L g1089 ( .A(n_534), .Y(n_1089) );
INVx2_ASAP7_75t_L g1364 ( .A(n_534), .Y(n_1364) );
INVx8_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g639 ( .A(n_535), .B(n_627), .Y(n_639) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_538), .A2(n_1082), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g599 ( .A(n_540), .Y(n_599) );
INVx2_ASAP7_75t_L g1291 ( .A(n_540), .Y(n_1291) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g601 ( .A(n_543), .Y(n_601) );
INVx2_ASAP7_75t_L g1356 ( .A(n_543), .Y(n_1356) );
OAI33xp33_ASAP7_75t_L g1210 ( .A1(n_544), .A2(n_1211), .A3(n_1212), .B1(n_1215), .B2(n_1219), .B3(n_1222), .Y(n_1210) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_546), .B(n_548), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_546), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g728 ( .A(n_546), .B(n_610), .Y(n_728) );
INVx4_ASAP7_75t_L g833 ( .A(n_546), .Y(n_833) );
INVx4_ASAP7_75t_L g1329 ( .A(n_546), .Y(n_1329) );
INVx1_ASAP7_75t_L g649 ( .A(n_547), .Y(n_649) );
AND2x4_ASAP7_75t_L g853 ( .A(n_547), .B(n_621), .Y(n_853) );
OR2x2_ASAP7_75t_L g562 ( .A(n_548), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g611 ( .A(n_548), .Y(n_611) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_548), .Y(n_681) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
BUFx6f_ASAP7_75t_L g1358 ( .A(n_551), .Y(n_1358) );
INVx2_ASAP7_75t_SL g1631 ( .A(n_551), .Y(n_1631) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_552), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_552), .A2(n_809), .B1(n_810), .B2(n_812), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_552), .A2(n_1191), .B1(n_1213), .B2(n_1214), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_552), .A2(n_1223), .B1(n_1225), .B2(n_1226), .Y(n_1222) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_682), .B2(n_758), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_615), .C(n_651), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_591), .Y(n_559) );
OAI33xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .A3(n_572), .B1(n_576), .B2(n_582), .B3(n_587), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx8_ASAP7_75t_L g868 ( .A(n_562), .Y(n_868) );
BUFx4f_ASAP7_75t_L g1021 ( .A(n_562), .Y(n_1021) );
BUFx2_ASAP7_75t_L g705 ( .A(n_563), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_569), .B2(n_570), .Y(n_564) );
OAI22xp5_ASAP7_75t_SL g592 ( .A1(n_565), .A2(n_588), .B1(n_593), .B2(n_596), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_566), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_587) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_568), .A2(n_570), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_569), .A2(n_590), .B1(n_603), .B2(n_606), .Y(n_602) );
HB1xp67_ASAP7_75t_L g1572 ( .A(n_570), .Y(n_1572) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g902 ( .A(n_571), .B(n_897), .Y(n_902) );
INVx4_ASAP7_75t_L g1065 ( .A(n_571), .Y(n_1065) );
INVx3_ASAP7_75t_L g1238 ( .A(n_571), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_571), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_573), .A2(n_578), .B1(n_599), .B2(n_600), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_574), .A2(n_581), .B1(n_593), .B2(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_575), .A2(n_1269), .B1(n_1270), .B2(n_1271), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_579), .B2(n_581), .Y(n_576) );
INVx2_ASAP7_75t_L g1309 ( .A(n_577), .Y(n_1309) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_579), .A2(n_696), .B1(n_700), .B2(n_701), .C(n_702), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_579), .A2(n_707), .B1(n_709), .B2(n_710), .C(n_711), .Y(n_706) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g896 ( .A(n_580), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI33xp33_ASAP7_75t_L g1932 ( .A1(n_583), .A2(n_1317), .A3(n_1933), .B1(n_1934), .B2(n_1935), .B3(n_1937), .Y(n_1932) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g968 ( .A(n_584), .Y(n_968) );
BUFx2_ASAP7_75t_L g1312 ( .A(n_584), .Y(n_1312) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g885 ( .A(n_585), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g1612 ( .A1(n_589), .A2(n_1420), .B1(n_1613), .B2(n_1614), .Y(n_1612) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_595), .A2(n_1057), .B1(n_1068), .B2(n_1082), .Y(n_1081) );
OAI211xp5_ASAP7_75t_L g1351 ( .A1(n_596), .A2(n_1352), .B(n_1353), .C(n_1354), .Y(n_1351) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g614 ( .A(n_597), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_597), .A2(n_780), .B1(n_804), .B2(n_805), .Y(n_803) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_601), .A2(n_1216), .B1(n_1217), .B2(n_1218), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g920 ( .A1(n_603), .A2(n_849), .B1(n_853), .B2(n_921), .C(n_922), .Y(n_920) );
OAI221xp5_ASAP7_75t_L g1359 ( .A1(n_603), .A2(n_1288), .B1(n_1360), .B2(n_1361), .C(n_1362), .Y(n_1359) );
INVx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g1287 ( .A1(n_605), .A2(n_1262), .B1(n_1270), .B2(n_1288), .C(n_1289), .Y(n_1287) );
OAI33xp33_ASAP7_75t_L g1550 ( .A1(n_607), .A2(n_743), .A3(n_1551), .B1(n_1556), .B2(n_1560), .B3(n_1565), .Y(n_1550) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22xp5_ASAP7_75t_SL g1286 ( .A1(n_609), .A2(n_1211), .B1(n_1287), .B2(n_1290), .Y(n_1286) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g1629 ( .A1(n_613), .A2(n_1611), .B1(n_1619), .B2(n_1630), .C(n_1632), .Y(n_1629) );
OAI221xp5_ASAP7_75t_L g1639 ( .A1(n_613), .A2(n_1613), .B1(n_1640), .B2(n_1642), .C(n_1643), .Y(n_1639) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI31xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_632), .A3(n_640), .B(n_647), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g1290 ( .A1(n_617), .A2(n_1261), .B1(n_1266), .B2(n_1291), .C(n_1292), .Y(n_1290) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_617), .A2(n_1557), .B1(n_1558), .B2(n_1559), .Y(n_1556) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g644 ( .A(n_621), .Y(n_644) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_622), .Y(n_727) );
INVx1_ASAP7_75t_L g799 ( .A(n_622), .Y(n_799) );
BUFx3_ASAP7_75t_L g807 ( .A(n_622), .Y(n_807) );
BUFx3_ASAP7_75t_L g830 ( .A(n_622), .Y(n_830) );
BUFx3_ASAP7_75t_L g985 ( .A(n_622), .Y(n_985) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_622), .Y(n_1003) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g1128 ( .A(n_623), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_628), .B2(n_629), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_625), .A2(n_661), .B1(n_665), .B2(n_668), .Y(n_660) );
BUFx3_ASAP7_75t_L g1582 ( .A(n_626), .Y(n_1582) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g1585 ( .A(n_631), .Y(n_1585) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g1588 ( .A(n_634), .Y(n_1588) );
OR2x6_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OR2x6_ASAP7_75t_L g643 ( .A(n_635), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g811 ( .A(n_635), .Y(n_811) );
BUFx4f_ASAP7_75t_L g1191 ( .A(n_635), .Y(n_1191) );
INVxp67_ASAP7_75t_L g1224 ( .A(n_635), .Y(n_1224) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g1590 ( .A(n_639), .Y(n_1590) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_642), .B(n_1664), .Y(n_1663) );
AND2x4_ASAP7_75t_SL g1940 ( .A(n_642), .B(n_1941), .Y(n_1940) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx3_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
CKINVDCx16_ASAP7_75t_R g1592 ( .A(n_646), .Y(n_1592) );
OAI31xp33_ASAP7_75t_L g1578 ( .A1(n_647), .A2(n_1579), .A3(n_1586), .B(n_1591), .Y(n_1578) );
BUFx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g1664 ( .A(n_649), .Y(n_1664) );
NOR2xp33_ASAP7_75t_L g1941 ( .A(n_649), .B(n_1656), .Y(n_1941) );
OAI31xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_657), .A3(n_669), .B(n_676), .Y(n_651) );
INVx2_ASAP7_75t_SL g1536 ( .A(n_653), .Y(n_1536) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g1537 ( .A(n_655), .Y(n_1537) );
CKINVDCx8_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
BUFx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx3_ASAP7_75t_L g1542 ( .A(n_662), .Y(n_1542) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x4_ASAP7_75t_L g666 ( .A(n_663), .B(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_665), .A2(n_1542), .B1(n_1543), .B2(n_1544), .Y(n_1541) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g1546 ( .A(n_672), .Y(n_1546) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g1548 ( .A(n_674), .Y(n_1548) );
INVx1_ASAP7_75t_L g873 ( .A(n_675), .Y(n_873) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_675), .Y(n_1061) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_678), .B(n_680), .Y(n_677) );
AND2x4_ASAP7_75t_L g1532 ( .A(n_678), .B(n_680), .Y(n_1532) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_683), .Y(n_758) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_718), .Y(n_685) );
INVx1_ASAP7_75t_L g1146 ( .A(n_690), .Y(n_1146) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_706), .C(n_715), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g1577 ( .A1(n_698), .A2(n_1237), .B1(n_1555), .B2(n_1564), .Y(n_1577) );
OR2x2_ASAP7_75t_L g1622 ( .A(n_698), .B(n_1623), .Y(n_1622) );
INVx2_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g1070 ( .A(n_699), .Y(n_1070) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_700), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_738) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g1409 ( .A(n_708), .Y(n_1409) );
BUFx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g1166 ( .A(n_713), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_713), .B(n_1278), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_745), .Y(n_718) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g1002 ( .A(n_722), .Y(n_1002) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_723), .Y(n_737) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g1517 ( .A(n_724), .Y(n_1517) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_727), .Y(n_1197) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_728), .Y(n_1084) );
NAND3xp33_ASAP7_75t_L g1121 ( .A(n_728), .B(n_1122), .C(n_1125), .Y(n_1121) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_SL g835 ( .A(n_731), .Y(n_835) );
INVx1_ASAP7_75t_L g855 ( .A(n_731), .Y(n_855) );
INVx2_ASAP7_75t_L g1091 ( .A(n_731), .Y(n_1091) );
INVx2_ASAP7_75t_L g1331 ( .A(n_731), .Y(n_1331) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_734), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
BUFx3_ASAP7_75t_L g1332 ( .A(n_734), .Y(n_1332) );
HB1xp67_ASAP7_75t_L g1917 ( .A(n_734), .Y(n_1917) );
OAI221xp5_ASAP7_75t_L g1484 ( .A1(n_739), .A2(n_1088), .B1(n_1485), .B2(n_1486), .C(n_1487), .Y(n_1484) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
XNOR2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_817), .Y(n_761) );
OR2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_789), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .C(n_775), .Y(n_765) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx8_ASAP7_75t_L g875 ( .A(n_769), .Y(n_875) );
INVx2_ASAP7_75t_L g907 ( .A(n_769), .Y(n_907) );
INVx3_ASAP7_75t_L g1052 ( .A(n_769), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1573 ( .A1(n_772), .A2(n_1557), .B1(n_1567), .B2(n_1574), .Y(n_1573) );
INVx2_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
INVx5_ASAP7_75t_L g1027 ( .A(n_773), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_773), .Y(n_1059) );
INVx3_ASAP7_75t_L g1269 ( .A(n_773), .Y(n_1269) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g1129 ( .A1(n_787), .A2(n_859), .B1(n_1130), .B2(n_1147), .Y(n_1129) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND4xp25_ASAP7_75t_L g789 ( .A(n_790), .B(n_795), .C(n_813), .D(n_815), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g1118 ( .A1(n_791), .A2(n_793), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_791), .A2(n_793), .B1(n_1183), .B2(n_1184), .Y(n_1182) );
AOI222xp33_ASAP7_75t_L g1428 ( .A1(n_791), .A2(n_793), .B1(n_1402), .B2(n_1429), .C1(n_1430), .C2(n_1431), .Y(n_1428) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1633 ( .A(n_799), .Y(n_1633) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_802), .Y(n_1198) );
INVx1_ASAP7_75t_L g1554 ( .A(n_810), .Y(n_1554) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND4x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_860), .C(n_893), .D(n_905), .Y(n_818) );
OAI21xp33_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_838), .B(n_857), .Y(n_819) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_824), .A2(n_826), .B1(n_906), .B2(n_909), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_825), .A2(n_827), .B1(n_939), .B2(n_940), .Y(n_938) );
HB1xp67_ASAP7_75t_L g1324 ( .A(n_825), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_825), .A2(n_827), .B1(n_1521), .B2(n_1522), .Y(n_1520) );
INVx1_ASAP7_75t_L g1645 ( .A(n_825), .Y(n_1645) );
AOI22xp33_ASAP7_75t_L g1918 ( .A1(n_825), .A2(n_1326), .B1(n_1919), .B2(n_1920), .Y(n_1918) );
BUFx6f_ASAP7_75t_L g1326 ( .A(n_827), .Y(n_1326) );
INVx1_ASAP7_75t_L g1481 ( .A(n_827), .Y(n_1481) );
HB1xp67_ASAP7_75t_L g1637 ( .A(n_827), .Y(n_1637) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_834), .B(n_837), .Y(n_828) );
INVx1_ASAP7_75t_L g1338 ( .A(n_831), .Y(n_1338) );
HB1xp67_ASAP7_75t_L g1440 ( .A(n_831), .Y(n_1440) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_837), .A2(n_934), .B(n_935), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_837), .A2(n_931), .B1(n_1298), .B2(n_1328), .C(n_1330), .Y(n_1327) );
AOI21xp5_ASAP7_75t_SL g1471 ( .A1(n_837), .A2(n_1472), .B(n_1476), .Y(n_1471) );
AOI221xp5_ASAP7_75t_L g1515 ( .A1(n_837), .A2(n_931), .B1(n_1494), .B2(n_1516), .C(n_1518), .Y(n_1515) );
INVx1_ASAP7_75t_L g1634 ( .A(n_837), .Y(n_1634) );
AOI21xp5_ASAP7_75t_L g1914 ( .A1(n_837), .A2(n_1915), .B(n_1916), .Y(n_1914) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g1483 ( .A(n_840), .Y(n_1483) );
INVx2_ASAP7_75t_L g1902 ( .A(n_840), .Y(n_1902) );
INVx4_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_842), .Y(n_1334) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g1638 ( .A(n_844), .Y(n_1638) );
NOR2x1_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g993 ( .A(n_846), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B(n_850), .C(n_854), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_848), .A2(n_877), .B1(n_879), .B2(n_880), .C(n_881), .Y(n_876) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_851), .Y(n_1188) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx3_ASAP7_75t_L g1004 ( .A(n_853), .Y(n_1004) );
INVx1_ASAP7_75t_L g1339 ( .A(n_853), .Y(n_1339) );
INVx2_ASAP7_75t_L g1907 ( .A(n_853), .Y(n_1907) );
A2O1A1Ixp33_ASAP7_75t_L g1257 ( .A1(n_857), .A2(n_1258), .B(n_1272), .C(n_1280), .Y(n_1257) );
A2O1A1Ixp33_ASAP7_75t_SL g1400 ( .A1(n_857), .A2(n_1401), .B(n_1405), .C(n_1425), .Y(n_1400) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx2_ASAP7_75t_L g1387 ( .A(n_858), .Y(n_1387) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_SL g1175 ( .A(n_859), .Y(n_1175) );
NOR3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .C(n_886), .Y(n_860) );
INVx3_ASAP7_75t_L g969 ( .A(n_861), .Y(n_969) );
INVx3_ASAP7_75t_L g1306 ( .A(n_861), .Y(n_1306) );
NOR3xp33_ASAP7_75t_L g1451 ( .A(n_861), .B(n_1452), .C(n_1468), .Y(n_1451) );
AND2x4_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_862), .A2(n_1052), .B1(n_1108), .B2(n_1120), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1467 ( .A(n_862), .Y(n_1467) );
AND2x4_ASAP7_75t_SL g890 ( .A(n_863), .B(n_891), .Y(n_890) );
A2O1A1Ixp33_ASAP7_75t_L g1018 ( .A1(n_863), .A2(n_875), .B(n_984), .C(n_1019), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_863), .B(n_891), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_869), .B1(n_876), .B2(n_884), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_868), .Y(n_867) );
OAI21xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B(n_874), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_871), .A2(n_1068), .B1(n_1069), .B2(n_1071), .Y(n_1067) );
INVx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g1028 ( .A(n_873), .Y(n_1028) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g1047 ( .A(n_883), .Y(n_1047) );
INVx2_ASAP7_75t_L g1310 ( .A(n_883), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_885), .Y(n_884) );
AOI33xp33_ASAP7_75t_L g1459 ( .A1(n_885), .A2(n_1317), .A3(n_1460), .B1(n_1461), .B2(n_1463), .B3(n_1466), .Y(n_1459) );
INVx2_ASAP7_75t_L g1576 ( .A(n_885), .Y(n_1576) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g951 ( .A1(n_890), .A2(n_952), .B1(n_953), .B2(n_955), .Y(n_951) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_899), .B(n_900), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_894), .B(n_949), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g1297 ( .A1(n_894), .A2(n_958), .B1(n_1298), .B2(n_1299), .C(n_1300), .Y(n_1297) );
AOI221xp5_ASAP7_75t_L g1493 ( .A1(n_894), .A2(n_958), .B1(n_1494), .B2(n_1495), .C(n_1496), .Y(n_1493) );
AOI21xp5_ASAP7_75t_L g1624 ( .A1(n_894), .A2(n_1625), .B(n_1626), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1923 ( .A(n_894), .B(n_1924), .Y(n_1923) );
INVx8_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AND2x4_ASAP7_75t_L g895 ( .A(n_896), .B(n_898), .Y(n_895) );
INVx1_ASAP7_75t_L g908 ( .A(n_897), .Y(n_908) );
INVx1_ASAP7_75t_L g946 ( .A(n_897), .Y(n_946) );
INVx1_ASAP7_75t_L g1097 ( .A(n_898), .Y(n_1097) );
INVx2_ASAP7_75t_L g1015 ( .A(n_902), .Y(n_1015) );
INVx3_ASAP7_75t_L g958 ( .A(n_903), .Y(n_958) );
INVx5_ASAP7_75t_L g1931 ( .A(n_903), .Y(n_1931) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_906), .A2(n_939), .B1(n_940), .B2(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_906), .A2(n_944), .B1(n_1521), .B2(n_1522), .Y(n_1526) );
AND2x4_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_907), .B(n_908), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_909), .A2(n_1012), .B1(n_1323), .B2(n_1325), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_909), .A2(n_1012), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
INVx2_ASAP7_75t_L g1602 ( .A(n_909), .Y(n_1602) );
AOI22xp33_ASAP7_75t_L g1922 ( .A1(n_909), .A2(n_1012), .B1(n_1919), .B2(n_1920), .Y(n_1922) );
AOI22x1_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_1394), .B1(n_1651), .B2(n_1652), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
AO22x2_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_970), .B2(n_971), .Y(n_912) );
AO22x1_ASAP7_75t_L g1652 ( .A1(n_913), .A2(n_914), .B1(n_970), .B2(n_971), .Y(n_1652) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NOR2x1p5_ASAP7_75t_L g916 ( .A(n_917), .B(n_947), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_SL g918 ( .A1(n_919), .A2(n_929), .B(n_941), .C(n_942), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_925), .B1(n_926), .B2(n_927), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g1565 ( .A1(n_927), .A2(n_1566), .B1(n_1567), .B2(n_1568), .Y(n_1565) );
BUFx3_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx3_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_932), .Y(n_1008) );
INVx1_ASAP7_75t_L g1124 ( .A(n_932), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx3_ASAP7_75t_L g991 ( .A(n_937), .Y(n_991) );
OAI31xp33_ASAP7_75t_L g1627 ( .A1(n_941), .A2(n_1628), .A3(n_1635), .B(n_1644), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_944), .A2(n_999), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
INVx2_ASAP7_75t_L g1031 ( .A(n_945), .Y(n_1031) );
INVx2_ASAP7_75t_L g1275 ( .A(n_945), .Y(n_1275) );
INVxp67_ASAP7_75t_L g1623 ( .A(n_946), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_950), .Y(n_947) );
AND4x1_ASAP7_75t_L g950 ( .A(n_951), .B(n_956), .C(n_959), .D(n_969), .Y(n_950) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .Y(n_956) );
AOI33xp33_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .A3(n_963), .B1(n_965), .B2(n_967), .B3(n_968), .Y(n_959) );
BUFx3_ASAP7_75t_L g1317 ( .A(n_960), .Y(n_1317) );
AOI33xp33_ASAP7_75t_L g1497 ( .A1(n_960), .A2(n_1498), .A3(n_1500), .B1(n_1502), .B2(n_1503), .B3(n_1504), .Y(n_1497) );
BUFx2_ASAP7_75t_L g1319 ( .A(n_964), .Y(n_1319) );
NAND3xp33_ASAP7_75t_L g1496 ( .A(n_969), .B(n_1497), .C(n_1506), .Y(n_1496) );
AND4x1_ASAP7_75t_SL g1925 ( .A(n_969), .B(n_1926), .C(n_1929), .D(n_1932), .Y(n_1925) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
XOR2x2_ASAP7_75t_L g971 ( .A(n_972), .B(n_1202), .Y(n_971) );
XNOR2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_1102), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_1038), .Y(n_974) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
OR2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_1009), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_987), .B(n_988), .Y(n_980) );
INVx2_ASAP7_75t_SL g1641 ( .A(n_982), .Y(n_1641) );
A2O1A1Ixp33_ASAP7_75t_L g989 ( .A1(n_985), .A2(n_990), .B(n_992), .C(n_993), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_994), .Y(n_988) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g1519 ( .A(n_991), .Y(n_1519) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_997), .B1(n_998), .B2(n_999), .Y(n_994) );
INVx1_ASAP7_75t_L g1341 ( .A(n_995), .Y(n_1341) );
AOI222xp33_ASAP7_75t_L g1512 ( .A1(n_995), .A2(n_1334), .B1(n_1507), .B2(n_1509), .C1(n_1513), .C2(n_1514), .Y(n_1512) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1005), .B1(n_1006), .B2(n_1007), .Y(n_1000) );
NAND3xp33_ASAP7_75t_SL g1009 ( .A(n_1010), .B(n_1013), .C(n_1016), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
NOR2xp33_ASAP7_75t_SL g1016 ( .A(n_1017), .B(n_1020), .Y(n_1016) );
OAI33xp33_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1022), .A3(n_1025), .B1(n_1030), .B2(n_1034), .B3(n_1037), .Y(n_1020) );
BUFx3_ASAP7_75t_L g1570 ( .A(n_1021), .Y(n_1570) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .B1(n_1028), .B2(n_1029), .Y(n_1025) );
INVx8_ASAP7_75t_L g1139 ( .A(n_1027), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_1028), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1575 ( .A1(n_1031), .A2(n_1061), .B1(n_1559), .B2(n_1568), .Y(n_1575) );
NAND4xp75_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1078), .C(n_1095), .D(n_1099), .Y(n_1039) );
OAI21x1_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1055), .B(n_1076), .Y(n_1040) );
OAI21xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1045), .B(n_1050), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1043), .A2(n_1112), .B1(n_1143), .B2(n_1146), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
A2O1A1Ixp33_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1052), .B(n_1053), .C(n_1054), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1062), .B1(n_1067), .B2(n_1072), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1060), .B2(n_1061), .Y(n_1056) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_1060), .A2(n_1073), .B1(n_1086), .B2(n_1088), .C(n_1090), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1607 ( .A1(n_1061), .A2(n_1608), .B1(n_1609), .B2(n_1611), .Y(n_1607) );
OAI221xp5_ASAP7_75t_L g1615 ( .A1(n_1061), .A2(n_1616), .B1(n_1617), .B2(n_1619), .C(n_1620), .Y(n_1615) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1065), .Y(n_1074) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1065), .Y(n_1162) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1065), .Y(n_1379) );
BUFx4f_ASAP7_75t_SL g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
AOI211x1_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1080), .B(n_1083), .C(n_1092), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1580 ( .A(n_1082), .Y(n_1580) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx6_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx5_ASAP7_75t_L g1193 ( .A(n_1089), .Y(n_1193) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVxp67_ASAP7_75t_L g1429 ( .A(n_1098), .Y(n_1429) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_1103), .A2(n_1149), .B1(n_1150), .B2(n_1201), .Y(n_1102) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1103), .Y(n_1201) );
OAI21x1_ASAP7_75t_SL g1103 ( .A1(n_1104), .A2(n_1105), .B(n_1148), .Y(n_1103) );
NAND4xp25_ASAP7_75t_L g1148 ( .A(n_1104), .B(n_1107), .C(n_1109), .D(n_1129), .Y(n_1148) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
NAND3xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1109), .C(n_1129), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1114), .Y(n_1109) );
NAND3xp33_ASAP7_75t_SL g1114 ( .A(n_1115), .B(n_1118), .C(n_1121), .Y(n_1114) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx2_ASAP7_75t_L g1475 ( .A(n_1127), .Y(n_1475) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND3xp33_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1136), .C(n_1142), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1135), .Y(n_1131) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
NOR3xp33_ASAP7_75t_L g1240 ( .A(n_1135), .B(n_1241), .C(n_1246), .Y(n_1240) );
NOR3xp33_ASAP7_75t_L g1258 ( .A(n_1135), .B(n_1259), .C(n_1264), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1138), .B1(n_1140), .B2(n_1141), .Y(n_1136) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
NOR2x1_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1178), .Y(n_1151) );
A2O1A1Ixp33_ASAP7_75t_L g1152 ( .A1(n_1153), .A2(n_1157), .B(n_1175), .C(n_1176), .Y(n_1152) );
NOR3xp33_ASAP7_75t_SL g1157 ( .A(n_1158), .B(n_1168), .C(n_1169), .Y(n_1157) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1164), .Y(n_1462) );
INVx2_ASAP7_75t_L g1465 ( .A(n_1164), .Y(n_1465) );
INVx2_ASAP7_75t_R g1501 ( .A(n_1164), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1167), .A2(n_1191), .B1(n_1192), .B2(n_1193), .Y(n_1190) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
O2A1O1Ixp5_ASAP7_75t_L g1900 ( .A1(n_1175), .A2(n_1901), .B(n_1913), .C(n_1921), .Y(n_1900) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1186), .Y(n_1178) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_1191), .A2(n_1193), .B1(n_1442), .B2(n_1443), .Y(n_1441) );
OAI22xp33_ASAP7_75t_L g1551 ( .A1(n_1193), .A2(n_1552), .B1(n_1553), .B2(n_1555), .Y(n_1551) );
XNOR2xp5_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1294), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
XNOR2x1_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1253), .Y(n_1204) );
XNOR2x1_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
NOR2x1_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1234), .Y(n_1207) );
NAND3xp33_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1228), .C(n_1232), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1227), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_1216), .A2(n_1226), .B1(n_1249), .B2(n_1250), .Y(n_1248) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1238), .Y(n_1276) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1249), .Y(n_1464) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
XNOR2x1_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1256), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1281), .Y(n_1256) );
INVx2_ASAP7_75t_L g1618 ( .A(n_1269), .Y(n_1618) );
OAI221xp5_ASAP7_75t_L g1903 ( .A1(n_1291), .A2(n_1562), .B1(n_1904), .B2(n_1905), .C(n_1906), .Y(n_1903) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_1295), .A2(n_1345), .B1(n_1392), .B2(n_1393), .Y(n_1294) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1295), .Y(n_1393) );
NAND2xp67_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1320), .Y(n_1296) );
NAND3xp33_ASAP7_75t_SL g1300 ( .A(n_1301), .B(n_1306), .C(n_1307), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1303), .B1(n_1304), .B2(n_1305), .Y(n_1301) );
AOI222xp33_ASAP7_75t_L g1333 ( .A1(n_1302), .A2(n_1304), .B1(n_1334), .B2(n_1335), .C1(n_1336), .C2(n_1340), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_1303), .A2(n_1305), .B1(n_1454), .B2(n_1455), .Y(n_1453) );
AOI22xp5_ASAP7_75t_L g1926 ( .A1(n_1303), .A2(n_1305), .B1(n_1927), .B2(n_1928), .Y(n_1926) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_1305), .A2(n_1507), .B1(n_1508), .B2(n_1509), .Y(n_1506) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1305), .Y(n_1605) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1311), .B1(n_1315), .B2(n_1318), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
NAND3xp33_ASAP7_75t_SL g1321 ( .A(n_1322), .B(n_1327), .C(n_1333), .Y(n_1321) );
AOI22xp5_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1324), .B1(n_1325), .B2(n_1326), .Y(n_1322) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1345), .Y(n_1392) );
XOR2x2_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1391), .Y(n_1345) );
NOR2x1_ASAP7_75t_SL g1346 ( .A(n_1347), .B(n_1370), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1359), .Y(n_1350) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVxp33_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
BUFx6f_ASAP7_75t_L g1911 ( .A(n_1364), .Y(n_1911) );
INVx2_ASAP7_75t_SL g1437 ( .A(n_1365), .Y(n_1437) );
A2O1A1Ixp33_ASAP7_75t_SL g1370 ( .A1(n_1371), .A2(n_1374), .B(n_1385), .C(n_1388), .Y(n_1370) );
NOR3xp33_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1381), .C(n_1384), .Y(n_1374) );
OAI21xp5_ASAP7_75t_L g1469 ( .A1(n_1385), .A2(n_1470), .B(n_1482), .Y(n_1469) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1387), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1390), .Y(n_1388) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1394), .Y(n_1651) );
AOI22xp5_ASAP7_75t_SL g1394 ( .A1(n_1395), .A2(n_1488), .B1(n_1649), .B2(n_1650), .Y(n_1394) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1395), .Y(n_1649) );
OA22x2_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1397), .B1(n_1448), .B2(n_1449), .Y(n_1395) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
NOR3xp33_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1417), .C(n_1418), .Y(n_1405) );
NOR3xp33_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1410), .C(n_1416), .Y(n_1406) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1409), .Y(n_1407) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1408), .B(n_1435), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1414), .Y(n_1410) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g1571 ( .A1(n_1420), .A2(n_1552), .B1(n_1561), .B2(n_1572), .Y(n_1571) );
INVx2_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
NAND3xp33_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1432), .C(n_1446), .Y(n_1427) );
AOI22xp5_ASAP7_75t_L g1432 ( .A1(n_1433), .A2(n_1438), .B1(n_1444), .B2(n_1445), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_1434), .A2(n_1439), .B1(n_1440), .B2(n_1441), .Y(n_1438) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1469), .Y(n_1450) );
NAND3xp33_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1456), .C(n_1459), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_1457), .A2(n_1458), .B1(n_1478), .B2(n_1480), .Y(n_1477) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx2_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1488), .Y(n_1650) );
XOR2xp5_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1527), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
HB1xp67_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1510), .Y(n_1492) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1508), .Y(n_1604) );
AOI21xp5_ASAP7_75t_L g1510 ( .A1(n_1511), .A2(n_1523), .B(n_1525), .Y(n_1510) );
NAND3xp33_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1515), .C(n_1520), .Y(n_1511) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
AOI22x1_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1529), .B1(n_1595), .B2(n_1647), .Y(n_1527) );
INVx2_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1530), .Y(n_1593) );
OAI211xp5_ASAP7_75t_L g1530 ( .A1(n_1531), .A2(n_1533), .B(n_1549), .C(n_1578), .Y(n_1530) );
CKINVDCx14_ASAP7_75t_R g1531 ( .A(n_1532), .Y(n_1531) );
NOR3xp33_ASAP7_75t_SL g1533 ( .A(n_1534), .B(n_1538), .C(n_1545), .Y(n_1533) );
INVx2_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g1581 ( .A1(n_1543), .A2(n_1582), .B1(n_1583), .B2(n_1584), .Y(n_1581) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1569), .Y(n_1549) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
OAI22xp5_ASAP7_75t_L g1560 ( .A1(n_1558), .A2(n_1561), .B1(n_1562), .B2(n_1564), .Y(n_1560) );
INVx5_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
OAI33xp33_ASAP7_75t_L g1569 ( .A1(n_1570), .A2(n_1571), .A3(n_1573), .B1(n_1575), .B2(n_1576), .B3(n_1577), .Y(n_1569) );
INVx2_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
HB1xp67_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVxp67_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
INVx2_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
AND3x2_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1624), .C(n_1627), .Y(n_1598) );
AOI211xp5_ASAP7_75t_SL g1599 ( .A1(n_1600), .A2(n_1601), .B(n_1603), .C(n_1606), .Y(n_1599) );
INVxp67_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
OAI22xp5_ASAP7_75t_L g1908 ( .A1(n_1630), .A2(n_1909), .B1(n_1910), .B2(n_1912), .Y(n_1908) );
INVx2_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVxp67_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
BUFx3_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx3_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
OR2x2_ASAP7_75t_L g1655 ( .A(n_1656), .B(n_1662), .Y(n_1655) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1660), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1949 ( .A(n_1658), .B(n_1661), .Y(n_1949) );
INVx1_ASAP7_75t_L g1953 ( .A(n_1658), .Y(n_1953) );
HB1xp67_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
NOR2xp33_ASAP7_75t_L g1955 ( .A(n_1661), .B(n_1953), .Y(n_1955) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
OAI221xp5_ASAP7_75t_L g1665 ( .A1(n_1666), .A2(n_1895), .B1(n_1898), .B2(n_1939), .C(n_1942), .Y(n_1665) );
AOI21xp5_ASAP7_75t_L g1666 ( .A1(n_1667), .A2(n_1809), .B(n_1862), .Y(n_1666) );
NAND4xp25_ASAP7_75t_L g1667 ( .A(n_1668), .B(n_1779), .C(n_1795), .D(n_1801), .Y(n_1667) );
NOR5xp2_ASAP7_75t_L g1668 ( .A(n_1669), .B(n_1733), .C(n_1746), .D(n_1753), .E(n_1776), .Y(n_1668) );
OAI21xp5_ASAP7_75t_SL g1669 ( .A1(n_1670), .A2(n_1690), .B(n_1709), .Y(n_1669) );
NOR2xp33_ASAP7_75t_L g1710 ( .A(n_1670), .B(n_1691), .Y(n_1710) );
OAI31xp33_ASAP7_75t_L g1887 ( .A1(n_1670), .A2(n_1888), .A3(n_1889), .B(n_1890), .Y(n_1887) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1808 ( .A(n_1671), .B(n_1766), .Y(n_1808) );
AOI221xp5_ASAP7_75t_L g1825 ( .A1(n_1671), .A2(n_1749), .B1(n_1826), .B2(n_1827), .C(n_1829), .Y(n_1825) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1672), .B(n_1686), .Y(n_1671) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1672), .Y(n_1736) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1672), .Y(n_1748) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1672), .Y(n_1794) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1672), .B(n_1724), .Y(n_1798) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1680), .Y(n_1672) );
AND2x6_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1676), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1675), .B(n_1679), .Y(n_1678) );
AND2x4_ASAP7_75t_L g1681 ( .A(n_1675), .B(n_1682), .Y(n_1681) );
AND2x6_ASAP7_75t_L g1684 ( .A(n_1675), .B(n_1685), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1675), .B(n_1679), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1770 ( .A(n_1675), .B(n_1679), .Y(n_1770) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1677), .B(n_1683), .Y(n_1682) );
INVx2_ASAP7_75t_L g1897 ( .A(n_1684), .Y(n_1897) );
HB1xp67_ASAP7_75t_L g1952 ( .A(n_1685), .Y(n_1952) );
CKINVDCx5p33_ASAP7_75t_R g1724 ( .A(n_1686), .Y(n_1724) );
OR2x2_ASAP7_75t_L g1745 ( .A(n_1686), .B(n_1721), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1686), .B(n_1736), .Y(n_1773) );
HB1xp67_ASAP7_75t_SL g1791 ( .A(n_1686), .Y(n_1791) );
NAND2xp5_ASAP7_75t_L g1855 ( .A(n_1686), .B(n_1766), .Y(n_1855) );
NAND2xp5_ASAP7_75t_L g1867 ( .A(n_1686), .B(n_1693), .Y(n_1867) );
AND2x4_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1689), .Y(n_1686) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1690), .Y(n_1878) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1696), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1802 ( .A(n_1691), .B(n_1728), .Y(n_1802) );
NAND2xp5_ASAP7_75t_L g1885 ( .A(n_1691), .B(n_1774), .Y(n_1885) );
CKINVDCx14_ASAP7_75t_R g1691 ( .A(n_1692), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1692), .B(n_1744), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1692), .B(n_1721), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1692), .B(n_1713), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1805 ( .A(n_1692), .B(n_1741), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1819 ( .A(n_1692), .B(n_1820), .Y(n_1819) );
NOR2xp33_ASAP7_75t_L g1831 ( .A(n_1692), .B(n_1745), .Y(n_1831) );
NOR2xp33_ASAP7_75t_L g1851 ( .A(n_1692), .B(n_1787), .Y(n_1851) );
NOR2xp33_ASAP7_75t_L g1861 ( .A(n_1692), .B(n_1754), .Y(n_1861) );
INVx3_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
CKINVDCx5p33_ASAP7_75t_R g1725 ( .A(n_1693), .Y(n_1725) );
NOR2xp33_ASAP7_75t_L g1762 ( .A(n_1693), .B(n_1730), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1693), .B(n_1698), .Y(n_1765) );
NAND2xp5_ASAP7_75t_L g1800 ( .A(n_1693), .B(n_1714), .Y(n_1800) );
AND2x2_ASAP7_75t_L g1835 ( .A(n_1693), .B(n_1807), .Y(n_1835) );
NAND2xp5_ASAP7_75t_L g1857 ( .A(n_1693), .B(n_1816), .Y(n_1857) );
NAND2xp5_ASAP7_75t_L g1859 ( .A(n_1693), .B(n_1741), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1889 ( .A(n_1693), .B(n_1787), .Y(n_1889) );
AND2x4_ASAP7_75t_SL g1693 ( .A(n_1694), .B(n_1695), .Y(n_1693) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1701), .Y(n_1697) );
INVx2_ASAP7_75t_L g1713 ( .A(n_1698), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1698), .B(n_1706), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1698), .B(n_1715), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1698), .B(n_1714), .Y(n_1790) );
AND2x2_ASAP7_75t_L g1813 ( .A(n_1698), .B(n_1814), .Y(n_1813) );
NAND2xp5_ASAP7_75t_L g1828 ( .A(n_1698), .B(n_1703), .Y(n_1828) );
OAI322xp33_ASAP7_75t_L g1829 ( .A1(n_1698), .A2(n_1712), .A3(n_1807), .B1(n_1830), .B2(n_1832), .C1(n_1836), .C2(n_1838), .Y(n_1829) );
OR2x2_ASAP7_75t_L g1865 ( .A(n_1698), .B(n_1800), .Y(n_1865) );
OR2x2_ASAP7_75t_L g1876 ( .A(n_1698), .B(n_1703), .Y(n_1876) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
OR2x2_ASAP7_75t_L g1775 ( .A(n_1701), .B(n_1713), .Y(n_1775) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1701), .Y(n_1816) );
OR2x2_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1706), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1702), .B(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
OR2x2_ASAP7_75t_L g1730 ( .A(n_1703), .B(n_1731), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1703), .B(n_1706), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1703), .B(n_1713), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1705), .Y(n_1703) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1706), .Y(n_1715) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1706), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1848 ( .A(n_1706), .B(n_1713), .Y(n_1848) );
NAND2x1_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1708), .Y(n_1706) );
AOI22xp33_ASAP7_75t_L g1709 ( .A1(n_1710), .A2(n_1711), .B1(n_1717), .B2(n_1726), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1716), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1713), .B(n_1714), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1713), .B(n_1729), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1713), .B(n_1741), .Y(n_1740) );
OR2x2_ASAP7_75t_L g1785 ( .A(n_1713), .B(n_1786), .Y(n_1785) );
OR2x2_ASAP7_75t_L g1821 ( .A(n_1713), .B(n_1730), .Y(n_1821) );
NOR2xp33_ASAP7_75t_L g1833 ( .A(n_1713), .B(n_1834), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1714), .B(n_1758), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1714), .B(n_1765), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1814 ( .A(n_1714), .B(n_1725), .Y(n_1814) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1716), .Y(n_1778) );
OAI21xp5_ASAP7_75t_L g1866 ( .A1(n_1716), .A2(n_1867), .B(n_1868), .Y(n_1866) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1725), .Y(n_1718) );
INVx1_ASAP7_75t_L g1894 ( .A(n_1719), .Y(n_1894) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
OR2x2_ASAP7_75t_L g1734 ( .A(n_1720), .B(n_1735), .Y(n_1734) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1724), .Y(n_1720) );
INVx2_ASAP7_75t_SL g1755 ( .A(n_1721), .Y(n_1755) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1721), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1722), .B(n_1723), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1754 ( .A(n_1724), .B(n_1755), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1724), .B(n_1748), .Y(n_1761) );
NOR2xp33_ASAP7_75t_L g1780 ( .A(n_1724), .B(n_1781), .Y(n_1780) );
OAI22xp5_ASAP7_75t_L g1811 ( .A1(n_1724), .A2(n_1791), .B1(n_1812), .B2(n_1815), .Y(n_1811) );
NAND3xp33_ASAP7_75t_L g1850 ( .A(n_1724), .B(n_1741), .C(n_1851), .Y(n_1850) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1725), .Y(n_1739) );
NAND2xp5_ASAP7_75t_L g1846 ( .A(n_1725), .B(n_1847), .Y(n_1846) );
INVxp33_ASAP7_75t_SL g1726 ( .A(n_1727), .Y(n_1726) );
NOR2xp33_ASAP7_75t_SL g1727 ( .A(n_1728), .B(n_1732), .Y(n_1727) );
INVx2_ASAP7_75t_L g1752 ( .A(n_1728), .Y(n_1752) );
AOI222xp33_ASAP7_75t_L g1801 ( .A1(n_1729), .A2(n_1802), .B1(n_1803), .B2(n_1804), .C1(n_1806), .C2(n_1808), .Y(n_1801) );
NOR2xp33_ASAP7_75t_L g1837 ( .A(n_1729), .B(n_1816), .Y(n_1837) );
A2O1A1Ixp33_ASAP7_75t_L g1890 ( .A1(n_1729), .A2(n_1739), .B(n_1808), .C(n_1820), .Y(n_1890) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
A2O1A1Ixp33_ASAP7_75t_L g1891 ( .A1(n_1732), .A2(n_1803), .B(n_1831), .C(n_1892), .Y(n_1891) );
OAI21xp5_ASAP7_75t_SL g1733 ( .A1(n_1734), .A2(n_1737), .B(n_1742), .Y(n_1733) );
INVx1_ASAP7_75t_L g1886 ( .A(n_1734), .Y(n_1886) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1736), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1824 ( .A(n_1736), .B(n_1783), .Y(n_1824) );
AND2x2_ASAP7_75t_L g1826 ( .A(n_1736), .B(n_1744), .Y(n_1826) );
NAND2xp5_ASAP7_75t_L g1873 ( .A(n_1736), .B(n_1874), .Y(n_1873) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1739), .B(n_1740), .Y(n_1738) );
AOI221xp5_ASAP7_75t_L g1877 ( .A1(n_1740), .A2(n_1843), .B1(n_1878), .B2(n_1879), .C(n_1880), .Y(n_1877) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1741), .B(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1741), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1870 ( .A(n_1741), .B(n_1765), .Y(n_1870) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1743), .B(n_1778), .Y(n_1777) );
NAND2xp5_ASAP7_75t_L g1792 ( .A(n_1743), .B(n_1793), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1844 ( .A(n_1744), .B(n_1803), .Y(n_1844) );
INVx2_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
AOI21xp33_ASAP7_75t_L g1810 ( .A1(n_1745), .A2(n_1811), .B(n_1817), .Y(n_1810) );
INVxp67_ASAP7_75t_SL g1746 ( .A(n_1747), .Y(n_1746) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1748), .B(n_1749), .Y(n_1747) );
NOR2xp33_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1752), .Y(n_1749) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
OAI21xp33_ASAP7_75t_L g1772 ( .A1(n_1751), .A2(n_1773), .B(n_1774), .Y(n_1772) );
OAI211xp5_ASAP7_75t_SL g1753 ( .A1(n_1754), .A2(n_1756), .B(n_1760), .C(n_1772), .Y(n_1753) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1754), .Y(n_1879) );
INVx2_ASAP7_75t_L g1787 ( .A(n_1755), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1869 ( .A(n_1755), .B(n_1870), .Y(n_1869) );
O2A1O1Ixp33_ASAP7_75t_SL g1880 ( .A1(n_1755), .A2(n_1822), .B(n_1881), .C(n_1882), .Y(n_1880) );
CKINVDCx14_ASAP7_75t_R g1756 ( .A(n_1757), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1815 ( .A(n_1758), .B(n_1816), .Y(n_1815) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
OR2x2_ASAP7_75t_L g1822 ( .A(n_1759), .B(n_1786), .Y(n_1822) );
AOI211xp5_ASAP7_75t_L g1871 ( .A1(n_1759), .A2(n_1872), .B(n_1873), .C(n_1875), .Y(n_1871) );
AOI221xp5_ASAP7_75t_L g1760 ( .A1(n_1761), .A2(n_1762), .B1(n_1763), .B2(n_1766), .C(n_1767), .Y(n_1760) );
NOR2xp33_ASAP7_75t_L g1784 ( .A(n_1761), .B(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1761), .Y(n_1838) );
O2A1O1Ixp33_ASAP7_75t_L g1883 ( .A1(n_1762), .A2(n_1884), .B(n_1886), .C(n_1887), .Y(n_1883) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1782 ( .A(n_1764), .B(n_1783), .Y(n_1782) );
INVx2_ASAP7_75t_L g1783 ( .A(n_1766), .Y(n_1783) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1767), .B(n_1850), .Y(n_1849) );
INVx3_ASAP7_75t_L g1767 ( .A(n_1768), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1768 ( .A(n_1769), .B(n_1771), .Y(n_1768) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1773), .Y(n_1882) );
INVx2_ASAP7_75t_L g1774 ( .A(n_1775), .Y(n_1774) );
INVxp67_ASAP7_75t_SL g1776 ( .A(n_1777), .Y(n_1776) );
O2A1O1Ixp33_ASAP7_75t_L g1779 ( .A1(n_1780), .A2(n_1784), .B(n_1787), .C(n_1788), .Y(n_1779) );
OAI31xp33_ASAP7_75t_L g1795 ( .A1(n_1780), .A2(n_1784), .A3(n_1796), .B(n_1799), .Y(n_1795) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1783), .B(n_1807), .Y(n_1806) );
OR2x2_ASAP7_75t_L g1842 ( .A(n_1783), .B(n_1807), .Y(n_1842) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1785), .Y(n_1840) );
NAND2xp5_ASAP7_75t_L g1797 ( .A(n_1787), .B(n_1798), .Y(n_1797) );
O2A1O1Ixp33_ASAP7_75t_L g1788 ( .A1(n_1789), .A2(n_1791), .B(n_1792), .C(n_1794), .Y(n_1788) );
AOI21xp33_ASAP7_75t_L g1892 ( .A1(n_1789), .A2(n_1893), .B(n_1894), .Y(n_1892) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1860 ( .A(n_1793), .B(n_1861), .Y(n_1860) );
CKINVDCx14_ASAP7_75t_R g1888 ( .A(n_1793), .Y(n_1888) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1794), .Y(n_1803) );
AOI221xp5_ASAP7_75t_L g1863 ( .A1(n_1794), .A2(n_1826), .B1(n_1864), .B2(n_1866), .C(n_1871), .Y(n_1863) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1799), .Y(n_1881) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1802), .Y(n_1893) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
AOI222xp33_ASAP7_75t_L g1852 ( .A1(n_1806), .A2(n_1841), .B1(n_1853), .B2(n_1854), .C1(n_1856), .C2(n_1858), .Y(n_1852) );
NAND5xp2_ASAP7_75t_L g1809 ( .A(n_1810), .B(n_1825), .C(n_1839), .D(n_1852), .E(n_1860), .Y(n_1809) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVxp67_ASAP7_75t_SL g1872 ( .A(n_1814), .Y(n_1872) );
AOI21xp33_ASAP7_75t_L g1817 ( .A1(n_1818), .A2(n_1822), .B(n_1823), .Y(n_1817) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1822), .Y(n_1853) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
INVxp67_ASAP7_75t_SL g1830 ( .A(n_1831), .Y(n_1830) );
INVxp67_ASAP7_75t_L g1832 ( .A(n_1833), .Y(n_1832) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
HB1xp67_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
AOI221xp5_ASAP7_75t_L g1839 ( .A1(n_1840), .A2(n_1841), .B1(n_1843), .B2(n_1845), .C(n_1849), .Y(n_1839) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1844), .Y(n_1843) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1855), .Y(n_1874) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1857), .Y(n_1856) );
INVxp67_ASAP7_75t_SL g1858 ( .A(n_1859), .Y(n_1858) );
NAND4xp25_ASAP7_75t_L g1862 ( .A(n_1863), .B(n_1877), .C(n_1883), .D(n_1891), .Y(n_1862) );
INVxp67_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1876), .Y(n_1875) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
CKINVDCx20_ASAP7_75t_R g1895 ( .A(n_1896), .Y(n_1895) );
CKINVDCx20_ASAP7_75t_R g1896 ( .A(n_1897), .Y(n_1896) );
INVx1_ASAP7_75t_L g1945 ( .A(n_1899), .Y(n_1945) );
NAND3x1_ASAP7_75t_L g1899 ( .A(n_1900), .B(n_1923), .C(n_1925), .Y(n_1899) );
INVx1_ASAP7_75t_L g1906 ( .A(n_1907), .Y(n_1906) );
BUFx2_ASAP7_75t_L g1910 ( .A(n_1911), .Y(n_1910) );
NAND2xp5_ASAP7_75t_L g1929 ( .A(n_1930), .B(n_1931), .Y(n_1929) );
INVx3_ASAP7_75t_L g1939 ( .A(n_1940), .Y(n_1939) );
INVxp33_ASAP7_75t_L g1943 ( .A(n_1944), .Y(n_1943) );
HB1xp67_ASAP7_75t_L g1947 ( .A(n_1948), .Y(n_1947) );
BUFx3_ASAP7_75t_L g1948 ( .A(n_1949), .Y(n_1948) );
HB1xp67_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
OAI21xp5_ASAP7_75t_L g1951 ( .A1(n_1952), .A2(n_1953), .B(n_1954), .Y(n_1951) );
INVx1_ASAP7_75t_L g1954 ( .A(n_1955), .Y(n_1954) );
endmodule