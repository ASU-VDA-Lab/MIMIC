module fake_jpeg_6923_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_27),
.B2(n_32),
.Y(n_48)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_62),
.B1(n_46),
.B2(n_24),
.Y(n_99)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_41),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_27),
.B1(n_26),
.B2(n_20),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_24),
.B(n_18),
.C(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_79),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_87),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_43),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_54),
.B1(n_37),
.B2(n_51),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_73),
.B1(n_72),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_104),
.B1(n_115),
.B2(n_97),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_61),
.C(n_56),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_126),
.C(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_61),
.B1(n_60),
.B2(n_45),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_127),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_17),
.B(n_19),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_79),
.B(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_92),
.B1(n_84),
.B2(n_89),
.Y(n_129)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_113),
.Y(n_145)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_40),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_54),
.B1(n_37),
.B2(n_51),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_43),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_125),
.B(n_28),
.Y(n_142)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_18),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_31),
.Y(n_150)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_43),
.B(n_20),
.C(n_33),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_40),
.C(n_39),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_131),
.B1(n_137),
.B2(n_143),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_144),
.C(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_87),
.B1(n_89),
.B2(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_116),
.B1(n_110),
.B2(n_101),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_24),
.B1(n_26),
.B2(n_20),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_33),
.B(n_25),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_136),
.A2(n_139),
.B(n_142),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_55),
.B1(n_52),
.B2(n_26),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_R g139 ( 
.A(n_123),
.B(n_40),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_40),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_40),
.C(n_44),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_152),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_33),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_106),
.Y(n_175)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_156),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_25),
.B(n_28),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_182),
.C(n_25),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_154),
.B1(n_139),
.B2(n_151),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_174),
.B1(n_128),
.B2(n_44),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_108),
.Y(n_170)
);

BUFx4f_ASAP7_75t_SL g171 ( 
.A(n_148),
.Y(n_171)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_173),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_124),
.B1(n_112),
.B2(n_113),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_177),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_103),
.B1(n_122),
.B2(n_117),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_149),
.B1(n_105),
.B2(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_44),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_134),
.B(n_140),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_187),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_21),
.B(n_28),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_31),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_39),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_193),
.A2(n_198),
.B1(n_167),
.B2(n_171),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_178),
.A2(n_160),
.B(n_181),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_202),
.B1(n_203),
.B2(n_211),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_149),
.B1(n_105),
.B2(n_156),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_210),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_29),
.B(n_128),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_138),
.B1(n_29),
.B2(n_31),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_179),
.C(n_166),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_174),
.C(n_161),
.Y(n_235)
);

OAI22x1_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_31),
.B1(n_69),
.B2(n_39),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_30),
.B1(n_23),
.B2(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_29),
.B(n_31),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_171),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_185),
.A2(n_100),
.B(n_69),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_176),
.B1(n_211),
.B2(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_222),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_164),
.Y(n_227)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_230),
.B1(n_204),
.B2(n_187),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_233),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_173),
.B1(n_161),
.B2(n_157),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_196),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_202),
.B(n_191),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_30),
.C(n_1),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_159),
.C(n_158),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_243),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_226),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_197),
.B1(n_205),
.B2(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_220),
.B(n_227),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_190),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_260),
.C(n_264),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_205),
.B1(n_199),
.B2(n_188),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_256),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_203),
.B1(n_30),
.B2(n_23),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_30),
.B1(n_1),
.B2(n_3),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_215),
.B1(n_238),
.B2(n_221),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_262),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_240),
.B1(n_228),
.B2(n_214),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_0),
.C(n_1),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_263),
.B(n_219),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_281),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_217),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_249),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_273),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_232),
.C(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_280),
.C(n_282),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_222),
.B(n_10),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_253),
.B1(n_256),
.B2(n_254),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_247),
.B(n_10),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_3),
.C(n_4),
.Y(n_282)
);

INVxp33_ASAP7_75t_SL g286 ( 
.A(n_277),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_252),
.B1(n_255),
.B2(n_245),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_261),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_296),
.B(n_12),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_244),
.B1(n_254),
.B2(n_250),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_257),
.B1(n_248),
.B2(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_260),
.C(n_243),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_4),
.C(n_5),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_264),
.Y(n_296)
);

OAI321xp33_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_267),
.A3(n_280),
.B1(n_272),
.B2(n_270),
.C(n_283),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_303),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_270),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_306),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_11),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_310),
.C(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_4),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_16),
.B(n_15),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_308),
.B(n_312),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_284),
.B(n_15),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_15),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_299),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_5),
.C(n_6),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_12),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_293),
.Y(n_317)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_285),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_303),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_5),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_311),
.B(n_13),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_326),
.B(n_330),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_331),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_305),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_13),
.C(n_6),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_335),
.C(n_336),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_329),
.B(n_315),
.C(n_322),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_333),
.Y(n_339)
);

OAI321xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_337),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_5),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.B(n_7),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_7),
.B(n_8),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_8),
.B(n_341),
.Y(n_343)
);


endmodule