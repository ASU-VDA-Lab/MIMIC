module fake_jpeg_28063_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_17),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_6),
.B1(n_13),
.B2(n_21),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_5),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_23),
.C(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_9),
.B(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_21),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_28),
.B1(n_15),
.B2(n_19),
.Y(n_34)
);

XNOR2x1_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_30),
.B1(n_24),
.B2(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_34),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_26),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.C(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_39),
.C(n_36),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_28),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_43),
.B(n_40),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_29),
.C(n_16),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_23),
.B(n_6),
.Y(n_46)
);


endmodule