module fake_jpeg_20433_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_27),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_57),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_53),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_10),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_23),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_40),
.B1(n_28),
.B2(n_21),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_29),
.B1(n_43),
.B2(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_71),
.B(n_78),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_26),
.C(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_18),
.B1(n_30),
.B2(n_15),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_74),
.A2(n_86),
.B(n_83),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_31),
.B1(n_23),
.B2(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_76),
.B(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_18),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_30),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_62),
.B(n_63),
.C(n_15),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_84),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_11),
.B1(n_13),
.B2(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_45),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_11),
.B1(n_55),
.B2(n_60),
.Y(n_114)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_8),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_60),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_1),
.B1(n_8),
.B2(n_9),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_11),
.B1(n_13),
.B2(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_9),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx6f_ASAP7_75t_SL g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_115),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_97),
.B1(n_82),
.B2(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_87),
.B1(n_69),
.B2(n_67),
.Y(n_128)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_97),
.C(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_66),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_72),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_132),
.B1(n_135),
.B2(n_141),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_79),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_135),
.C(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_68),
.B1(n_76),
.B2(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_89),
.B1(n_82),
.B2(n_66),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_85),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_86),
.B1(n_121),
.B2(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_105),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_147),
.B(n_104),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_111),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_122),
.C(n_118),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_127),
.C(n_132),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_109),
.B(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_99),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_100),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_163),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_128),
.B1(n_142),
.B2(n_144),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_164),
.B1(n_131),
.B2(n_109),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_122),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_107),
.B1(n_103),
.B2(n_114),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_170),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_127),
.CI(n_116),
.CON(n_167),
.SN(n_167)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_172),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_107),
.B(n_131),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_150),
.B(n_164),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_131),
.B1(n_133),
.B2(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_175),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_101),
.C(n_106),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_113),
.C(n_103),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_115),
.C(n_109),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_148),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_175),
.B1(n_148),
.B2(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_176),
.B(n_178),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

XOR2x1_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_162),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_154),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_167),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_170),
.C(n_174),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_188),
.C(n_187),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_197),
.B(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_158),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_161),
.B1(n_180),
.B2(n_182),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_161),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_190),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_204),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_203),
.C(n_193),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_208),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_198),
.C(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

OAI221xp5_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_166),
.B1(n_155),
.B2(n_156),
.C(n_201),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_191),
.B(n_200),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_191),
.B(n_205),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_210),
.B(n_125),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_108),
.Y(n_216)
);


endmodule