module fake_aes_5639_n_494 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_494);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_494;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g70 ( .A(n_23), .Y(n_70) );
HB1xp67_ASAP7_75t_L g71 ( .A(n_65), .Y(n_71) );
INVxp67_ASAP7_75t_SL g72 ( .A(n_56), .Y(n_72) );
CKINVDCx16_ASAP7_75t_R g73 ( .A(n_2), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_47), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_52), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_60), .Y(n_76) );
OR2x2_ASAP7_75t_L g77 ( .A(n_39), .B(n_17), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_26), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_51), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_18), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_33), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_68), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_48), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_18), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_32), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_38), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_17), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_37), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_30), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_40), .B(n_2), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_45), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_10), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_66), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_11), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_100), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_86), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_80), .B(n_0), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_80), .B(n_1), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_100), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_100), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_86), .Y(n_115) );
INVx3_ASAP7_75t_L g116 ( .A(n_101), .Y(n_116) );
CKINVDCx8_ASAP7_75t_R g117 ( .A(n_73), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_100), .B(n_3), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_90), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
INVx6_ASAP7_75t_L g122 ( .A(n_100), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_75), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_81), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_71), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_103), .B(n_3), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_94), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_76), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_117), .A2(n_81), .B1(n_93), .B2(n_107), .Y(n_131) );
BUFx4f_ASAP7_75t_L g132 ( .A(n_120), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_120), .B(n_78), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_121), .B(n_77), .Y(n_134) );
INVx8_ASAP7_75t_L g135 ( .A(n_116), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_123), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_123), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g141 ( .A(n_121), .B(n_77), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_125), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_123), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
INVx2_ASAP7_75t_SL g146 ( .A(n_116), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_124), .A2(n_107), .B1(n_108), .B2(n_98), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_109), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_126), .B(n_101), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_123), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_110), .B(n_93), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
NOR3xp33_ASAP7_75t_SL g156 ( .A(n_131), .B(n_115), .C(n_128), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_136), .A2(n_126), .B1(n_127), .B2(n_111), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_134), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_143), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_136), .B(n_127), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_154), .A2(n_112), .B1(n_94), .B2(n_119), .Y(n_164) );
OR2x6_ASAP7_75t_L g165 ( .A(n_134), .B(n_112), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_149), .B(n_124), .Y(n_166) );
NOR3xp33_ASAP7_75t_SL g167 ( .A(n_131), .B(n_118), .C(n_97), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_132), .B(n_129), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_132), .A2(n_130), .B1(n_129), .B2(n_88), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_132), .B(n_87), .Y(n_173) );
OR2x6_ASAP7_75t_L g174 ( .A(n_141), .B(n_117), .Y(n_174) );
AND2x6_ASAP7_75t_L g175 ( .A(n_153), .B(n_78), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_149), .B(n_129), .Y(n_178) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_132), .B(n_105), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_154), .Y(n_180) );
NAND2x2_ASAP7_75t_L g181 ( .A(n_153), .B(n_4), .Y(n_181) );
NOR2x1_ASAP7_75t_L g182 ( .A(n_149), .B(n_130), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_133), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_169), .A2(n_132), .B(n_146), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_155), .A2(n_133), .B1(n_138), .B2(n_140), .Y(n_190) );
INVx5_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_160), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_158), .A2(n_162), .B1(n_170), .B2(n_177), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_168), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_186), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_184), .B(n_146), .Y(n_197) );
INVx5_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_160), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_185), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_169), .A2(n_146), .B(n_135), .Y(n_201) );
CKINVDCx8_ASAP7_75t_R g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_172), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_176), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_165), .A2(n_138), .B1(n_140), .B2(n_135), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_160), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_165), .A2(n_138), .B1(n_140), .B2(n_135), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_185), .Y(n_209) );
AOI221xp5_ASAP7_75t_L g210 ( .A1(n_166), .A2(n_147), .B1(n_130), .B2(n_79), .C(n_82), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_163), .B(n_140), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_175), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_182), .Y(n_215) );
AOI21xp5_ASAP7_75t_SL g216 ( .A1(n_165), .A2(n_72), .B(n_140), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_175), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_191), .Y(n_218) );
AO31x2_ASAP7_75t_L g219 ( .A1(n_188), .A2(n_166), .A3(n_113), .B(n_83), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
OAI211xp5_ASAP7_75t_SL g221 ( .A1(n_210), .A2(n_156), .B(n_164), .C(n_157), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_202), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_210), .A2(n_174), .B1(n_175), .B2(n_181), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_188), .A2(n_150), .B(n_145), .Y(n_225) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_201), .A2(n_173), .B(n_179), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_194), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_194), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_187), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_209), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_209), .B(n_163), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_209), .B(n_204), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g233 ( .A1(n_204), .A2(n_174), .B1(n_175), .B2(n_180), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_205), .A2(n_174), .B1(n_171), .B2(n_147), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g235 ( .A1(n_213), .A2(n_173), .B1(n_179), .B2(n_82), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_209), .B(n_171), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_213), .A2(n_183), .B1(n_79), .B2(n_83), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_187), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_191), .B(n_156), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_201), .A2(n_85), .B(n_106), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_193), .A2(n_167), .B1(n_84), .B2(n_85), .Y(n_243) );
OAI211xp5_ASAP7_75t_SL g244 ( .A1(n_223), .A2(n_167), .B(n_202), .C(n_215), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_231), .B(n_205), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_232), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g247 ( .A1(n_238), .A2(n_213), .B1(n_198), .B2(n_191), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_214), .B1(n_215), .B2(n_211), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_231), .B(n_214), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_220), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_238), .A2(n_216), .B(n_195), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_233), .A2(n_213), .B1(n_208), .B2(n_206), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_225), .A2(n_216), .B(n_212), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g254 ( .A1(n_221), .A2(n_190), .B1(n_192), .B2(n_207), .C(n_199), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_229), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_232), .B(n_192), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_191), .B1(n_198), .B2(n_196), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g258 ( .A1(n_243), .A2(n_191), .B1(n_198), .B2(n_217), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_232), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_220), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_218), .B(n_191), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_231), .B(n_198), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_229), .Y(n_264) );
OAI211xp5_ASAP7_75t_SL g265 ( .A1(n_234), .A2(n_70), .B(n_104), .C(n_89), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_246), .B(n_219), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_251), .A2(n_225), .B(n_242), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_262), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_244), .A2(n_233), .B1(n_243), .B2(n_237), .Y(n_269) );
OAI221xp5_ASAP7_75t_L g270 ( .A1(n_265), .A2(n_234), .B1(n_244), .B2(n_257), .C(n_248), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_260), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_255), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_265), .A2(n_263), .B1(n_247), .B2(n_259), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_262), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_255), .B(n_236), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_247), .A2(n_235), .B1(n_237), .B2(n_239), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_264), .B(n_219), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_246), .A2(n_237), .B1(n_240), .B2(n_235), .Y(n_278) );
NOR2xp33_ASAP7_75t_R g279 ( .A(n_263), .B(n_222), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_250), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_263), .A2(n_240), .B1(n_230), .B2(n_218), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_245), .A2(n_227), .B1(n_228), .B2(n_240), .C(n_239), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_259), .A2(n_236), .B1(n_240), .B2(n_230), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_260), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_250), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_285), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_275), .B(n_245), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_281), .B(n_272), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_281), .B(n_219), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_268), .B(n_261), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_266), .B(n_219), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_275), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g295 ( .A(n_277), .B(n_99), .C(n_91), .Y(n_295) );
AOI211x1_ASAP7_75t_L g296 ( .A1(n_270), .A2(n_277), .B(n_276), .C(n_254), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_276), .A2(n_258), .B1(n_252), .B2(n_256), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_272), .B(n_219), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_266), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_269), .B(n_102), .C(n_92), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_279), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_271), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_267), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_278), .B(n_106), .C(n_84), .D(n_96), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_219), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
AO31x2_ASAP7_75t_L g311 ( .A1(n_284), .A2(n_251), .A3(n_252), .B(n_241), .Y(n_311) );
AOI31xp33_ASAP7_75t_L g312 ( .A1(n_273), .A2(n_240), .A3(n_258), .B(n_262), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_268), .B(n_219), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_304), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_302), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_300), .B(n_274), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_300), .B(n_274), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_294), .B(n_274), .Y(n_320) );
NAND2xp33_ASAP7_75t_SL g321 ( .A(n_303), .B(n_284), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_296), .B(n_273), .Y(n_322) );
NAND4xp25_ASAP7_75t_SL g323 ( .A(n_303), .B(n_283), .C(n_270), .D(n_282), .Y(n_323) );
AOI33xp33_ASAP7_75t_L g324 ( .A1(n_306), .A2(n_95), .A3(n_249), .B1(n_113), .B2(n_228), .B3(n_227), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_289), .B(n_219), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_288), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_298), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_307), .B(n_254), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_313), .B(n_287), .Y(n_329) );
AND2x4_ASAP7_75t_SL g330 ( .A(n_292), .B(n_250), .Y(n_330) );
NOR2x1_ASAP7_75t_L g331 ( .A(n_295), .B(n_261), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_293), .B(n_267), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_312), .A2(n_297), .B(n_267), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_290), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_291), .B(n_249), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_313), .B(n_267), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_291), .B(n_261), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_290), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_299), .B(n_280), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_309), .B(n_280), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_309), .B(n_250), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_299), .B(n_250), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_314), .Y(n_346) );
CKINVDCx16_ASAP7_75t_R g347 ( .A(n_292), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_305), .B(n_250), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_310), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_301), .B(n_4), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_292), .A2(n_262), .B1(n_250), .B2(n_218), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_311), .Y(n_353) );
OAI221xp5_ASAP7_75t_SL g354 ( .A1(n_334), .A2(n_230), .B1(n_311), .B2(n_113), .C(n_224), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_316), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_315), .B(n_5), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_339), .B(n_311), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_347), .B(n_311), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_339), .B(n_311), .Y(n_359) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_335), .A2(n_152), .B(n_150), .C(n_145), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_338), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_330), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_323), .B(n_242), .C(n_253), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_318), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g365 ( .A1(n_351), .A2(n_230), .B(n_224), .C(n_241), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_336), .B(n_280), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_330), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_350), .B(n_280), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_327), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_321), .B(n_280), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_328), .A2(n_242), .B1(n_253), .B2(n_241), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_341), .Y(n_374) );
OAI22xp33_ASAP7_75t_SL g375 ( .A1(n_322), .A2(n_230), .B1(n_122), .B2(n_224), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_341), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_332), .B(n_253), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_328), .A2(n_226), .B1(n_199), .B2(n_207), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_325), .A2(n_144), .B(n_137), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_320), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_331), .A2(n_212), .B1(n_198), .B2(n_217), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_321), .Y(n_382) );
AOI322xp5_ASAP7_75t_L g383 ( .A1(n_351), .A2(n_109), .A3(n_114), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_12), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_329), .B(n_5), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g385 ( .A1(n_332), .A2(n_198), .B1(n_212), .B2(n_8), .C1(n_9), .C2(n_13), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_349), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_337), .B(n_109), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_344), .A2(n_226), .B1(n_212), .B2(n_203), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_317), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_329), .B(n_6), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_324), .B(n_6), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_324), .B(n_7), .Y(n_392) );
OAI32xp33_ASAP7_75t_L g393 ( .A1(n_344), .A2(n_340), .A3(n_343), .B1(n_319), .B2(n_353), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_327), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_345), .B(n_13), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_343), .B(n_14), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_333), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_SL g398 ( .A1(n_353), .A2(n_14), .B(n_15), .C(n_16), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_333), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_342), .B(n_15), .Y(n_400) );
XOR2x2_ASAP7_75t_L g401 ( .A(n_356), .B(n_352), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_361), .A2(n_348), .B1(n_122), .B2(n_109), .C(n_114), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_380), .B(n_16), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_362), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_358), .B(n_114), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_389), .B(n_114), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_371), .B(n_114), .Y(n_410) );
NOR2xp33_ASAP7_75t_R g411 ( .A(n_382), .B(n_21), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_384), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_368), .B(n_114), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_386), .B(n_109), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_375), .A2(n_226), .B(n_198), .Y(n_415) );
NOR2xp33_ASAP7_75t_SL g416 ( .A(n_384), .B(n_189), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_357), .B(n_144), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_372), .A2(n_189), .B(n_203), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_364), .B(n_122), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_394), .Y(n_421) );
NOR4xp25_ASAP7_75t_SL g422 ( .A(n_354), .B(n_122), .C(n_137), .D(n_27), .Y(n_422) );
XOR2x2_ASAP7_75t_L g423 ( .A(n_390), .B(n_22), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_366), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_383), .B(n_148), .C(n_151), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_400), .A2(n_189), .B1(n_200), .B2(n_196), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_387), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_396), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_395), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_397), .B(n_24), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_399), .B(n_28), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
AOI21xp33_ASAP7_75t_SL g433 ( .A1(n_393), .A2(n_29), .B(n_31), .Y(n_433) );
OA22x2_ASAP7_75t_L g434 ( .A1(n_359), .A2(n_197), .B1(n_203), .B2(n_195), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_359), .B(n_151), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_407), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_401), .A2(n_363), .B1(n_392), .B2(n_391), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_407), .B(n_377), .Y(n_441) );
OAI21xp33_ASAP7_75t_SL g442 ( .A1(n_434), .A2(n_388), .B(n_377), .Y(n_442) );
OAI22xp33_ASAP7_75t_L g443 ( .A1(n_416), .A2(n_378), .B1(n_381), .B2(n_385), .Y(n_443) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_411), .B(n_381), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_401), .A2(n_423), .B1(n_429), .B2(n_434), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_406), .B(n_365), .C(n_398), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_404), .B(n_360), .C(n_151), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_409), .B(n_379), .Y(n_448) );
XNOR2xp5_ASAP7_75t_L g449 ( .A(n_423), .B(n_373), .Y(n_449) );
XOR2xp5_ASAP7_75t_L g450 ( .A(n_429), .B(n_35), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_411), .A2(n_200), .B(n_196), .C(n_195), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_435), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_433), .B(n_200), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_412), .A2(n_148), .B1(n_142), .B2(n_152), .C(n_139), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_437), .A2(n_200), .B1(n_196), .B2(n_197), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_421), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_428), .A2(n_139), .B1(n_152), .B2(n_197), .C(n_200), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_454), .B(n_406), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_444), .A2(n_405), .B1(n_437), .B2(n_432), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_445), .A2(n_428), .B1(n_406), .B2(n_427), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_442), .A2(n_438), .B1(n_426), .B2(n_408), .C(n_425), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_455), .Y(n_465) );
OAI32xp33_ASAP7_75t_L g466 ( .A1(n_446), .A2(n_403), .A3(n_410), .B1(n_417), .B2(n_419), .Y(n_466) );
AOI322xp5_ASAP7_75t_L g467 ( .A1(n_443), .A2(n_421), .A3(n_420), .B1(n_413), .B2(n_414), .C1(n_430), .C2(n_431), .Y(n_467) );
NAND2x1_ASAP7_75t_SL g468 ( .A(n_439), .B(n_420), .Y(n_468) );
OAI322xp33_ASAP7_75t_L g469 ( .A1(n_440), .A2(n_415), .A3(n_418), .B1(n_422), .B2(n_139), .C1(n_46), .C2(n_49), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_449), .A2(n_197), .B1(n_139), .B2(n_42), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_452), .B(n_36), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_441), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_450), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_447), .A2(n_41), .B1(n_43), .B2(n_53), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_448), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_451), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_456), .A2(n_54), .B(n_55), .C(n_57), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_460), .B(n_58), .C(n_59), .D(n_62), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_453), .A2(n_67), .B1(n_69), .B2(n_458), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g480 ( .A1(n_459), .A2(n_442), .B1(n_444), .B2(n_449), .C1(n_356), .C2(n_401), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g481 ( .A1(n_457), .A2(n_442), .B1(n_444), .B2(n_449), .C1(n_356), .C2(n_401), .Y(n_481) );
NAND5xp2_ASAP7_75t_L g482 ( .A(n_481), .B(n_480), .C(n_464), .D(n_463), .E(n_462), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_467), .B(n_464), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_461), .B(n_475), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_465), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_475), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_482), .A2(n_466), .B1(n_469), .B2(n_473), .C(n_472), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_483), .A2(n_461), .B1(n_471), .B2(n_470), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_486), .A2(n_468), .B1(n_474), .B2(n_478), .C(n_479), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_488), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_489), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_490), .Y(n_492) );
AOI22xp5_ASAP7_75t_SL g493 ( .A1(n_492), .A2(n_491), .B1(n_486), .B2(n_487), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_493), .A2(n_484), .B1(n_485), .B2(n_476), .C(n_477), .Y(n_494) );
endmodule