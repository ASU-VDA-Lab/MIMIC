module fake_jpeg_28609_n_82 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_1),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_1),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_27),
.B1(n_17),
.B2(n_20),
.C(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_3),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

XNOR2x2_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_21),
.B(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_21),
.B1(n_15),
.B2(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_12),
.B1(n_15),
.B2(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_14),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_19),
.B1(n_20),
.B2(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_36),
.C(n_19),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_41),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_8),
.B(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_52),
.C(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_6),
.C(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_58),
.B1(n_54),
.B2(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_42),
.B1(n_32),
.B2(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_15),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_60),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_74),
.C(n_6),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_69),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_70),
.C(n_66),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_77),
.C(n_71),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_81),
.Y(n_82)
);


endmodule