module fake_jpeg_5308_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_0),
.B(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_27),
.B(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_39),
.B1(n_13),
.B2(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_10),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_56),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_15),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_29),
.A2(n_13),
.B1(n_15),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_59),
.B1(n_48),
.B2(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_34),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_53),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_73),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_66),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_55),
.C(n_41),
.Y(n_65)
);

NAND2x1p5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_62),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_72),
.B(n_68),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.C(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_70),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_69),
.B1(n_72),
.B2(n_68),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_86),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_71),
.B(n_63),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_67),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_87),
.C(n_85),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_86),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_93),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_96),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_100),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_103),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_105),
.Y(n_110)
);


endmodule