module fake_jpeg_13977_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_10),
.B(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_23),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_48),
.B(n_45),
.C(n_59),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_45),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_19),
.B1(n_42),
.B2(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_57),
.B1(n_51),
.B2(n_55),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_63),
.B1(n_61),
.B2(n_58),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_2),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_49),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_72),
.B1(n_71),
.B2(n_73),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_97),
.B1(n_95),
.B2(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_9),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_17),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_99),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_20),
.B1(n_40),
.B2(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

AO21x2_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_30),
.B(n_37),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_12),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_6),
.B(n_7),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_8),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_9),
.C(n_10),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_113),
.B1(n_31),
.B2(n_44),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_96),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_126),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_107),
.C(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_104),
.B(n_110),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_131),
.C(n_125),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_120),
.C(n_117),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_134),
.B(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_123),
.B1(n_129),
.B2(n_122),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_118),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_116),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_106),
.C(n_127),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_136),
.Y(n_140)
);


endmodule