module fake_jpeg_9306_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_28),
.B1(n_32),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_24),
.B1(n_37),
.B2(n_34),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_40),
.B1(n_41),
.B2(n_28),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_61),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_22),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_59),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_32),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_47),
.B1(n_45),
.B2(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_70),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_21),
.B1(n_37),
.B2(n_34),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_57),
.B1(n_63),
.B2(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_59),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_51),
.B1(n_63),
.B2(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_16),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_60),
.C(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_53),
.Y(n_137)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_110),
.B(n_118),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_105),
.B1(n_118),
.B2(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_56),
.B1(n_43),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_46),
.B1(n_53),
.B2(n_42),
.Y(n_142)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_114),
.Y(n_147)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_79),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_47),
.B1(n_45),
.B2(n_31),
.Y(n_118)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_122),
.A2(n_148),
.B1(n_25),
.B2(n_29),
.Y(n_181)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_124),
.Y(n_176)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_90),
.B1(n_64),
.B2(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_127),
.A2(n_136),
.B1(n_132),
.B2(n_124),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_132),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_64),
.B(n_97),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_130),
.B(n_133),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_111),
.B(n_94),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_143),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_76),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_67),
.B1(n_71),
.B2(n_81),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_150),
.C(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_69),
.B1(n_68),
.B2(n_46),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_149),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_0),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_38),
.B1(n_42),
.B2(n_31),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_0),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_46),
.B1(n_18),
.B2(n_16),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_84),
.C(n_72),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_160),
.C(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_154),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_1),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_167),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_93),
.C(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_170),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_104),
.B1(n_114),
.B2(n_106),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_171),
.B1(n_91),
.B2(n_80),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_106),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_104),
.B1(n_107),
.B2(n_101),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_178),
.B1(n_121),
.B2(n_139),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_R g174 ( 
.A1(n_137),
.A2(n_29),
.B(n_33),
.C(n_18),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_143),
.A3(n_146),
.B1(n_133),
.B2(n_144),
.C1(n_26),
.C2(n_30),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_19),
.B(n_25),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_131),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_123),
.A2(n_120),
.B(n_26),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_26),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_107),
.C(n_101),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_138),
.C(n_147),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_29),
.B1(n_109),
.B2(n_9),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_191),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_193),
.C(n_199),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_198),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_133),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_204),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_143),
.C(n_139),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_184),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_169),
.B1(n_153),
.B2(n_158),
.Y(n_226)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_109),
.C(n_74),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_207),
.B1(n_212),
.B2(n_183),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_109),
.C(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_208),
.C(n_210),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_R g204 ( 
.A1(n_155),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_179),
.C(n_152),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_228),
.B1(n_237),
.B2(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_227),
.B(n_233),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_173),
.B1(n_152),
.B2(n_171),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_228),
.A2(n_236),
.B1(n_212),
.B2(n_207),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_164),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_164),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_234),
.C(n_237),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_210),
.C(n_189),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_235),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_163),
.B1(n_155),
.B2(n_170),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_163),
.C(n_178),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g251 ( 
.A(n_238),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_196),
.B1(n_187),
.B2(n_185),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_257),
.B(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_201),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_253),
.C(n_254),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_206),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_218),
.C(n_221),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_190),
.C(n_209),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_175),
.C(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_162),
.C(n_211),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_225),
.C(n_253),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_206),
.B(n_2),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_206),
.B1(n_9),
.B2(n_10),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_257),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_266),
.C(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_242),
.C(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_273),
.B1(n_248),
.B2(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_223),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_4),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_264),
.B1(n_246),
.B2(n_271),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_231),
.C(n_224),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_239),
.B(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_1),
.C(n_4),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_4),
.C(n_6),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_240),
.B1(n_244),
.B2(n_249),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_270),
.B1(n_11),
.B2(n_10),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_15),
.B1(n_7),
.B2(n_8),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_284),
.Y(n_290)
);

AOI21x1_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_246),
.B(n_5),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_265),
.B(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_286),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_6),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_9),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_6),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_296),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_263),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_278),
.C(n_285),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_280),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_287),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_277),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_311),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_285),
.B(n_306),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_290),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_290),
.B(n_299),
.C(n_282),
.D(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_315),
.B(n_313),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_316),
.B(n_310),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_314),
.B(n_7),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_8),
.B(n_6),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_7),
.Y(n_322)
);


endmodule