module fake_jpeg_2058_n_511 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_511);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_511;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_59),
.Y(n_153)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g180 ( 
.A(n_60),
.Y(n_180)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_61),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_69),
.Y(n_122)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_65),
.B(n_78),
.Y(n_155)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_27),
.B(n_16),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_77),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_13),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_23),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_102),
.Y(n_167)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_33),
.B(n_13),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_33),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_113),
.Y(n_172)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_32),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_120),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_18),
.Y(n_117)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_35),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_119),
.B(n_28),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_31),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_127),
.B(n_129),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_30),
.B1(n_52),
.B2(n_29),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_149),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_132),
.B(n_145),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_91),
.A2(n_30),
.B1(n_37),
.B2(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_42),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_78),
.A2(n_44),
.B1(n_48),
.B2(n_52),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_65),
.A2(n_20),
.B1(n_47),
.B2(n_43),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_160),
.A2(n_189),
.B1(n_134),
.B2(n_149),
.Y(n_237)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_48),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_164),
.B(n_178),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_57),
.A2(n_18),
.B1(n_41),
.B2(n_29),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_168),
.A2(n_181),
.B1(n_183),
.B2(n_188),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_80),
.B(n_47),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_116),
.B(n_43),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_5),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_41),
.B1(n_28),
.B2(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_103),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_22),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_184),
.B(n_187),
.C(n_173),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_75),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_81),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_87),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_191),
.A2(n_198),
.B1(n_138),
.B2(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_89),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_213),
.Y(n_271)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_205),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_88),
.B1(n_56),
.B2(n_58),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_208),
.B(n_215),
.Y(n_309)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_209),
.Y(n_295)
);

BUFx2_ASAP7_75t_SL g210 ( 
.A(n_166),
.Y(n_210)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_59),
.B1(n_62),
.B2(n_7),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_211),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_10),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_212),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_5),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_166),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_216),
.A2(n_218),
.B1(n_221),
.B2(n_227),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_8),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_217),
.B(n_223),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_155),
.A2(n_8),
.B1(n_10),
.B2(n_194),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_144),
.A2(n_8),
.B1(n_10),
.B2(n_150),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_140),
.Y(n_224)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_122),
.B(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_244),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_143),
.A2(n_176),
.B1(n_180),
.B2(n_151),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_228),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_125),
.B(n_142),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_237),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_123),
.B(n_131),
.Y(n_232)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_124),
.Y(n_235)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_235),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_180),
.A2(n_169),
.B1(n_174),
.B2(n_133),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_236),
.A2(n_252),
.B1(n_263),
.B2(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_156),
.Y(n_241)
);

INVx11_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_139),
.B(n_147),
.Y(n_242)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_243),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_148),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_245),
.Y(n_289)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_251),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_181),
.A2(n_130),
.B(n_189),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_249),
.A2(n_262),
.B(n_261),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_171),
.B(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_254),
.B(n_255),
.Y(n_310)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_128),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_138),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_259),
.B1(n_265),
.B2(n_266),
.Y(n_277)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_257),
.B(n_258),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_135),
.B(n_165),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_124),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_268),
.Y(n_279)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_154),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_185),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_186),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_121),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_157),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_254),
.B1(n_239),
.B2(n_203),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_196),
.A2(n_152),
.B1(n_153),
.B2(n_165),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_214),
.B1(n_229),
.B2(n_213),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_197),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_256),
.B1(n_235),
.B2(n_255),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_244),
.A2(n_152),
.B1(n_170),
.B2(n_249),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_280),
.A2(n_288),
.B1(n_285),
.B2(n_303),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_284),
.Y(n_333)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_247),
.A2(n_253),
.B1(n_231),
.B2(n_204),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_291),
.A2(n_298),
.B1(n_307),
.B2(n_315),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_292),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_238),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_296),
.C(n_300),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_212),
.B(n_230),
.C(n_225),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_246),
.A2(n_250),
.B1(n_256),
.B2(n_258),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_230),
.B(n_219),
.C(n_207),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_212),
.A2(n_220),
.B(n_228),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_302),
.A2(n_306),
.B(n_290),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_224),
.B(n_248),
.C(n_266),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_282),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_260),
.A2(n_240),
.B1(n_234),
.B2(n_257),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_245),
.A2(n_205),
.B1(n_209),
.B2(n_243),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_291),
.A2(n_233),
.B1(n_265),
.B2(n_259),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_329),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_274),
.A2(n_222),
.B1(n_293),
.B2(n_288),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_294),
.B(n_293),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_339),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_280),
.A2(n_274),
.B1(n_303),
.B2(n_272),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_325),
.A2(n_345),
.B1(n_349),
.B2(n_356),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_274),
.A2(n_278),
.B1(n_301),
.B2(n_318),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_327),
.B(n_330),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_271),
.A2(n_306),
.B1(n_313),
.B2(n_279),
.Y(n_329)
);

AOI22x1_ASAP7_75t_L g330 ( 
.A1(n_299),
.A2(n_271),
.B1(n_313),
.B2(n_310),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_331),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_286),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_344),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_284),
.A2(n_299),
.B1(n_296),
.B2(n_316),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_334),
.A2(n_336),
.B1(n_358),
.B2(n_328),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_309),
.A2(n_289),
.B1(n_302),
.B2(n_295),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_335),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_315),
.A2(n_283),
.B1(n_320),
.B2(n_311),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_277),
.A2(n_283),
.B(n_300),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_341),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_340),
.A2(n_325),
.B(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_281),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_319),
.B1(n_312),
.B2(n_297),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_273),
.B(n_286),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_352),
.Y(n_374)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_275),
.B(n_308),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_351),
.C(n_342),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_308),
.A2(n_317),
.B1(n_305),
.B2(n_277),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_276),
.B(n_277),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_314),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_332),
.Y(n_362)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_355),
.B(n_337),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_280),
.B1(n_291),
.B2(n_274),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_291),
.A2(n_274),
.B1(n_293),
.B2(n_288),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_337),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_361),
.A2(n_386),
.B(n_363),
.Y(n_399)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_345),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_372),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_331),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_365),
.B(n_366),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_324),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_339),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_384),
.C(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_371),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_344),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_373),
.B(n_377),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_341),
.B(n_329),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_383),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_356),
.A2(n_323),
.B1(n_353),
.B2(n_328),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_385),
.A2(n_336),
.B1(n_348),
.B2(n_338),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_340),
.A2(n_358),
.B(n_330),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_330),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_398),
.C(n_400),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_369),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_390),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_369),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_360),
.A2(n_335),
.B1(n_328),
.B2(n_349),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_387),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_381),
.A2(n_357),
.B1(n_321),
.B2(n_326),
.Y(n_394)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_394),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_371),
.A2(n_354),
.B(n_326),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_395),
.A2(n_399),
.B(n_380),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_396),
.A2(n_406),
.B1(n_375),
.B2(n_361),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_347),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_365),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g401 ( 
.A(n_359),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_401),
.B(n_410),
.Y(n_430)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_374),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_408),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_383),
.B1(n_379),
.B2(n_387),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_384),
.C(n_380),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_359),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_411),
.Y(n_418)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_413),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_419),
.A2(n_426),
.B1(n_414),
.B2(n_392),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_433),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_388),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_427),
.Y(n_447)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_406),
.A2(n_392),
.B1(n_386),
.B2(n_414),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_376),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_395),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_428),
.Y(n_448)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_411),
.Y(n_433)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_399),
.B(n_376),
.CI(n_372),
.CON(n_434),
.SN(n_434)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_434),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_376),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_407),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_389),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_436),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_412),
.C(n_397),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_438),
.A2(n_439),
.B1(n_446),
.B2(n_449),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_405),
.B1(n_404),
.B2(n_391),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_432),
.B1(n_390),
.B2(n_416),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_441),
.A2(n_453),
.B1(n_418),
.B2(n_422),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_437),
.C(n_420),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_424),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_430),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_391),
.B1(n_393),
.B2(n_396),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_432),
.A2(n_426),
.B1(n_394),
.B2(n_375),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_452),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_427),
.B(n_397),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_435),
.A2(n_364),
.B1(n_413),
.B2(n_378),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_456),
.B(n_460),
.Y(n_472)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_457),
.A2(n_459),
.B1(n_463),
.B2(n_444),
.Y(n_477)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_423),
.C(n_420),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_450),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_439),
.A2(n_421),
.B(n_434),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_466),
.Y(n_475)
);

INVx11_ASAP7_75t_L g463 ( 
.A(n_454),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_434),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_467),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_443),
.A2(n_422),
.B1(n_429),
.B2(n_425),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_418),
.Y(n_467)
);

XNOR2x1_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_453),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_431),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_455),
.Y(n_480)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_456),
.B(n_442),
.CI(n_441),
.CON(n_471),
.SN(n_471)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_471),
.A2(n_478),
.B1(n_468),
.B2(n_438),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_480),
.Y(n_482)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_466),
.Y(n_474)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_469),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_479),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_458),
.A2(n_445),
.B1(n_451),
.B2(n_449),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_464),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_SL g481 ( 
.A1(n_474),
.A2(n_451),
.B1(n_458),
.B2(n_455),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_486),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_471),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_485),
.A2(n_489),
.B(n_446),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_462),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_464),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_475),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_460),
.B(n_467),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_461),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_491),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_488),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_496),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_473),
.C(n_475),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_494),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_457),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_501),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_487),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_459),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_504),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_499),
.B(n_493),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_500),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_497),
.B(n_482),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_505),
.C(n_486),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_481),
.C(n_444),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_417),
.C(n_433),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_510),
.Y(n_511)
);


endmodule