module fake_jpeg_182_n_87 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_87);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_40),
.B1(n_0),
.B2(n_1),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_37),
.B(n_36),
.C(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_50),
.B1(n_38),
.B2(n_43),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_27),
.B(n_30),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_10),
.A3(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_60),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_57),
.B1(n_55),
.B2(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_23),
.C(n_17),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_16),
.C(n_15),
.Y(n_65)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_69),
.C(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_3),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_14),
.C(n_12),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_11),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_77),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_1),
.C(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_73),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_75),
.C(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_79),
.B1(n_78),
.B2(n_6),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_4),
.B(n_5),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_4),
.B(n_6),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_8),
.Y(n_87)
);


endmodule