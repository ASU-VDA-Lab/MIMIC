module fake_jpeg_16196_n_62 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_19),
.A2(n_7),
.B1(n_18),
.B2(n_26),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_19),
.A2(n_26),
.B1(n_25),
.B2(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_27),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_21),
.B1(n_36),
.B2(n_37),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_33),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_34),
.B1(n_19),
.B2(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_50),
.B1(n_40),
.B2(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_42),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_50),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_48),
.B(n_45),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_47),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_23),
.B(n_46),
.Y(n_62)
);


endmodule