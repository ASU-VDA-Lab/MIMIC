module fake_jpeg_17416_n_303 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_36),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_28),
.B1(n_33),
.B2(n_27),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_51),
.B(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_31),
.B1(n_23),
.B2(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_55),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_13),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_23),
.B1(n_15),
.B2(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_69),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_20),
.B(n_29),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_20),
.C(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_44),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_23),
.B1(n_32),
.B2(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_37),
.B1(n_17),
.B2(n_14),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_45),
.C(n_44),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_13),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_46),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_53),
.B1(n_51),
.B2(n_50),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_99),
.B(n_106),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_73),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_101),
.B(n_89),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_82),
.B1(n_77),
.B2(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_100),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_58),
.B1(n_63),
.B2(n_68),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NAND2x1_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_57),
.B1(n_46),
.B2(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_113),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_119),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_89),
.B(n_79),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_102),
.Y(n_142)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_130),
.Y(n_148)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_79),
.B(n_76),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_108),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_93),
.B(n_101),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_72),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_127),
.B(n_81),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_98),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_80),
.C(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_70),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_76),
.C(n_111),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_157),
.C(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_79),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_90),
.C(n_93),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_109),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_161),
.C(n_20),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_109),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_87),
.Y(n_179)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_178),
.B(n_25),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_128),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_155),
.B(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_122),
.B1(n_132),
.B2(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_182),
.Y(n_190)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_119),
.B(n_125),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_115),
.B1(n_119),
.B2(n_122),
.Y(n_180)
);

AOI22x1_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_115),
.B1(n_120),
.B2(n_113),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_84),
.B1(n_86),
.B2(n_79),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_20),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_69),
.B1(n_59),
.B2(n_25),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_142),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_12),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_11),
.C(n_10),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_39),
.C(n_48),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_147),
.C(n_148),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_193),
.C(n_201),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_204),
.B(n_164),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_195),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_183),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_18),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_148),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_159),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_210),
.C(n_185),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_166),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_170),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_199),
.A2(n_196),
.B1(n_178),
.B2(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_216),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_224),
.B(n_210),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_176),
.B1(n_173),
.B2(n_163),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_217),
.B(n_11),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_228),
.C(n_230),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_184),
.B1(n_186),
.B2(n_177),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_224),
.B1(n_227),
.B2(n_214),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_11),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_180),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

FAx1_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_180),
.CI(n_164),
.CON(n_227),
.SN(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_21),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_167),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_180),
.B1(n_175),
.B2(n_188),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_189),
.B1(n_208),
.B2(n_15),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_193),
.B1(n_198),
.B2(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_246),
.B1(n_234),
.B2(n_232),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_234),
.B(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_9),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_227),
.A2(n_22),
.B(n_24),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_221),
.C(n_235),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_223),
.B(n_219),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_39),
.C(n_48),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_220),
.C(n_228),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_251),
.C(n_259),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_220),
.B1(n_15),
.B2(n_24),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_261),
.C(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_48),
.C(n_43),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_21),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_21),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_9),
.C(n_2),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_245),
.B(n_256),
.C(n_24),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_48),
.C(n_43),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_270),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_267),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_247),
.C(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_238),
.B(n_246),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_21),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_272),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_21),
.C(n_43),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_43),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_257),
.B(n_260),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_0),
.CI(n_3),
.CON(n_279),
.SN(n_279)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_280),
.C(n_283),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_39),
.C(n_20),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_22),
.B(n_39),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_20),
.C(n_22),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_263),
.C(n_20),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_287),
.C(n_289),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_3),
.C(n_4),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_279),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_277),
.B1(n_276),
.B2(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_3),
.C(n_4),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_278),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_286),
.B(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_293),
.C(n_5),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_4),
.B(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_295),
.C(n_5),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_4),
.C(n_5),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_6),
.C(n_7),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_7),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_7),
.C(n_296),
.Y(n_303)
);


endmodule