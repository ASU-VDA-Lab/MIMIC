module fake_jpeg_29227_n_492 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_492);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_492;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_8),
.B(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_62),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_64),
.B(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_69),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_14),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_32),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_84),
.B(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_13),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_23),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_93),
.B1(n_21),
.B2(n_40),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_98),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_28),
.B(n_13),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_44),
.A3(n_24),
.B1(n_39),
.B2(n_33),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_109),
.A2(n_144),
.B(n_45),
.C(n_29),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_39),
.B1(n_24),
.B2(n_22),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_110),
.A2(n_126),
.B1(n_133),
.B2(n_142),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_39),
.B1(n_33),
.B2(n_42),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_45),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_33),
.B1(n_37),
.B2(n_30),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_73),
.B1(n_76),
.B2(n_52),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_28),
.B1(n_23),
.B2(n_42),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_130),
.B1(n_137),
.B2(n_45),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_18),
.B1(n_40),
.B2(n_21),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_50),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_35),
.B1(n_34),
.B2(n_42),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_18),
.B1(n_40),
.B2(n_21),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_59),
.A2(n_35),
.B1(n_34),
.B2(n_42),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_50),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_91),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_66),
.A2(n_30),
.B(n_26),
.C(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_68),
.B(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_70),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_49),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_199),
.B(n_170),
.Y(n_213)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_61),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_51),
.B(n_64),
.C(n_74),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_53),
.B(n_86),
.C(n_55),
.Y(n_237)
);

OR2x2_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_81),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_196),
.C(n_131),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_38),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_170),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_90),
.Y(n_171)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_80),
.B1(n_78),
.B2(n_65),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_174),
.B1(n_189),
.B2(n_151),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_86),
.B(n_30),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_176),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_116),
.A2(n_67),
.B1(n_94),
.B2(n_89),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_38),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_181),
.Y(n_203)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_104),
.B(n_26),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_200),
.B1(n_125),
.B2(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_115),
.B(n_31),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_187),
.Y(n_219)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_195),
.B(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_192),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_97),
.B(n_54),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_77),
.B(n_72),
.Y(n_221)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_194),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_27),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_101),
.B(n_67),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_176),
.B(n_160),
.Y(n_207)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_139),
.B(n_86),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_113),
.A2(n_71),
.B1(n_83),
.B2(n_29),
.Y(n_200)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_202),
.B1(n_99),
.B2(n_153),
.Y(n_243)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_204),
.A2(n_220),
.B1(n_222),
.B2(n_200),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_209),
.B1(n_214),
.B2(n_216),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_55),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_162),
.A2(n_124),
.B1(n_113),
.B2(n_143),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_227),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_164),
.A2(n_124),
.B1(n_143),
.B2(n_125),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_103),
.B1(n_105),
.B2(n_134),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_169),
.B1(n_167),
.B2(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_217),
.A2(n_218),
.B1(n_225),
.B2(n_231),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_159),
.A2(n_103),
.B1(n_105),
.B2(n_134),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_112),
.B1(n_107),
.B2(n_145),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_191),
.B(n_196),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_172),
.A2(n_112),
.B1(n_131),
.B2(n_114),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_167),
.A2(n_81),
.B1(n_34),
.B2(n_35),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_114),
.B1(n_75),
.B2(n_79),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_237),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_160),
.A2(n_153),
.B1(n_106),
.B2(n_146),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_238),
.A2(n_244),
.B1(n_99),
.B2(n_179),
.Y(n_276)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_106),
.B1(n_60),
.B2(n_147),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_168),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_259),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_154),
.B(n_165),
.C(n_175),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_248),
.A2(n_282),
.B(n_246),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_249),
.A2(n_272),
.B(n_212),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_199),
.C(n_166),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_255),
.C(n_215),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_190),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_283),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_253),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_188),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_254),
.B(n_256),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_184),
.C(n_193),
.Y(n_255)
);

OAI32xp33_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_200),
.A3(n_174),
.B1(n_177),
.B2(n_161),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_188),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_258),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_226),
.B(n_201),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_261),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_178),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_265),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_223),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_229),
.B(n_186),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_267),
.Y(n_313)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_274),
.B1(n_206),
.B2(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

AO21x2_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_200),
.B(n_155),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_SL g274 ( 
.A1(n_221),
.A2(n_180),
.B(n_202),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_220),
.B1(n_204),
.B2(n_222),
.Y(n_291)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_281),
.A2(n_284),
.B1(n_212),
.B2(n_236),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_228),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_238),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_302),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_205),
.C(n_215),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_294),
.C(n_299),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_306),
.B1(n_272),
.B2(n_277),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_205),
.C(n_215),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_296),
.A2(n_307),
.B1(n_319),
.B2(n_155),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_298),
.B(n_240),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_210),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_314),
.B(n_267),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_210),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_228),
.C(n_232),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_318),
.C(n_321),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_277),
.A2(n_219),
.B1(n_231),
.B2(n_213),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_266),
.B1(n_268),
.B2(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_282),
.A2(n_237),
.B(n_203),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_264),
.B(n_276),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_251),
.A2(n_232),
.B(n_203),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_260),
.A2(n_243),
.B(n_223),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_316),
.A2(n_121),
.B(n_48),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_209),
.C(n_214),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_266),
.A2(n_218),
.B1(n_216),
.B2(n_225),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_236),
.C(n_240),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_249),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_331),
.C(n_344),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_323),
.A2(n_325),
.B1(n_335),
.B2(n_297),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_324),
.A2(n_326),
.B(n_333),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_268),
.B1(n_272),
.B2(n_247),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_303),
.A2(n_272),
.B1(n_248),
.B2(n_269),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_328),
.B(n_349),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_271),
.Y(n_329)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_247),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_298),
.B(n_229),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_332),
.B(n_295),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_306),
.A2(n_272),
.B1(n_279),
.B2(n_278),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_272),
.A3(n_281),
.B1(n_275),
.B2(n_253),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_345),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_252),
.B1(n_261),
.B2(n_259),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_280),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_263),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_305),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_245),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_342),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_245),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_317),
.B1(n_315),
.B2(n_308),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_234),
.C(n_195),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_300),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g346 ( 
.A1(n_307),
.A2(n_192),
.A3(n_234),
.B1(n_29),
.B2(n_48),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_257),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_241),
.C(n_239),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_352),
.C(n_344),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_321),
.B(n_48),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_353),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_311),
.A2(n_198),
.B(n_188),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_350),
.A2(n_288),
.B1(n_315),
.B2(n_308),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g378 ( 
.A(n_351),
.B(n_292),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_294),
.B(n_239),
.C(n_257),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_288),
.B(n_316),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_SL g355 ( 
.A1(n_324),
.A2(n_296),
.B(n_319),
.C(n_318),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_355),
.A2(n_0),
.B(n_1),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_337),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_369),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_330),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_346),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_361),
.A2(n_382),
.B1(n_333),
.B2(n_340),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_363),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_304),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_366),
.B(n_375),
.Y(n_389)
);

AO22x1_ASAP7_75t_SL g367 ( 
.A1(n_327),
.A2(n_317),
.B1(n_293),
.B2(n_285),
.Y(n_367)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_332),
.A2(n_293),
.B1(n_314),
.B2(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_312),
.B1(n_285),
.B2(n_287),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_372),
.B(n_329),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_379),
.C(n_338),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_330),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_325),
.A2(n_287),
.B1(n_297),
.B2(n_292),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_339),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_378),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_331),
.B(n_295),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_350),
.B1(n_343),
.B2(n_354),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_353),
.B(n_326),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_371),
.B(n_377),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_345),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_385),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_386),
.A2(n_397),
.B1(n_404),
.B2(n_400),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_357),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_391),
.B1(n_392),
.B2(n_359),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_399),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_383),
.A2(n_335),
.B1(n_341),
.B2(n_334),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_383),
.A2(n_365),
.B1(n_382),
.B2(n_361),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_338),
.C(n_347),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_393),
.B(n_394),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_380),
.B(n_352),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_354),
.B1(n_351),
.B2(n_348),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_328),
.C(n_349),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_408),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_403),
.B(n_395),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_364),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_0),
.C(n_2),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_402),
.A2(n_371),
.B1(n_364),
.B2(n_362),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_409),
.A2(n_422),
.B1(n_395),
.B2(n_405),
.Y(n_439)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_411),
.Y(n_430)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_391),
.A2(n_378),
.B(n_355),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_416),
.B(n_428),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_355),
.B(n_380),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_419),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_357),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_406),
.B1(n_407),
.B2(n_388),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_424),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_374),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_426),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_379),
.Y(n_426)
);

A2O1A1O1Ixp25_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_356),
.B(n_355),
.C(n_358),
.D(n_360),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_403),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_367),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_417),
.B(n_390),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_432),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_433),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_389),
.C(n_398),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_437),
.C(n_410),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_408),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_440),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_389),
.C(n_397),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_356),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_409),
.A2(n_395),
.B(n_405),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_443),
.A2(n_413),
.B(n_416),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_453),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_455),
.B(n_443),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_430),
.A2(n_422),
.B1(n_411),
.B2(n_421),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

INVx11_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_439),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_418),
.C(n_427),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_451),
.C(n_454),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_386),
.C(n_415),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_412),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_441),
.A2(n_425),
.B(n_414),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_441),
.A2(n_444),
.B1(n_430),
.B2(n_442),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_453),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_414),
.C(n_355),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_458),
.B(n_450),
.C(n_447),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_446),
.A2(n_431),
.B(n_429),
.Y(n_460)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_460),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_461),
.B(n_463),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_458),
.C(n_451),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_465),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_452),
.B(n_456),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_469),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_457),
.A2(n_431),
.B(n_438),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_10),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_10),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_SL g471 ( 
.A1(n_463),
.A2(n_367),
.B(n_448),
.C(n_444),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g480 ( 
.A1(n_471),
.A2(n_462),
.B(n_459),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_468),
.A2(n_449),
.B1(n_404),
.B2(n_11),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_475),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_2),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_2),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_479),
.A2(n_459),
.B(n_3),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_L g486 ( 
.A1(n_480),
.A2(n_482),
.B(n_473),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_481),
.A2(n_483),
.B(n_479),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_464),
.C(n_3),
.Y(n_483)
);

OAI221xp5_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_486),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_488)
);

AOI321xp33_ASAP7_75t_L g487 ( 
.A1(n_484),
.A2(n_473),
.A3(n_478),
.B1(n_476),
.B2(n_464),
.C(n_6),
.Y(n_487)
);

AOI321xp33_ASAP7_75t_L g489 ( 
.A1(n_487),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_489)
);

OAI321xp33_ASAP7_75t_L g490 ( 
.A1(n_488),
.A2(n_489),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_490),
.A2(n_6),
.B(n_7),
.Y(n_491)
);

FAx1_ASAP7_75t_SL g492 ( 
.A(n_491),
.B(n_6),
.CI(n_345),
.CON(n_492),
.SN(n_492)
);


endmodule