module fake_jpeg_8219_n_247 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_15),
.B1(n_23),
.B2(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_43),
.B1(n_54),
.B2(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_15),
.B1(n_23),
.B2(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_15),
.B(n_38),
.C(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_15),
.B1(n_28),
.B2(n_14),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_25),
.B1(n_14),
.B2(n_28),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_38),
.B(n_19),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_19),
.C(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_66),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_38),
.B1(n_26),
.B2(n_16),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_68),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_37),
.B(n_30),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_64),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_61),
.B(n_59),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_93),
.C(n_77),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.C(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_61),
.C(n_67),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_105),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_30),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_71),
.C(n_58),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_76),
.C(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_75),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_66),
.B1(n_64),
.B2(n_33),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_64),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_66),
.B1(n_33),
.B2(n_41),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_56),
.B1(n_46),
.B2(n_75),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_84),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_85),
.B(n_89),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_121),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_89),
.B(n_85),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_123),
.B(n_132),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_87),
.C(n_74),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_27),
.B(n_14),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_126),
.B(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_65),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_97),
.C(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_65),
.B(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_124),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_139),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_154),
.Y(n_173)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_103),
.B1(n_100),
.B2(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_141),
.B1(n_151),
.B2(n_153),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_125),
.B1(n_133),
.B2(n_134),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_106),
.B(n_63),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_149),
.B(n_17),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_29),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_1),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_88),
.B1(n_60),
.B2(n_46),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_88),
.B1(n_63),
.B2(n_60),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_88),
.C(n_34),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_153),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_160),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_161),
.B1(n_171),
.B2(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_153),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_121),
.B1(n_130),
.B2(n_129),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_136),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_56),
.B1(n_28),
.B2(n_25),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_25),
.B1(n_27),
.B2(n_63),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_20),
.B1(n_24),
.B2(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_138),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_182),
.C(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_135),
.C(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_188),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_145),
.B1(n_149),
.B2(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_149),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_145),
.C(n_34),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_169),
.B(n_160),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_196),
.B(n_198),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_162),
.B(n_157),
.Y(n_196)
);

AO221x1_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_158),
.B1(n_24),
.B2(n_20),
.C(n_22),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_21),
.B(n_30),
.C(n_29),
.D(n_34),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_201),
.B(n_176),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_187),
.A2(n_1),
.B(n_2),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_203),
.A2(n_183),
.B(n_179),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_29),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_191),
.C(n_202),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_213),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_182),
.C(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_215),
.C(n_216),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_214),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_203),
.B(n_197),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_199),
.B(n_24),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_8),
.C(n_13),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_17),
.C(n_20),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_193),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_2),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_207),
.A2(n_193),
.B(n_206),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_10),
.B(n_2),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_216),
.A2(n_200),
.B1(n_7),
.B2(n_9),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_223),
.A2(n_225),
.B1(n_10),
.B2(n_2),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_12),
.C(n_11),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_1),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_17),
.B1(n_12),
.B2(n_11),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_233),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_226),
.B1(n_4),
.B2(n_5),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_3),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_232),
.B(n_220),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_3),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_241),
.B1(n_238),
.B2(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_235),
.B(n_229),
.Y(n_241)
);

OAI21x1_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_236),
.B(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_243),
.C2(n_242),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_6),
.Y(n_247)
);


endmodule