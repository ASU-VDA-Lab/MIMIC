module fake_jpeg_24592_n_25 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_17;
wire n_15;

INVx11_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.C(n_14),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B1(n_13),
.B2(n_2),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_2),
.Y(n_21)
);

AOI31xp67_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_22),
.A3(n_4),
.B(n_5),
.Y(n_24)
);

OAI321xp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_3),
.A3(n_6),
.B1(n_7),
.B2(n_10),
.C(n_12),
.Y(n_25)
);


endmodule