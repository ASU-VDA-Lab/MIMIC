module real_jpeg_9543_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_0),
.A2(n_1),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_0),
.A2(n_26),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_1),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_21),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_42),
.B1(n_45),
.B2(n_51),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_9),
.B(n_42),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_6),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_24),
.B(n_30),
.C(n_34),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_5),
.B(n_24),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_6),
.A3(n_24),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_6),
.B(n_51),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_9),
.B1(n_27),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_10),
.B1(n_32),
.B2(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_8),
.B1(n_32),
.B2(n_48),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_27),
.B(n_51),
.C(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

HAxp5_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_27),
.CON(n_26),
.SN(n_26)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_24),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_24),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_27),
.B1(n_42),
.B2(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_9),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_30),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_10),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_86),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_84),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_72),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_14),
.B(n_72),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_56),
.C(n_64),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_15),
.B(n_56),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_39),
.B2(n_55),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_16),
.A2(n_17),
.B1(n_99),
.B2(n_104),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_16),
.A2(n_17),
.B1(n_65),
.B2(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_18),
.A2(n_37),
.B1(n_57),
.B2(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_18),
.A2(n_37),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_23),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_25),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_27),
.B(n_53),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_27),
.B(n_43),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_28),
.A2(n_79),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_79),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_28),
.A2(n_38),
.B1(n_49),
.B2(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_103),
.C(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_28),
.A2(n_38),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_31),
.B(n_32),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_36),
.Y(n_148)
);

AOI211xp5_ASAP7_75t_SL g92 ( 
.A1(n_37),
.A2(n_49),
.B(n_71),
.C(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_94),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_38),
.A2(n_94),
.B(n_151),
.C(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_39),
.A2(n_68),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_49),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_40),
.A2(n_49),
.B1(n_94),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_41),
.A2(n_43),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_45),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_66),
.B1(n_94),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_49),
.A2(n_94),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_49),
.A2(n_94),
.B1(n_125),
.B2(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_49),
.B(n_103),
.C(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_49),
.A2(n_94),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_157),
.C(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_54),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_53),
.B1(n_62),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_64),
.B(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_68),
.B(n_70),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_65),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_69),
.A2(n_71),
.B(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_82),
.B2(n_83),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_186),
.B(n_190),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_118),
.B(n_174),
.C(n_185),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_105),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_89),
.B(n_105),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_91),
.B(n_96),
.C(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_103),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_112),
.B1(n_128),
.B2(n_131),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_112),
.B1(n_147),
.B2(n_150),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_103),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_103),
.B(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_114),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_106),
.A2(n_107),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_109),
.B1(n_146),
.B2(n_151),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_140),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_173),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_166),
.B(n_172),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_153),
.B(n_165),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_143),
.B(n_152),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_132),
.B(n_142),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_127),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_147),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_156),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_176),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_183),
.C(n_184),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);


endmodule