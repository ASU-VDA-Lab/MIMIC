module fake_ariane_2399_n_1883 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1883);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1883;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_104),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_34),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_2),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_90),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_39),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_81),
.Y(n_199)
);

BUFx8_ASAP7_75t_SL g200 ( 
.A(n_32),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_4),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_32),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_113),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_83),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_103),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_35),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_66),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_12),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_38),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_33),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_136),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_7),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_51),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_33),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_38),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_8),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_42),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_74),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_111),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_85),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_40),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_124),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_150),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_66),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_72),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_21),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_126),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_152),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_47),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_78),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_172),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_98),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_40),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_12),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_30),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_123),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_39),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_36),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_108),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_16),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_17),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_88),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_143),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_0),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_169),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_158),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_50),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_87),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_47),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_118),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_131),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_95),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_106),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_30),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_101),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_162),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_77),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_37),
.Y(n_283)
);

BUFx2_ASAP7_75t_SL g284 ( 
.A(n_122),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_34),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_107),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_89),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_159),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_105),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_164),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_25),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_19),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_84),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_43),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_112),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_24),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_99),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_138),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_154),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_116),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_160),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_42),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_26),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_91),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_135),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_167),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_20),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_53),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_46),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_27),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_109),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_45),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_173),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_63),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_49),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_48),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_61),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_4),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_10),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_5),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_63),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_64),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_114),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_110),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_56),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_146),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_23),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_14),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_144),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_139),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_9),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_68),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_117),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_56),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_59),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_11),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_48),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_76),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_100),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_168),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_45),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_43),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_171),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_51),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_35),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_11),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_141),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_67),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_79),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_44),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_54),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_200),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_213),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_237),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_0),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_259),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_291),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_301),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_309),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_344),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_213),
.B(n_269),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_213),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_287),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_191),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_213),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_209),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_213),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_221),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_191),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_249),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_213),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_213),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_213),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_182),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_182),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_303),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_186),
.B(n_1),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_182),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_270),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_188),
.B(n_1),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_238),
.B(n_2),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_182),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_182),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_193),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_211),
.B(n_129),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_222),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_226),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_231),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_222),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_222),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_287),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_222),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_222),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_197),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_285),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_285),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_280),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_285),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_314),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_250),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_314),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_314),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_285),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_285),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_253),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_229),
.B(n_3),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_235),
.B(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_254),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_212),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_212),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_256),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_261),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_302),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_214),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_302),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_197),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_197),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_332),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_268),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_214),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_272),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_217),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_217),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_192),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_274),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_192),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_185),
.B(n_5),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_193),
.B(n_6),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_278),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_198),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_220),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_283),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_220),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_295),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_361),
.B(n_284),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_187),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_239),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_440),
.A2(n_356),
.B1(n_311),
.B2(n_349),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_245),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_248),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_369),
.B(n_289),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_369),
.B(n_230),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_370),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_377),
.B(n_251),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_377),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_383),
.B(n_252),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_385),
.B(n_257),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_386),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_376),
.B(n_292),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_203),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_398),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_363),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_372),
.B(n_266),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

CKINVDCx8_ASAP7_75t_R g489 ( 
.A(n_357),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_425),
.B(n_198),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_372),
.B(n_271),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

CKINVDCx6p67_ASAP7_75t_R g500 ( 
.A(n_411),
.Y(n_500)
);

CKINVDCx8_ASAP7_75t_R g501 ( 
.A(n_358),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_378),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_273),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_403),
.B(n_276),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_436),
.B(n_288),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_361),
.B(n_295),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_436),
.B(n_234),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_438),
.B(n_308),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_382),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_446),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_445),
.B(n_327),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_422),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_422),
.B(n_328),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_524),
.B(n_400),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_457),
.B(n_373),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_459),
.B(n_234),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_449),
.A2(n_457),
.B1(n_459),
.B2(n_510),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_449),
.A2(n_389),
.B1(n_419),
.B2(n_368),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_452),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_455),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_524),
.B(n_412),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_472),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_475),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_524),
.B(n_417),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_464),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_449),
.B(n_392),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_449),
.A2(n_392),
.B1(n_418),
.B2(n_355),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_388),
.Y(n_542)
);

AO21x2_ASAP7_75t_L g543 ( 
.A1(n_463),
.A2(n_418),
.B(n_342),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_524),
.B(n_420),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_472),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_449),
.A2(n_439),
.B1(n_442),
.B2(n_396),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_464),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_455),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_475),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_511),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_455),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_449),
.A2(n_439),
.B1(n_380),
.B2(n_393),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_510),
.A2(n_393),
.B1(n_427),
.B2(n_315),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_464),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_502),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_473),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_473),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_502),
.B(n_448),
.Y(n_562)
);

AO22x1_ASAP7_75t_L g563 ( 
.A1(n_450),
.A2(n_406),
.B1(n_201),
.B2(n_205),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_476),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_447),
.B(n_424),
.C(n_423),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_477),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_464),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_447),
.B(n_431),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_501),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_502),
.B(n_433),
.Y(n_570)
);

AND3x1_ASAP7_75t_L g571 ( 
.A(n_453),
.B(n_223),
.C(n_218),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_448),
.B(n_437),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_478),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_475),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_478),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_503),
.B(n_441),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_464),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_490),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_479),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_468),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_490),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_503),
.B(n_444),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_458),
.B(n_379),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_458),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_486),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_479),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_513),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_468),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_485),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_460),
.B(n_462),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_451),
.B(n_413),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_453),
.A2(n_440),
.B1(n_355),
.B2(n_350),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_495),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_486),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_495),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_450),
.B(n_234),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_450),
.B(n_360),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_460),
.B(n_282),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_493),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_462),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_511),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_495),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_481),
.A2(n_205),
.B1(n_201),
.B2(n_336),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_466),
.B(n_179),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_481),
.B(n_234),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_500),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_468),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_468),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_495),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_468),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_466),
.B(n_179),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_481),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_489),
.B(n_362),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_501),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_468),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_501),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_468),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_461),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_491),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_474),
.B(n_234),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_467),
.B(n_299),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_461),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_461),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_461),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_491),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_480),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_508),
.B(n_432),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_492),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_489),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_489),
.B(n_180),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_487),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_467),
.B(n_299),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_492),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_497),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_500),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_470),
.B(n_180),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_480),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_515),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_520),
.A2(n_244),
.B1(n_225),
.B2(n_353),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_497),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_498),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_498),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_508),
.B(n_432),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_515),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_470),
.B(n_181),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_451),
.B(n_414),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_SL g658 ( 
.A(n_463),
.B(n_397),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_454),
.B(n_181),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_454),
.B(n_183),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_505),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_480),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_487),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_505),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_515),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_515),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_500),
.B(n_336),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_515),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_520),
.A2(n_346),
.B1(n_322),
.B2(n_313),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_518),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_456),
.B(n_183),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_518),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_R g674 ( 
.A(n_496),
.B(n_364),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_518),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_496),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_504),
.B(n_338),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_592),
.B(n_428),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_592),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_456),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_642),
.B(n_504),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_591),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_594),
.B(n_429),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_664),
.B(n_506),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_608),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_664),
.B(n_506),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_608),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_527),
.A2(n_469),
.B1(n_465),
.B2(n_517),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_529),
.B(n_465),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_630),
.A2(n_509),
.B1(n_516),
.B2(n_514),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_535),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_604),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_569),
.B(n_365),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_570),
.B(n_661),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_598),
.B(n_469),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_535),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_626),
.A2(n_635),
.B(n_632),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_657),
.B(n_542),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_572),
.B(n_514),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_554),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_540),
.A2(n_630),
.B1(n_539),
.B2(n_620),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_603),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_601),
.B(n_184),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_597),
.A2(n_258),
.B(n_233),
.C(n_241),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_557),
.B(n_184),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_620),
.B(n_517),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_548),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_563),
.B(n_265),
.C(n_260),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_SL g710 ( 
.A(n_525),
.B(n_339),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_563),
.B(n_293),
.C(n_277),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_548),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_677),
.B(n_660),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_601),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_630),
.B(n_518),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_606),
.B(n_522),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_638),
.B(n_522),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_638),
.B(n_509),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_559),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_633),
.B(n_518),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_559),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_677),
.B(n_672),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_560),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_633),
.B(n_512),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_560),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_632),
.B(n_509),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_601),
.B(n_189),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_561),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_633),
.B(n_512),
.Y(n_729)
);

NAND3x1_ASAP7_75t_L g730 ( 
.A(n_599),
.B(n_381),
.C(n_375),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_561),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_564),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_539),
.A2(n_516),
.B1(n_518),
.B2(n_521),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_601),
.B(n_430),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_565),
.B(n_189),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_638),
.B(n_516),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_633),
.B(n_518),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_564),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_640),
.B(n_549),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_629),
.B(n_519),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_539),
.A2(n_243),
.B1(n_230),
.B2(n_246),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_566),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_539),
.A2(n_345),
.B1(n_340),
.B2(n_348),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_637),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_532),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_668),
.B(n_366),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_566),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_638),
.B(n_521),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_532),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_638),
.B(n_521),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_637),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_SL g753 ( 
.A1(n_599),
.A2(n_409),
.B1(n_391),
.B2(n_367),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_573),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_654),
.B(n_519),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_523),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_648),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_573),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_569),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_574),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_654),
.B(n_523),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_622),
.B(n_624),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_654),
.B(n_190),
.Y(n_763)
);

NAND2x1_ASAP7_75t_L g764 ( 
.A(n_554),
.B(n_511),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_654),
.B(n_190),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_640),
.B(n_332),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_SL g767 ( 
.A(n_614),
.B(n_332),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_629),
.B(n_194),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_574),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_580),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_551),
.B(n_337),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_568),
.B(n_482),
.Y(n_772)
);

INVxp33_ASAP7_75t_L g773 ( 
.A(n_668),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_654),
.B(n_194),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_580),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_555),
.B(n_195),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_632),
.B(n_195),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_533),
.B(n_196),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_635),
.B(n_196),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_537),
.B(n_294),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_663),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_635),
.B(n_199),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_590),
.B(n_199),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_663),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_612),
.B(n_204),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_547),
.B(n_296),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_526),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_539),
.A2(n_297),
.B1(n_246),
.B2(n_243),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_646),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_551),
.B(n_352),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_204),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_605),
.B(n_298),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_530),
.B(n_345),
.C(n_348),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_647),
.B(n_206),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_626),
.B(n_206),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_557),
.B(n_207),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_586),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_586),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_557),
.B(n_207),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_593),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_656),
.B(n_305),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_611),
.B(n_350),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_557),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_641),
.B(n_310),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_526),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_543),
.B(n_208),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_604),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_593),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_543),
.B(n_208),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_543),
.B(n_347),
.Y(n_810)
);

INVx8_ASAP7_75t_L g811 ( 
.A(n_604),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_557),
.B(n_347),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_587),
.B(n_351),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_604),
.B(n_351),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_658),
.A2(n_297),
.B1(n_354),
.B2(n_216),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_607),
.B(n_317),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_582),
.B(n_589),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_676),
.B(n_434),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_676),
.B(n_434),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_604),
.B(n_354),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_571),
.B(n_312),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_554),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_SL g823 ( 
.A1(n_571),
.A2(n_320),
.B1(n_319),
.B2(n_318),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_604),
.B(n_613),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_545),
.B(n_321),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_531),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_545),
.B(n_323),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_596),
.Y(n_828)
);

BUFx8_ASAP7_75t_L g829 ( 
.A(n_604),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_613),
.B(n_482),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_531),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_536),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_558),
.B(n_324),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_613),
.B(n_558),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_613),
.B(n_482),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_596),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_621),
.B(n_325),
.C(n_331),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_613),
.B(n_483),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_613),
.B(n_483),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_613),
.B(n_483),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_536),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_545),
.B(n_326),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_544),
.B(n_484),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_587),
.B(n_329),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_674),
.A2(n_335),
.B1(n_499),
.B2(n_494),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_544),
.B(n_484),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_627),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_696),
.B(n_556),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_679),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_702),
.B(n_587),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_741),
.A2(n_562),
.B(n_623),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_699),
.B(n_627),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_695),
.A2(n_581),
.B(n_584),
.C(n_585),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_713),
.A2(n_722),
.B1(n_817),
.B2(n_801),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_681),
.B(n_628),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_759),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_693),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_713),
.B(n_636),
.C(n_628),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_682),
.B(n_636),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_741),
.A2(n_625),
.B(n_623),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_744),
.A2(n_617),
.B(n_581),
.C(n_584),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_756),
.A2(n_625),
.B(n_546),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_685),
.B(n_639),
.Y(n_863)
);

AO21x1_ASAP7_75t_L g864 ( 
.A1(n_690),
.A2(n_644),
.B(n_639),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_724),
.B(n_587),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_684),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_740),
.B(n_545),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_753),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_722),
.A2(n_644),
.B(n_645),
.C(n_651),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_746),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_822),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_687),
.B(n_645),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_689),
.B(n_651),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_692),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_756),
.A2(n_546),
.B(n_538),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_724),
.A2(n_546),
.B(n_538),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_SL g877 ( 
.A1(n_768),
.A2(n_653),
.B(n_652),
.C(n_662),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_697),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_678),
.B(n_734),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_729),
.A2(n_538),
.B(n_550),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_729),
.A2(n_602),
.B(n_552),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_698),
.A2(n_602),
.B(n_552),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_694),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_720),
.A2(n_575),
.B(n_576),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_720),
.A2(n_550),
.B(n_618),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_762),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_738),
.A2(n_550),
.B(n_618),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_693),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_822),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_738),
.A2(n_595),
.B(n_618),
.Y(n_891)
);

AND2x6_ASAP7_75t_L g892 ( 
.A(n_824),
.B(n_575),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_700),
.B(n_652),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_707),
.A2(n_617),
.B(n_610),
.C(n_576),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_807),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_747),
.B(n_650),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_768),
.A2(n_595),
.B(n_583),
.Y(n_897)
);

AO21x1_ASAP7_75t_L g898 ( 
.A1(n_715),
.A2(n_665),
.B(n_653),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_766),
.B(n_670),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_801),
.B(n_662),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_803),
.B(n_587),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_832),
.A2(n_595),
.B(n_583),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_819),
.B(n_665),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_832),
.A2(n_583),
.B(n_615),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_716),
.B(n_528),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_755),
.B(n_528),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_761),
.B(n_528),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_701),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_807),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_829),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_712),
.A2(n_600),
.B1(n_588),
.B2(n_610),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_803),
.B(n_616),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_817),
.B(n_567),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_841),
.A2(n_567),
.B(n_615),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_841),
.A2(n_846),
.B(n_843),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_773),
.B(n_577),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_787),
.A2(n_567),
.B(n_615),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_816),
.B(n_528),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_703),
.B(n_577),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_L g920 ( 
.A1(n_780),
.A2(n_786),
.B(n_783),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_787),
.A2(n_567),
.B(n_615),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_816),
.B(n_528),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_805),
.A2(n_578),
.B(n_579),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_L g924 ( 
.A1(n_780),
.A2(n_578),
.B(n_579),
.Y(n_924)
);

AO21x2_ASAP7_75t_L g925 ( 
.A1(n_715),
.A2(n_809),
.B(n_806),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_805),
.A2(n_585),
.B(n_588),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_714),
.B(n_554),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_826),
.A2(n_600),
.B(n_616),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_719),
.B(n_528),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_804),
.A2(n_711),
.B1(n_709),
.B2(n_786),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_750),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_721),
.B(n_528),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_826),
.A2(n_616),
.B(n_666),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_804),
.A2(n_649),
.B1(n_673),
.B2(n_659),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_803),
.B(n_616),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_829),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_723),
.B(n_725),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_834),
.A2(n_675),
.B(n_666),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_731),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_802),
.A2(n_659),
.B(n_673),
.C(n_649),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_789),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_818),
.Y(n_942)
);

BUFx2_ASAP7_75t_SL g943 ( 
.A(n_772),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_732),
.B(n_659),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_680),
.B(n_683),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_739),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_831),
.A2(n_616),
.B(n_667),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_831),
.A2(n_675),
.B(n_671),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_782),
.A2(n_671),
.B(n_669),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_686),
.B(n_673),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_743),
.A2(n_669),
.B(n_667),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_750),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_701),
.B(n_541),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_748),
.A2(n_655),
.B(n_634),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_754),
.B(n_634),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_758),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_760),
.A2(n_655),
.B(n_634),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_704),
.B(n_727),
.Y(n_958)
);

BUFx4f_ASAP7_75t_L g959 ( 
.A(n_771),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_750),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_769),
.Y(n_961)
);

OAI321xp33_ASAP7_75t_L g962 ( 
.A1(n_793),
.A2(n_484),
.A3(n_499),
.B1(n_494),
.B2(n_471),
.C(n_507),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_770),
.A2(n_655),
.B(n_634),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_775),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_735),
.B(n_499),
.C(n_494),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_803),
.B(n_750),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_733),
.B(n_634),
.Y(n_967)
);

AOI33xp33_ASAP7_75t_L g968 ( 
.A1(n_821),
.A2(n_847),
.A3(n_800),
.B1(n_797),
.B2(n_836),
.B3(n_828),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_798),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_742),
.A2(n_655),
.B1(n_290),
.B2(n_286),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_808),
.B(n_655),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_736),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_718),
.A2(n_643),
.B(n_631),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_777),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_693),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_777),
.A2(n_281),
.B(n_227),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_688),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_815),
.A2(n_236),
.B(n_232),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_779),
.A2(n_300),
.B(n_228),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_779),
.A2(n_307),
.B(n_240),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_785),
.B(n_631),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_830),
.A2(n_643),
.B(n_631),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_767),
.B(n_471),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_791),
.B(n_13),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_833),
.A2(n_316),
.B(n_242),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_825),
.A2(n_219),
.B(n_247),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_794),
.B(n_631),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_717),
.B(n_631),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_810),
.A2(n_334),
.B(n_471),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_825),
.A2(n_333),
.B(n_262),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_827),
.B(n_631),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_827),
.A2(n_255),
.B(n_263),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_795),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_726),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_842),
.A2(n_264),
.B(n_267),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_842),
.A2(n_275),
.B(n_279),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_796),
.A2(n_609),
.B(n_553),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_763),
.B(n_643),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_796),
.A2(n_609),
.B(n_553),
.Y(n_999)
);

BUFx2_ASAP7_75t_SL g1000 ( 
.A(n_726),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_733),
.A2(n_507),
.B1(n_471),
.B2(n_609),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_776),
.B(n_792),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_788),
.A2(n_507),
.B1(n_471),
.B2(n_609),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_771),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_812),
.A2(n_609),
.B(n_553),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_812),
.A2(n_609),
.B(n_553),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_765),
.B(n_643),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_813),
.A2(n_553),
.B(n_541),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_792),
.A2(n_471),
.B(n_507),
.C(n_343),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_774),
.B(n_643),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_691),
.A2(n_471),
.B1(n_507),
.B2(n_541),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_795),
.A2(n_15),
.B(n_18),
.C(n_19),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_745),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_752),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_737),
.A2(n_751),
.B(n_749),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_752),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_790),
.B(n_643),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_813),
.A2(n_778),
.B(n_784),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_L g1019 ( 
.A(n_790),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_757),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_811),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_691),
.B(n_643),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_730),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_757),
.A2(n_553),
.B(n_541),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_SL g1025 ( 
.A(n_823),
.B(n_541),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_781),
.B(n_507),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_781),
.B(n_20),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_726),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_837),
.B(n_21),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_705),
.B(n_22),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_784),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_726),
.A2(n_511),
.B(n_541),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_726),
.A2(n_511),
.B(n_334),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_835),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_1004),
.B(n_764),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_920),
.A2(n_710),
.B(n_820),
.C(n_814),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_854),
.B(n_845),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_942),
.B(n_811),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_874),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_941),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1002),
.B(n_840),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_900),
.A2(n_844),
.B(n_799),
.C(n_706),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_878),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_903),
.B(n_811),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_890),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_852),
.A2(n_839),
.B1(n_838),
.B2(n_343),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_848),
.B(n_22),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_855),
.B(n_24),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_880),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_890),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_893),
.A2(n_299),
.B(n_330),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_899),
.B(n_26),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_856),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_946),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_956),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_961),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_964),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_975),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_873),
.A2(n_299),
.B1(n_330),
.B2(n_343),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_865),
.A2(n_299),
.B(n_330),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_969),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_866),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_977),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_866),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_865),
.A2(n_330),
.B(n_343),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_913),
.A2(n_330),
.B1(n_343),
.B2(n_37),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_972),
.Y(n_1067)
);

INVx6_ASAP7_75t_L g1068 ( 
.A(n_994),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_930),
.B(n_334),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_877),
.A2(n_334),
.B(n_31),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_945),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_975),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1016),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_945),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_959),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_937),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_869),
.A2(n_28),
.B(n_41),
.C(n_44),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_870),
.B(n_511),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_959),
.B(n_334),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_939),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_984),
.A2(n_28),
.B(n_49),
.C(n_50),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_877),
.A2(n_334),
.B(n_53),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_883),
.A2(n_334),
.B(n_511),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_859),
.A2(n_334),
.B(n_54),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1019),
.B(n_52),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_863),
.B(n_52),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_R g1087 ( 
.A(n_868),
.B(n_55),
.Y(n_1087)
);

AO21x2_ASAP7_75t_L g1088 ( 
.A1(n_864),
.A2(n_511),
.B(n_96),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_872),
.A2(n_55),
.B(n_57),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_968),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_968),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1020),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1002),
.B(n_57),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_913),
.B(n_887),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_869),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1031),
.Y(n_1096)
);

AOI22x1_ASAP7_75t_L g1097 ( 
.A1(n_875),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1013),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_SL g1099 ( 
.A1(n_984),
.A2(n_62),
.B(n_65),
.C(n_68),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_879),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_858),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_896),
.A2(n_82),
.B1(n_86),
.B2(n_92),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_849),
.B(n_102),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_919),
.Y(n_1104)
);

OA22x2_ASAP7_75t_L g1105 ( 
.A1(n_1023),
.A2(n_115),
.B1(n_120),
.B2(n_132),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_SL g1106 ( 
.A(n_974),
.B(n_134),
.C(n_140),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1019),
.B(n_142),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_851),
.A2(n_147),
.B(n_151),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_857),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_858),
.A2(n_153),
.B(n_156),
.C(n_161),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_890),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_867),
.A2(n_165),
.B(n_924),
.C(n_940),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_898),
.A2(n_1018),
.B(n_861),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_870),
.B(n_895),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_993),
.A2(n_1012),
.B(n_1030),
.C(n_849),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_967),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_860),
.A2(n_881),
.B(n_876),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_890),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_916),
.B(n_884),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_955),
.A2(n_971),
.B1(n_927),
.B2(n_1028),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1014),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_884),
.A2(n_895),
.B1(n_909),
.B2(n_910),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1015),
.B(n_867),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_989),
.A2(n_1009),
.B(n_850),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_882),
.A2(n_927),
.B(n_885),
.C(n_965),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_944),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_958),
.B(n_871),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_909),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_918),
.A2(n_922),
.B(n_905),
.C(n_853),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_931),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_934),
.A2(n_950),
.B1(n_857),
.B2(n_1021),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_950),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_983),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_910),
.B(n_936),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1027),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_954),
.A2(n_963),
.B(n_957),
.C(n_991),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_894),
.A2(n_911),
.B(n_965),
.C(n_1029),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_936),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_978),
.B(n_871),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_931),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_862),
.A2(n_949),
.B(n_902),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_889),
.B(n_1021),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_986),
.B(n_996),
.C(n_995),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_889),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_L g1145 ( 
.A(n_908),
.B(n_931),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_R g1146 ( 
.A(n_994),
.B(n_1025),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1000),
.A2(n_850),
.B1(n_992),
.B2(n_990),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1034),
.A2(n_925),
.B1(n_967),
.B2(n_943),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_952),
.B(n_960),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_952),
.B(n_960),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_952),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_952),
.B(n_960),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_914),
.A2(n_917),
.B(n_921),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1026),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1009),
.A2(n_981),
.B(n_987),
.C(n_926),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_904),
.A2(n_928),
.B(n_935),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_906),
.A2(n_907),
.B(n_962),
.C(n_1010),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_901),
.A2(n_912),
.B(n_935),
.Y(n_1158)
);

OR2x6_ASAP7_75t_SL g1159 ( 
.A(n_1017),
.B(n_1003),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_938),
.A2(n_912),
.B(n_901),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_948),
.A2(n_886),
.B(n_888),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_973),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_970),
.A2(n_908),
.B1(n_932),
.B2(n_929),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_966),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_925),
.B(n_923),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_891),
.A2(n_915),
.B(n_897),
.Y(n_1166)
);

AND2x2_ASAP7_75t_SL g1167 ( 
.A(n_1022),
.B(n_988),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_933),
.A2(n_947),
.B(n_951),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_998),
.B(n_1007),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_892),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_966),
.A2(n_980),
.B1(n_976),
.B2(n_979),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_892),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1001),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_892),
.B(n_985),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_892),
.B(n_1011),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_953),
.B(n_1032),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_982),
.A2(n_1024),
.B(n_1005),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_953),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_892),
.A2(n_1033),
.B1(n_999),
.B2(n_1006),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_997),
.A2(n_527),
.B(n_699),
.C(n_696),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1008),
.B(n_594),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_920),
.A2(n_854),
.B(n_1002),
.C(n_984),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_874),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_975),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_900),
.A2(n_852),
.B(n_893),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_942),
.B(n_594),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_854),
.B(n_594),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_849),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1165),
.A2(n_1129),
.A3(n_1157),
.B(n_1112),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1109),
.B(n_1172),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1076),
.B(n_1080),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1156),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_1093),
.B(n_1052),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1182),
.A2(n_1185),
.B(n_1180),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1185),
.B(n_1123),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_SL g1196 ( 
.A1(n_1095),
.A2(n_1077),
.B1(n_1089),
.B2(n_1115),
.C(n_1066),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1109),
.B(n_1172),
.Y(n_1197)
);

INVxp67_ASAP7_75t_SL g1198 ( 
.A(n_1188),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1132),
.A2(n_1125),
.B(n_1094),
.C(n_1180),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1039),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1068),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1047),
.A2(n_1137),
.B(n_1069),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1117),
.A2(n_1141),
.B(n_1166),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1117),
.A2(n_1141),
.B(n_1166),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1115),
.A2(n_1041),
.B(n_1137),
.C(n_1181),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_SL g1206 ( 
.A1(n_1059),
.A2(n_1091),
.B(n_1090),
.C(n_1135),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1081),
.A2(n_1099),
.B(n_1085),
.C(n_1101),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_1075),
.B(n_1040),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1048),
.A2(n_1086),
.B(n_1071),
.C(n_1074),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1186),
.B(n_1100),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1043),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1173),
.Y(n_1212)
);

BUFx8_ASAP7_75t_SL g1213 ( 
.A(n_1053),
.Y(n_1213)
);

NAND3x1_ASAP7_75t_L g1214 ( 
.A(n_1134),
.B(n_1103),
.C(n_1119),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1062),
.B(n_1064),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1049),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1153),
.A2(n_1156),
.B(n_1168),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_1132),
.A2(n_1110),
.B(n_1107),
.C(n_1106),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_1106),
.A2(n_1174),
.B(n_1131),
.C(n_1044),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1089),
.A2(n_1084),
.B(n_1070),
.C(n_1082),
.Y(n_1220)
);

BUFx2_ASAP7_75t_R g1221 ( 
.A(n_1159),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1173),
.A2(n_1061),
.B1(n_1057),
.B2(n_1183),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1168),
.A2(n_1161),
.B(n_1136),
.Y(n_1223)
);

OAI22x1_ASAP7_75t_L g1224 ( 
.A1(n_1097),
.A2(n_1138),
.B1(n_1128),
.B2(n_1114),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1042),
.A2(n_1070),
.B(n_1082),
.C(n_1084),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1054),
.A2(n_1055),
.B1(n_1056),
.B2(n_1105),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1104),
.B(n_1114),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1158),
.A2(n_1036),
.B(n_1175),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1045),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_SL g1230 ( 
.A(n_1143),
.B(n_1127),
.C(n_1139),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1051),
.A2(n_1113),
.B(n_1065),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1063),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1121),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1144),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1161),
.A2(n_1136),
.B(n_1083),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1098),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1150),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1126),
.B(n_1038),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_R g1239 ( 
.A(n_1068),
.B(n_1058),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1060),
.A2(n_1065),
.B(n_1160),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1042),
.A2(n_1120),
.B(n_1147),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1155),
.A2(n_1060),
.B(n_1158),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1051),
.A2(n_1116),
.B(n_1148),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1155),
.A2(n_1179),
.B(n_1108),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1108),
.A2(n_1171),
.B(n_1124),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1068),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1133),
.B(n_1035),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1167),
.B(n_1154),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1045),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1145),
.A2(n_1176),
.B(n_1143),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1102),
.B(n_1163),
.C(n_1169),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1067),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1073),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1072),
.B(n_1096),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1164),
.A2(n_1162),
.B(n_1170),
.C(n_1116),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1092),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1046),
.A2(n_1149),
.B(n_1124),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1088),
.A2(n_1151),
.A3(n_1172),
.B(n_1105),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1150),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1079),
.A2(n_1184),
.B(n_1058),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1172),
.A2(n_1152),
.B(n_1109),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1045),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_L g1263 ( 
.A(n_1050),
.B(n_1118),
.C(n_1111),
.Y(n_1263)
);

OA22x2_ASAP7_75t_L g1264 ( 
.A1(n_1122),
.A2(n_1087),
.B1(n_1078),
.B2(n_1152),
.Y(n_1264)
);

NAND3x1_ASAP7_75t_L g1265 ( 
.A(n_1184),
.B(n_1146),
.C(n_1111),
.Y(n_1265)
);

BUFx4_ASAP7_75t_SL g1266 ( 
.A(n_1109),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1050),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1088),
.A2(n_1144),
.A3(n_1178),
.B(n_1130),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1130),
.A2(n_1140),
.A3(n_1111),
.B(n_1118),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1140),
.A2(n_1142),
.B(n_1118),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1140),
.A2(n_1050),
.B(n_1078),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1182),
.A2(n_527),
.B(n_699),
.C(n_1093),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1165),
.A2(n_989),
.A3(n_864),
.B(n_898),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1165),
.A2(n_989),
.A3(n_864),
.B(n_898),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1076),
.B(n_854),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1182),
.A2(n_527),
.B1(n_563),
.B2(n_1093),
.C(n_571),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1093),
.A2(n_594),
.B1(n_527),
.B2(n_640),
.Y(n_1278)
);

OAI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1093),
.A2(n_599),
.B1(n_854),
.B2(n_930),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1165),
.A2(n_989),
.A3(n_864),
.B(n_898),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1039),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1093),
.B(n_630),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1075),
.B(n_1114),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1150),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1076),
.B(n_854),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1075),
.B(n_1114),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1186),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1182),
.A2(n_920),
.B(n_1002),
.C(n_854),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1094),
.B(n_854),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1182),
.A2(n_527),
.B(n_699),
.C(n_1093),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1100),
.B(n_887),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1134),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1039),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1076),
.B(n_854),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1187),
.B(n_594),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1053),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1156),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1182),
.A2(n_1095),
.B1(n_1093),
.B2(n_1070),
.C(n_1082),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1156),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1076),
.B(n_854),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_854),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_854),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1053),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1076),
.B(n_854),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1076),
.B(n_854),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1053),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1076),
.B(n_854),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1156),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_854),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1076),
.B(n_854),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1144),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1186),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_854),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1100),
.B(n_887),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1039),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1093),
.A2(n_594),
.B1(n_527),
.B2(n_640),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1156),
.Y(n_1322)
);

NAND2x1_ASAP7_75t_L g1323 ( 
.A(n_1150),
.B(n_1152),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1165),
.A2(n_989),
.A3(n_864),
.B(n_898),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_854),
.Y(n_1325)
);

AOI221x1_ASAP7_75t_L g1326 ( 
.A1(n_1182),
.A2(n_1095),
.B1(n_1093),
.B2(n_1070),
.C(n_1082),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1188),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1093),
.A2(n_854),
.B1(n_1182),
.B2(n_873),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1182),
.B(n_1180),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1076),
.B(n_854),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1186),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1185),
.B(n_1182),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1182),
.A2(n_920),
.B(n_1002),
.C(n_854),
.Y(n_1333)
);

INVx8_ASAP7_75t_L g1334 ( 
.A(n_1150),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1094),
.B(n_854),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1039),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1076),
.B(n_854),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1100),
.B(n_887),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1076),
.B(n_854),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1182),
.A2(n_920),
.B(n_1002),
.C(n_854),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1156),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1275),
.B(n_1286),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1279),
.A2(n_1316),
.B1(n_1303),
.B2(n_1304),
.Y(n_1343)
);

BUFx8_ASAP7_75t_L g1344 ( 
.A(n_1298),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1303),
.A2(n_1304),
.B1(n_1325),
.B2(n_1311),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1236),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1200),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1193),
.A2(n_1282),
.B1(n_1311),
.B2(n_1325),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1277),
.A2(n_1316),
.B1(n_1282),
.B2(n_1328),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1201),
.Y(n_1350)
);

CKINVDCx11_ASAP7_75t_R g1351 ( 
.A(n_1308),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1239),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1305),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1278),
.A2(n_1321),
.B1(n_1272),
.B2(n_1291),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1211),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1215),
.B(n_1292),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1289),
.A2(n_1333),
.B1(n_1340),
.B2(n_1205),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1226),
.A2(n_1264),
.B1(n_1222),
.B2(n_1251),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1213),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1290),
.A2(n_1335),
.B1(n_1331),
.B2(n_1251),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1293),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1296),
.A2(n_1337),
.B1(n_1312),
.B2(n_1306),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1221),
.A2(n_1297),
.B1(n_1246),
.B2(n_1287),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1216),
.Y(n_1364)
);

INVx4_ASAP7_75t_SL g1365 ( 
.A(n_1258),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1229),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1232),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1334),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1302),
.A2(n_1330),
.B1(n_1309),
.B2(n_1339),
.Y(n_1369)
);

BUFx4f_ASAP7_75t_L g1370 ( 
.A(n_1284),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1281),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1300),
.A2(n_1326),
.B1(n_1307),
.B2(n_1332),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1294),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1222),
.A2(n_1212),
.B1(n_1194),
.B2(n_1332),
.Y(n_1374)
);

BUFx8_ASAP7_75t_SL g1375 ( 
.A(n_1287),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1334),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1319),
.B(n_1338),
.Y(n_1377)
);

INVx8_ASAP7_75t_L g1378 ( 
.A(n_1334),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1214),
.A2(n_1209),
.B1(n_1198),
.B2(n_1327),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1202),
.A2(n_1194),
.B1(n_1191),
.B2(n_1331),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1293),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1234),
.Y(n_1382)
);

BUFx8_ASAP7_75t_SL g1383 ( 
.A(n_1210),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1202),
.A2(n_1248),
.B1(n_1336),
.B2(n_1320),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1276),
.A2(n_1317),
.B1(n_1295),
.B2(n_1329),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1233),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1227),
.B(n_1288),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1314),
.B(n_1248),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1267),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1285),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1266),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1247),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1196),
.A2(n_1208),
.B1(n_1224),
.B2(n_1218),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1283),
.A2(n_1315),
.B1(n_1318),
.B2(n_1252),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1323),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1253),
.A2(n_1238),
.B1(n_1256),
.B2(n_1195),
.Y(n_1397)
);

BUFx10_ASAP7_75t_L g1398 ( 
.A(n_1249),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1195),
.A2(n_1230),
.B1(n_1228),
.B2(n_1241),
.Y(n_1399)
);

INVx6_ASAP7_75t_L g1400 ( 
.A(n_1237),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1228),
.A2(n_1254),
.B1(n_1243),
.B2(n_1196),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1190),
.A2(n_1197),
.B1(n_1259),
.B2(n_1313),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1255),
.A2(n_1219),
.B1(n_1263),
.B2(n_1199),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1243),
.A2(n_1262),
.B1(n_1231),
.B2(n_1257),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1257),
.A2(n_1244),
.B1(n_1263),
.B2(n_1271),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1250),
.A2(n_1260),
.B1(n_1245),
.B2(n_1197),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1313),
.B(n_1206),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1223),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1269),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1225),
.A2(n_1207),
.B1(n_1220),
.B2(n_1203),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1258),
.A2(n_1189),
.B1(n_1268),
.B2(n_1270),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1204),
.A2(n_1261),
.B1(n_1240),
.B2(n_1189),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1189),
.A2(n_1242),
.B1(n_1268),
.B2(n_1217),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1235),
.A2(n_1192),
.B1(n_1322),
.B2(n_1310),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1299),
.A2(n_1301),
.B1(n_1341),
.B2(n_1274),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1268),
.A2(n_1273),
.B1(n_1274),
.B2(n_1280),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1273),
.A2(n_1274),
.B1(n_1280),
.B2(n_1324),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1324),
.A2(n_1277),
.B1(n_1279),
.B2(n_1311),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1324),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1277),
.A2(n_1279),
.B1(n_1304),
.B2(n_1303),
.Y(n_1420)
);

BUFx4_ASAP7_75t_R g1421 ( 
.A(n_1213),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1328),
.A2(n_1304),
.B(n_1303),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1229),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1277),
.A2(n_1279),
.B1(n_1304),
.B2(n_1303),
.Y(n_1424)
);

INVx3_ASAP7_75t_SL g1425 ( 
.A(n_1305),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1278),
.A2(n_1321),
.B1(n_1277),
.B2(n_854),
.Y(n_1426)
);

BUFx10_ASAP7_75t_L g1427 ( 
.A(n_1305),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1278),
.A2(n_1321),
.B1(n_1277),
.B2(n_854),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1239),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1236),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1212),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1213),
.Y(n_1432)
);

OAI22x1_ASAP7_75t_L g1433 ( 
.A1(n_1278),
.A2(n_1321),
.B1(n_599),
.B2(n_1093),
.Y(n_1433)
);

CKINVDCx11_ASAP7_75t_R g1434 ( 
.A(n_1308),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1278),
.A2(n_1321),
.B1(n_1277),
.B2(n_854),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1277),
.A2(n_1193),
.B1(n_1279),
.B2(n_753),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_1308),
.Y(n_1437)
);

CKINVDCx9p33_ASAP7_75t_R g1438 ( 
.A(n_1297),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1212),
.Y(n_1439)
);

BUFx2_ASAP7_75t_SL g1440 ( 
.A(n_1208),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1239),
.Y(n_1441)
);

CKINVDCx14_ASAP7_75t_R g1442 ( 
.A(n_1308),
.Y(n_1442)
);

BUFx8_ASAP7_75t_L g1443 ( 
.A(n_1298),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1265),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1213),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1308),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1277),
.A2(n_1321),
.B1(n_1278),
.B2(n_1193),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1213),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1193),
.A2(n_1282),
.B1(n_1304),
.B2(n_1303),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1282),
.A2(n_1037),
.B1(n_1226),
.B2(n_1278),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1213),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1239),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1213),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1334),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1277),
.A2(n_1279),
.B1(n_1304),
.B2(n_1303),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1334),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1236),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1265),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1277),
.A2(n_1279),
.B1(n_1304),
.B2(n_1303),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1236),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1193),
.A2(n_1282),
.B1(n_1304),
.B2(n_1303),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1212),
.Y(n_1462)
);

BUFx10_ASAP7_75t_L g1463 ( 
.A(n_1305),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1305),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1334),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1431),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1462),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1462),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1447),
.A2(n_1436),
.B1(n_1459),
.B2(n_1455),
.C(n_1424),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1439),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1439),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1409),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1342),
.B(n_1362),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1362),
.B(n_1369),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1377),
.B(n_1347),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1355),
.B(n_1364),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1367),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1371),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1373),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1365),
.B(n_1422),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1356),
.B(n_1345),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1426),
.A2(n_1428),
.B1(n_1435),
.B2(n_1345),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1387),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1417),
.A2(n_1404),
.B(n_1399),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1411),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1374),
.B(n_1401),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1408),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1365),
.B(n_1396),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1416),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1408),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1346),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1430),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1386),
.A2(n_1357),
.B(n_1410),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1379),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1457),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1421),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1460),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1369),
.B(n_1380),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_L g1499 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1450),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1343),
.B(n_1389),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1374),
.B(n_1401),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1399),
.B(n_1418),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1412),
.A2(n_1414),
.B(n_1413),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1418),
.B(n_1420),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1419),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1420),
.B(n_1424),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1453),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1372),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1372),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1394),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1354),
.A2(n_1459),
.B(n_1455),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1349),
.A2(n_1449),
.B(n_1348),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_SL g1513 ( 
.A(n_1445),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1390),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1400),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1417),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1375),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1407),
.Y(n_1518)
);

BUFx4f_ASAP7_75t_L g1519 ( 
.A(n_1391),
.Y(n_1519)
);

AO21x1_ASAP7_75t_SL g1520 ( 
.A1(n_1403),
.A2(n_1395),
.B(n_1406),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1395),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1397),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1397),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1344),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1388),
.Y(n_1525)
);

AOI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1415),
.A2(n_1414),
.B(n_1438),
.Y(n_1526)
);

AO21x1_ASAP7_75t_SL g1527 ( 
.A1(n_1385),
.A2(n_1380),
.B(n_1405),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1351),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1400),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1400),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1384),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1393),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1344),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1385),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1383),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1461),
.B(n_1358),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1358),
.B(n_1360),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1415),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1444),
.B(n_1458),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1363),
.A2(n_1458),
.B1(n_1444),
.B2(n_1370),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1398),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1443),
.B(n_1353),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1402),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1443),
.B(n_1464),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1402),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1350),
.Y(n_1546)
);

NOR3xp33_ASAP7_75t_L g1547 ( 
.A(n_1423),
.B(n_1361),
.C(n_1352),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1438),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1382),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1423),
.B(n_1366),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1475),
.B(n_1381),
.Y(n_1551)
);

AOI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1518),
.A2(n_1526),
.B(n_1509),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1482),
.A2(n_1442),
.B(n_1392),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1482),
.A2(n_1382),
.B1(n_1370),
.B2(n_1425),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1469),
.A2(n_1440),
.B1(n_1429),
.B2(n_1452),
.C(n_1441),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_SL g1556 ( 
.A1(n_1511),
.A2(n_1446),
.B(n_1434),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_1448),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1470),
.B(n_1427),
.Y(n_1558)
);

AND3x1_ASAP7_75t_L g1559 ( 
.A(n_1547),
.B(n_1437),
.C(n_1451),
.Y(n_1559)
);

OAI21xp33_ASAP7_75t_L g1560 ( 
.A1(n_1486),
.A2(n_1359),
.B(n_1432),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1493),
.A2(n_1378),
.B(n_1376),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1536),
.A2(n_1368),
.B1(n_1376),
.B2(n_1454),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_SL g1564 ( 
.A(n_1517),
.B(n_1378),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1496),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1481),
.B(n_1368),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_R g1567 ( 
.A(n_1528),
.B(n_1378),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1512),
.A2(n_1454),
.B(n_1456),
.C(n_1465),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1503),
.A2(n_1454),
.B(n_1456),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1481),
.B(n_1454),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1471),
.B(n_1456),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1503),
.A2(n_1456),
.B(n_1508),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1536),
.A2(n_1499),
.B(n_1537),
.C(n_1506),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1507),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1506),
.A2(n_1509),
.B1(n_1508),
.B2(n_1501),
.C(n_1486),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1488),
.B(n_1539),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1488),
.B(n_1539),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1501),
.A2(n_1521),
.B(n_1487),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_L g1579 ( 
.A(n_1494),
.B(n_1535),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1513),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1477),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1480),
.B(n_1548),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1466),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1476),
.B(n_1548),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1521),
.A2(n_1487),
.B(n_1490),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1537),
.A2(n_1498),
.B(n_1504),
.C(n_1502),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1534),
.B(n_1467),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1480),
.B(n_1468),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1527),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1480),
.B(n_1472),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1538),
.A2(n_1526),
.B(n_1485),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1534),
.B(n_1473),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1517),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1544),
.B(n_1546),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1504),
.A2(n_1502),
.B(n_1474),
.C(n_1485),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1510),
.A2(n_1500),
.B(n_1480),
.C(n_1538),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1510),
.B(n_1489),
.C(n_1500),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1478),
.B(n_1479),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1490),
.A2(n_1519),
.B(n_1484),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1515),
.B(n_1524),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1489),
.A2(n_1522),
.B1(n_1523),
.B2(n_1516),
.C(n_1479),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1543),
.A2(n_1545),
.B(n_1522),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1523),
.A2(n_1543),
.B(n_1545),
.C(n_1540),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1519),
.A2(n_1514),
.B(n_1484),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1527),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1581),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1583),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1569),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1575),
.A2(n_1484),
.B1(n_1520),
.B2(n_1516),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1483),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1578),
.B(n_1483),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1591),
.B(n_1576),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1484),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1585),
.B(n_1495),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1585),
.B(n_1495),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

OAI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1596),
.A2(n_1573),
.B1(n_1586),
.B2(n_1575),
.C(n_1604),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1590),
.A2(n_1531),
.B1(n_1533),
.B2(n_1497),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1576),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1582),
.B(n_1520),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1599),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1492),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1589),
.B(n_1492),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1587),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1587),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1590),
.A2(n_1532),
.B1(n_1491),
.B2(n_1513),
.Y(n_1627)
);

INVx8_ASAP7_75t_L g1628 ( 
.A(n_1577),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1606),
.A2(n_1531),
.B1(n_1533),
.B2(n_1491),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1552),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1558),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1592),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1556),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1617),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1617),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1608),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1618),
.A2(n_1602),
.B1(n_1560),
.B2(n_1606),
.C(n_1593),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1625),
.B(n_1593),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1617),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1618),
.A2(n_1602),
.B1(n_1598),
.B2(n_1555),
.C(n_1553),
.Y(n_1640)
);

OAI33xp33_ASAP7_75t_L g1641 ( 
.A1(n_1611),
.A2(n_1562),
.A3(n_1558),
.B1(n_1557),
.B2(n_1554),
.B3(n_1571),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1620),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1588),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1608),
.B(n_1614),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1608),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1618),
.A2(n_1555),
.B1(n_1597),
.B2(n_1603),
.C(n_1600),
.Y(n_1646)
);

BUFx2_ASAP7_75t_SL g1647 ( 
.A(n_1633),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1620),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1562),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1628),
.B(n_1600),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1615),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1607),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1607),
.Y(n_1655)
);

INVxp67_ASAP7_75t_SL g1656 ( 
.A(n_1615),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1625),
.B(n_1592),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1630),
.A2(n_1605),
.B(n_1505),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1613),
.B(n_1601),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1610),
.A2(n_1579),
.B1(n_1554),
.B2(n_1563),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1610),
.B(n_1568),
.C(n_1561),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1611),
.B(n_1570),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1607),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1612),
.B(n_1566),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1610),
.B(n_1561),
.C(n_1564),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_SL g1667 ( 
.A(n_1619),
.B(n_1629),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1651),
.B(n_1621),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1642),
.B(n_1631),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1626),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1594),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1642),
.B(n_1631),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1648),
.B(n_1623),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1634),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1648),
.B(n_1623),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1652),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1612),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1656),
.B(n_1622),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_1623),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1667),
.B(n_1623),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1634),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1634),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1643),
.B(n_1644),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1644),
.B(n_1624),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1612),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1653),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1653),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1635),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1635),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1649),
.B(n_1654),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1655),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1655),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1664),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1664),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1657),
.B(n_1616),
.Y(n_1697)
);

NAND2xp67_ASAP7_75t_L g1698 ( 
.A(n_1639),
.B(n_1550),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1649),
.B(n_1624),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1658),
.B(n_1622),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1657),
.B(n_1616),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1639),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1688),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1681),
.B(n_1649),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1678),
.B(n_1665),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1688),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1679),
.B(n_1665),
.Y(n_1709)
);

OR2x6_ASAP7_75t_L g1710 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1637),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1689),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1689),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1671),
.B(n_1637),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1693),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1649),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1693),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1683),
.Y(n_1718)
);

NOR2xp67_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1682),
.B(n_1647),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1694),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1682),
.B(n_1647),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1682),
.B(n_1660),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1679),
.B(n_1640),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1679),
.B(n_1645),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1694),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1669),
.B(n_1672),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1683),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1683),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1699),
.B(n_1651),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1695),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1669),
.B(n_1640),
.Y(n_1732)
);

INVx5_ASAP7_75t_L g1733 ( 
.A(n_1668),
.Y(n_1733)
);

INVx3_ASAP7_75t_SL g1734 ( 
.A(n_1668),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1695),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1692),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1636),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1668),
.B(n_1646),
.Y(n_1739)
);

NOR2x1p5_ASAP7_75t_SL g1740 ( 
.A(n_1676),
.B(n_1639),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1697),
.B(n_1636),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1690),
.Y(n_1742)
);

OAI22xp33_ASAP7_75t_SL g1743 ( 
.A1(n_1698),
.A2(n_1632),
.B1(n_1651),
.B2(n_1609),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1565),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1703),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1708),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1672),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1732),
.B(n_1711),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1712),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1739),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1719),
.B(n_1699),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1714),
.B(n_1672),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1733),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1713),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1704),
.B(n_1687),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1704),
.B(n_1687),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1706),
.B(n_1687),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1715),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1734),
.B(n_1673),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1739),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1720),
.A2(n_1692),
.B1(n_1670),
.B2(n_1701),
.C(n_1697),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1706),
.B(n_1686),
.Y(n_1762)
);

XNOR2xp5_ASAP7_75t_L g1763 ( 
.A(n_1710),
.B(n_1559),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1717),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1734),
.B(n_1673),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1707),
.B(n_1686),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1737),
.B(n_1673),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1721),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1726),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1718),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1707),
.B(n_1686),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1731),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1733),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1735),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1725),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1710),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1720),
.B(n_1692),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1718),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1737),
.B(n_1677),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1709),
.B(n_1701),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1763),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1763),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1745),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1750),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1753),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1745),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1746),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1760),
.A2(n_1748),
.B1(n_1776),
.B2(n_1710),
.Y(n_1788)
);

XNOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1747),
.B(n_1710),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1752),
.A2(n_1646),
.B1(n_1632),
.B2(n_1662),
.Y(n_1790)
);

OAI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1761),
.A2(n_1743),
.B1(n_1701),
.B2(n_1662),
.C(n_1670),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1746),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1775),
.A2(n_1729),
.B(n_1728),
.Y(n_1793)
);

AOI21xp33_ASAP7_75t_L g1794 ( 
.A1(n_1775),
.A2(n_1729),
.B(n_1728),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1751),
.A2(n_1733),
.B1(n_1727),
.B2(n_1661),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1780),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1751),
.A2(n_1641),
.B1(n_1632),
.B2(n_1659),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1773),
.A2(n_1722),
.B(n_1736),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1753),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1749),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1773),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1749),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1754),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1767),
.B(n_1723),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.B(n_1723),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1754),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1796),
.B(n_1780),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1781),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1804),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1784),
.B(n_1755),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1789),
.A2(n_1753),
.B(n_1777),
.Y(n_1811)
);

INVxp67_ASAP7_75t_SL g1812 ( 
.A(n_1784),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1797),
.A2(n_1755),
.B1(n_1756),
.B2(n_1757),
.C(n_1778),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1782),
.B(n_1779),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1791),
.A2(n_1764),
.B1(n_1758),
.B2(n_1774),
.C(n_1772),
.Y(n_1815)
);

OAI21xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1804),
.A2(n_1765),
.B(n_1759),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1805),
.B(n_1756),
.Y(n_1817)
);

NOR2x1_ASAP7_75t_L g1818 ( 
.A(n_1783),
.B(n_1546),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1783),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1790),
.A2(n_1733),
.B1(n_1771),
.B2(n_1766),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1786),
.B(n_1758),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1805),
.B(n_1779),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1789),
.A2(n_1632),
.B1(n_1778),
.B2(n_1770),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1788),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_SL g1825 ( 
.A(n_1798),
.B(n_1757),
.C(n_1759),
.Y(n_1825)
);

NOR2xp67_ASAP7_75t_L g1826 ( 
.A(n_1801),
.B(n_1733),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1817),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1813),
.A2(n_1795),
.B1(n_1786),
.B2(n_1787),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1808),
.B(n_1812),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1814),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1808),
.B(n_1801),
.Y(n_1831)
);

OAI21xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1815),
.A2(n_1799),
.B(n_1785),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1825),
.A2(n_1765),
.B(n_1722),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1823),
.A2(n_1794),
.B1(n_1793),
.B2(n_1802),
.C(n_1787),
.Y(n_1834)
);

AOI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1810),
.A2(n_1806),
.B(n_1800),
.Y(n_1835)
);

AOI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1824),
.A2(n_1802),
.B(n_1792),
.Y(n_1836)
);

XOR2xp5_ASAP7_75t_L g1837 ( 
.A(n_1811),
.B(n_1580),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1807),
.B(n_1762),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1821),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1829),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1831),
.B(n_1809),
.Y(n_1841)
);

AOI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1834),
.A2(n_1820),
.B(n_1826),
.C(n_1816),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1830),
.B(n_1822),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1827),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1838),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1828),
.B(n_1818),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1839),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_L g1848 ( 
.A(n_1837),
.B(n_1819),
.Y(n_1848)
);

NOR3x1_ASAP7_75t_L g1849 ( 
.A(n_1833),
.B(n_1803),
.C(n_1792),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_L g1850 ( 
.A(n_1832),
.B(n_1803),
.C(n_1769),
.Y(n_1850)
);

AOI222xp33_ASAP7_75t_L g1851 ( 
.A1(n_1840),
.A2(n_1740),
.B1(n_1770),
.B2(n_1836),
.C1(n_1772),
.C2(n_1769),
.Y(n_1851)
);

NAND5xp2_ASAP7_75t_L g1852 ( 
.A(n_1842),
.B(n_1835),
.C(n_1550),
.D(n_1716),
.E(n_1705),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1846),
.A2(n_1774),
.B1(n_1764),
.B2(n_1768),
.C(n_1738),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1850),
.A2(n_1742),
.B1(n_1676),
.B2(n_1684),
.C(n_1691),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_R g1855 ( 
.A(n_1844),
.B(n_1574),
.Y(n_1855)
);

AOI222xp33_ASAP7_75t_L g1856 ( 
.A1(n_1847),
.A2(n_1632),
.B1(n_1742),
.B2(n_1630),
.C1(n_1676),
.C2(n_1684),
.Y(n_1856)
);

AOI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1852),
.A2(n_1841),
.B(n_1845),
.C(n_1843),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1851),
.A2(n_1848),
.B(n_1849),
.Y(n_1858)
);

AOI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1853),
.A2(n_1736),
.B1(n_1684),
.B2(n_1676),
.C(n_1691),
.Y(n_1859)
);

OA22x2_ASAP7_75t_L g1860 ( 
.A1(n_1855),
.A2(n_1542),
.B1(n_1730),
.B2(n_1705),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1854),
.A2(n_1744),
.B(n_1741),
.C(n_1738),
.Y(n_1861)
);

AOI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1856),
.A2(n_1741),
.B(n_1730),
.C(n_1595),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1860),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1858),
.B(n_1709),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1857),
.B(n_1716),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1861),
.B(n_1725),
.Y(n_1866)
);

AO22x2_ASAP7_75t_SL g1867 ( 
.A1(n_1862),
.A2(n_1567),
.B1(n_1551),
.B2(n_1685),
.Y(n_1867)
);

NOR2x1_ASAP7_75t_L g1868 ( 
.A(n_1864),
.B(n_1863),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1865),
.B(n_1859),
.C(n_1730),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1866),
.A2(n_1684),
.B(n_1691),
.C(n_1702),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1868),
.B(n_1867),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1871),
.Y(n_1872)
);

AOI311xp33_ASAP7_75t_L g1873 ( 
.A1(n_1872),
.A2(n_1869),
.A3(n_1870),
.B(n_1696),
.C(n_1700),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1872),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1874),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1873),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1875),
.B(n_1876),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1876),
.A2(n_1680),
.B(n_1675),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1877),
.Y(n_1879)
);

OAI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_1878),
.B(n_1633),
.Y(n_1880)
);

INVxp67_ASAP7_75t_L g1881 ( 
.A(n_1880),
.Y(n_1881)
);

OAI221xp5_ASAP7_75t_R g1882 ( 
.A1(n_1881),
.A2(n_1627),
.B1(n_1661),
.B2(n_1674),
.C(n_1675),
.Y(n_1882)
);

AOI211xp5_ASAP7_75t_L g1883 ( 
.A1(n_1882),
.A2(n_1541),
.B(n_1549),
.C(n_1633),
.Y(n_1883)
);


endmodule