module fake_jpeg_1745_n_217 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_217);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_57),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_66),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_60),
.Y(n_98)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_82),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_54),
.B1(n_59),
.B2(n_68),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_96),
.B1(n_77),
.B2(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_67),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_69),
.B1(n_77),
.B2(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_62),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_98),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_70),
.B(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_107),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_80),
.B1(n_59),
.B2(n_68),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_117),
.B1(n_55),
.B2(n_64),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_116),
.Y(n_127)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_84),
.B1(n_55),
.B2(n_60),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_88),
.B1(n_92),
.B2(n_97),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_126),
.B1(n_76),
.B2(n_3),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_22),
.B1(n_48),
.B2(n_46),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_90),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_100),
.C(n_76),
.Y(n_144)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_58),
.B1(n_71),
.B2(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_0),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_20),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_82),
.B(n_64),
.C(n_63),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_0),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_63),
.B1(n_73),
.B2(n_76),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_52),
.B1(n_23),
.B2(n_24),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_1),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_135),
.B1(n_120),
.B2(n_125),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_156),
.B1(n_159),
.B2(n_8),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_160),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_157),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_26),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_138),
.Y(n_173)
);

OAI22x1_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_50),
.B1(n_43),
.B2(n_42),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_32),
.B(n_31),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_165),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_128),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_30),
.C(n_28),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_181),
.B1(n_182),
.B2(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_5),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_163),
.B1(n_142),
.B2(n_155),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_37),
.B(n_36),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_186),
.B1(n_170),
.B2(n_172),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_159),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_10),
.C(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

AOI221xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_166),
.B1(n_167),
.B2(n_171),
.C(n_175),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_199),
.B(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_187),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_181),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_190),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_201),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_188),
.B(n_194),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_204),
.A2(n_15),
.B(n_16),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_202),
.B(n_211),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_214),
.B(n_203),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_17),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_18),
.Y(n_217)
);


endmodule