module fake_jpeg_31410_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_1),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_20),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_6),
.C(n_3),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_3),
.B(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_11),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_11),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_22),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_36),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.C(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_39),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_44),
.C(n_37),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_28),
.Y(n_53)
);


endmodule