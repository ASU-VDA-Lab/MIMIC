module fake_jpeg_3703_n_188 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_56),
.B1(n_45),
.B2(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_1),
.Y(n_68)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_1),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_63),
.B1(n_50),
.B2(n_51),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_69),
.B1(n_51),
.B2(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_91),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_57),
.C(n_56),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_2),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_52),
.B1(n_20),
.B2(n_21),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_71),
.B1(n_60),
.B2(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_112),
.Y(n_135)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_54),
.B1(n_49),
.B2(n_48),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_116),
.B1(n_96),
.B2(n_93),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_52),
.B(n_64),
.C(n_49),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_116),
.Y(n_136)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_128),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_6),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_6),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_7),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_137),
.B1(n_136),
.B2(n_134),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_8),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_24),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_14),
.C(n_15),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_44),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_12),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_102),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_153),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_112),
.B(n_13),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_151),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_135),
.A2(n_28),
.B1(n_42),
.B2(n_39),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_26),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_29),
.C(n_38),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_124),
.C(n_31),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_16),
.B(n_17),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_19),
.B(n_22),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_154),
.C(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_155),
.B1(n_147),
.B2(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_33),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_172),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_174),
.C(n_149),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_143),
.C(n_141),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_167),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_145),
.B(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_180),
.C(n_179),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_177),
.B1(n_169),
.B2(n_168),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_161),
.C(n_176),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_35),
.B(n_37),
.Y(n_188)
);


endmodule