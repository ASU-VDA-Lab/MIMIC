module fake_jpeg_29506_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_7),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_61),
.B1(n_50),
.B2(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_52),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_58),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_0),
.C(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_52),
.B1(n_54),
.B2(n_44),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_60),
.B1(n_49),
.B2(n_46),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_44),
.B(n_53),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_4),
.C(n_6),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_8),
.Y(n_100)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_93),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_97),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_9),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_25),
.B1(n_42),
.B2(n_40),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_75),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_29),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_9),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_77),
.B1(n_11),
.B2(n_10),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_77),
.B1(n_10),
.B2(n_15),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_14),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_129),
.C(n_36),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_43),
.B1(n_18),
.B2(n_19),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_17),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_131),
.B(n_118),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_23),
.B(n_24),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_116),
.C(n_118),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.C(n_138),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_117),
.B1(n_108),
.B2(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_108),
.B1(n_117),
.B2(n_110),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_122),
.C(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_132),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_143),
.B(n_137),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_137),
.B(n_140),
.Y(n_147)
);

OAI221xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_128),
.B1(n_38),
.B2(n_39),
.C(n_37),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_103),
.Y(n_149)
);


endmodule