module fake_netlist_5_1128_n_1226 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1226);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1226;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_1222;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_284;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_443;
wire n_864;
wire n_173;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_1203;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1048;
wire n_946;
wire n_417;
wire n_932;
wire n_1008;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_212;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_252;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_1032;
wire n_929;
wire n_941;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_587;
wire n_191;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_171;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_204;
wire n_394;
wire n_250;
wire n_341;
wire n_1049;
wire n_992;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_1108;
wire n_908;
wire n_449;
wire n_325;
wire n_1073;
wire n_1100;
wire n_1214;
wire n_862;
wire n_1016;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_918;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_1077;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_1221;
wire n_654;
wire n_370;
wire n_1172;
wire n_1095;
wire n_1096;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_1208;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_1149;
wire n_882;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_1225;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_1020;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_897;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_181;
wire n_962;
wire n_1219;
wire n_1204;
wire n_1215;
wire n_1216;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_1218;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_1223;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_584;
wire n_336;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_168;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_1069;
wire n_969;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_1197;
wire n_1211;
wire n_306;
wire n_1093;
wire n_722;
wire n_907;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_466;
wire n_239;
wire n_1164;
wire n_630;
wire n_420;
wire n_1202;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_170;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_1190;
wire n_1224;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_1014;
wire n_917;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_1212;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_1217;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1131;
wire n_1059;
wire n_1084;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_180;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1220;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1207;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_1213;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_23),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_129),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_40),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_54),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_73),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_132),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_59),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_30),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_10),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_146),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_38),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_31),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_39),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_98),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_29),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_76),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_4),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_4),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_93),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_48),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_103),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_130),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_21),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_144),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_153),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_75),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_121),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_55),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_21),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_10),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_22),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_128),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_41),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_16),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_82),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_124),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_100),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_110),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_42),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_117),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_89),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_66),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_60),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_162),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_37),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_137),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_27),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_112),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_140),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_114),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_145),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_34),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_38),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_150),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_19),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_57),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_127),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_28),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_43),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_115),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_116),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_32),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_9),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_155),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_105),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_131),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_33),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_55),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_176),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_209),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_176),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_183),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_193),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_224),
.B(n_0),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_183),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_193),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_193),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_193),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_250),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_170),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_190),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_201),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_205),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_214),
.B(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_174),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_184),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_214),
.B(n_1),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_186),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_184),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_189),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_263),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_195),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_182),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_182),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_263),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_229),
.B(n_1),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_226),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_244),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_208),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_275),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_282),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_168),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_171),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_172),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_240),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_215),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_229),
.B(n_2),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_240),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_240),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_173),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_196),
.B(n_2),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_177),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_187),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_185),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_219),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_227),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_198),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_199),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_258),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_228),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_196),
.B(n_5),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_232),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_202),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_203),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_264),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_204),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_197),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_207),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_211),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_267),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_233),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_188),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_286),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_234),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_236),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_237),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_242),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_264),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_246),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_247),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_175),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_289),
.A2(n_285),
.B1(n_269),
.B2(n_268),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_291),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_365),
.B(n_243),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_300),
.Y(n_389)
);

OR2x6_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_288),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_303),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_304),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_305),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_350),
.B(n_175),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_305),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_308),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_352),
.B(n_258),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_361),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_169),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_308),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_319),
.A2(n_266),
.B(n_262),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_309),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_309),
.Y(n_411)
);

BUFx8_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_312),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_312),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_313),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_313),
.Y(n_416)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_292),
.B(n_288),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_314),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_293),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_297),
.B(n_290),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_362),
.B(n_265),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_178),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_294),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_358),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_347),
.A2(n_241),
.B1(n_272),
.B2(n_259),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_366),
.B(n_270),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_367),
.B(n_178),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_338),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_317),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_317),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_302),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_302),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_377),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_378),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_375),
.B(n_274),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_390),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_409),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_370),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_373),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_376),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_380),
.B(n_307),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_388),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_318),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_221),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_372),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_382),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_380),
.B(n_373),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_418),
.B(n_307),
.Y(n_476)
);

BUFx4f_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_417),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_445),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_439),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_383),
.B(n_321),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_310),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_387),
.B(n_346),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_406),
.B(n_325),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_387),
.B(n_310),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_311),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_325),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_428),
.B(n_311),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_399),
.B(n_339),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_394),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_390),
.B(n_329),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_390),
.B(n_332),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_390),
.A2(n_315),
.B1(n_295),
.B2(n_344),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_399),
.B(n_340),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_348),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_405),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_396),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_332),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_383),
.B(n_323),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_390),
.B(n_322),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_412),
.B(n_343),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_388),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_404),
.B(n_169),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_434),
.B(n_343),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_400),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_412),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_453),
.B(n_439),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_459),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_475),
.B(n_412),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_455),
.B(n_441),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_458),
.B(n_454),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_L g530 ( 
.A(n_476),
.B(n_354),
.C(n_353),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_465),
.B(n_460),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_L g532 ( 
.A(n_451),
.B(n_267),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_465),
.B(n_445),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_467),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_465),
.B(n_445),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_451),
.B(n_447),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_480),
.B(n_436),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_465),
.B(n_445),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_504),
.A2(n_500),
.B1(n_519),
.B2(n_502),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_453),
.B(n_441),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_467),
.B(n_445),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_453),
.B(n_169),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_472),
.B(n_445),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_514),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_458),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_472),
.B(n_485),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_485),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_519),
.B(n_351),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_500),
.A2(n_371),
.B1(n_337),
.B2(n_417),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_513),
.A2(n_333),
.B1(n_334),
.B2(n_328),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_499),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_506),
.B(n_448),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_506),
.B(n_448),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_448),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_509),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_500),
.A2(n_417),
.B1(n_434),
.B2(n_216),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_454),
.B(n_353),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_502),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_496),
.C(n_489),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_510),
.B(n_448),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_512),
.B(n_516),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_512),
.B(n_448),
.Y(n_566)
);

BUFx5_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_516),
.B(n_448),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_520),
.B(n_409),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_453),
.B(n_169),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_477),
.B(n_169),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_409),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_473),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_500),
.A2(n_417),
.B1(n_369),
.B2(n_360),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_514),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_514),
.B(n_354),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_479),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_481),
.Y(n_581)
);

BUFx6f_ASAP7_75t_SL g582 ( 
.A(n_514),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_498),
.A2(n_417),
.B1(n_360),
.B2(n_369),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_452),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_477),
.B(n_230),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_466),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_484),
.Y(n_588)
);

O2A1O1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_482),
.A2(n_433),
.B(n_405),
.C(n_447),
.Y(n_589)
);

BUFx5_ASAP7_75t_L g590 ( 
.A(n_450),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_487),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_477),
.A2(n_432),
.B(n_430),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_484),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_484),
.Y(n_594)
);

O2A1O1Ixp5_ASAP7_75t_L g595 ( 
.A1(n_477),
.A2(n_404),
.B(n_446),
.C(n_415),
.Y(n_595)
);

AOI22x1_ASAP7_75t_L g596 ( 
.A1(n_452),
.A2(n_456),
.B1(n_468),
.B2(n_457),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_491),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_466),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_505),
.B(n_400),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_487),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_468),
.B(n_230),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_468),
.B(n_230),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_507),
.B(n_401),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_500),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_497),
.A2(n_265),
.B1(n_404),
.B2(n_296),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_456),
.B(n_401),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_468),
.B(n_230),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_471),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_518),
.A2(n_349),
.B1(n_404),
.B2(n_424),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_494),
.B(n_402),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_464),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_457),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_464),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_402),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_533),
.A2(n_461),
.B(n_487),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_527),
.A2(n_515),
.B(n_492),
.C(n_478),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_576),
.B(n_483),
.Y(n_621)
);

O2A1O1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_522),
.A2(n_446),
.B(n_493),
.C(n_486),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_602),
.B(n_463),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_527),
.B(n_469),
.Y(n_624)
);

O2A1O1Ixp5_ASAP7_75t_L g625 ( 
.A1(n_542),
.A2(n_493),
.B(n_501),
.C(n_486),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_576),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_542),
.A2(n_495),
.B(n_491),
.Y(n_627)
);

AO22x1_ASAP7_75t_L g628 ( 
.A1(n_548),
.A2(n_481),
.B1(n_261),
.B2(n_273),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_535),
.A2(n_461),
.B(n_487),
.Y(n_629)
);

O2A1O1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_522),
.A2(n_446),
.B(n_503),
.C(n_501),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_544),
.B(n_545),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_606),
.B(n_463),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_529),
.B(n_513),
.Y(n_633)
);

AO21x1_ASAP7_75t_L g634 ( 
.A1(n_570),
.A2(n_495),
.B(n_503),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_531),
.B(n_463),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_538),
.A2(n_461),
.B(n_487),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g637 ( 
.A(n_563),
.B(n_324),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_539),
.B(n_181),
.C(n_179),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_540),
.A2(n_518),
.B1(n_517),
.B2(n_470),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_526),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_570),
.A2(n_461),
.B(n_487),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_571),
.A2(n_586),
.B(n_578),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_562),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_576),
.B(n_461),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_571),
.A2(n_586),
.B(n_572),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_589),
.A2(n_424),
.B(n_517),
.C(n_474),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_613),
.B(n_470),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_587),
.B(n_600),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_544),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_560),
.B(n_276),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_569),
.A2(n_461),
.B(n_470),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_L g653 ( 
.A(n_530),
.B(n_330),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_540),
.A2(n_284),
.B1(n_181),
.B2(n_280),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_523),
.B(n_470),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_525),
.A2(n_284),
.B1(n_280),
.B2(n_283),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_577),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_524),
.B(n_474),
.Y(n_658)
);

INVxp33_ASAP7_75t_SL g659 ( 
.A(n_537),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_528),
.B(n_474),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_547),
.B(n_474),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_582),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_521),
.B(n_179),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_536),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_546),
.A2(n_495),
.B(n_403),
.C(n_414),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_549),
.B(n_490),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_551),
.B(n_490),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_595),
.A2(n_517),
.B(n_490),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_554),
.B(n_490),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_592),
.A2(n_517),
.B(n_432),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_607),
.A2(n_283),
.B1(n_191),
.B2(n_225),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_553),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_532),
.A2(n_432),
.B(n_430),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_526),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_534),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_550),
.Y(n_677)
);

OAI321xp33_ASAP7_75t_L g678 ( 
.A1(n_559),
.A2(n_584),
.A3(n_575),
.B1(n_548),
.B2(n_565),
.C(n_552),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_614),
.B(n_617),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_532),
.A2(n_435),
.B(n_430),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_607),
.A2(n_192),
.B1(n_194),
.B2(n_200),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_536),
.B(n_278),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_604),
.A2(n_518),
.B(n_407),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_604),
.A2(n_435),
.B(n_410),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_550),
.B(n_438),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_536),
.Y(n_687)
);

AO21x1_ASAP7_75t_L g688 ( 
.A1(n_605),
.A2(n_414),
.B(n_403),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_558),
.A2(n_438),
.B(n_426),
.C(n_422),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_561),
.B(n_438),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_612),
.B(n_206),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_591),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_605),
.A2(n_518),
.B(n_407),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_608),
.B(n_561),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_610),
.A2(n_435),
.B(n_410),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_615),
.B(n_438),
.Y(n_696)
);

AND2x4_ASAP7_75t_SL g697 ( 
.A(n_581),
.B(n_243),
.Y(n_697)
);

AOI21xp33_ASAP7_75t_L g698 ( 
.A1(n_608),
.A2(n_279),
.B(n_212),
.Y(n_698)
);

AOI21x1_ASAP7_75t_L g699 ( 
.A1(n_610),
.A2(n_415),
.B(n_410),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_582),
.B(n_210),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_591),
.B(n_230),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_579),
.B(n_580),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_612),
.B(n_213),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_585),
.B(n_217),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_608),
.A2(n_518),
.B1(n_218),
.B2(n_222),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_591),
.A2(n_603),
.B(n_543),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_573),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_573),
.A2(n_518),
.B(n_407),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_541),
.A2(n_426),
.B(n_422),
.C(n_395),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_599),
.A2(n_220),
.B1(n_260),
.B2(n_271),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_591),
.B(n_223),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_603),
.A2(n_416),
.B(n_395),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_555),
.B(n_335),
.C(n_331),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_603),
.A2(n_557),
.B(n_556),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_SL g715 ( 
.A1(n_624),
.A2(n_611),
.B(n_616),
.C(n_597),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_646),
.A2(n_566),
.B(n_564),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_664),
.B(n_601),
.Y(n_717)
);

AO21x1_ASAP7_75t_L g718 ( 
.A1(n_638),
.A2(n_568),
.B(n_618),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_643),
.A2(n_624),
.B1(n_687),
.B2(n_620),
.Y(n_719)
);

BUFx12f_ASAP7_75t_L g720 ( 
.A(n_662),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_635),
.A2(n_609),
.B(n_603),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_714),
.A2(n_596),
.B(n_583),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_657),
.B(n_581),
.Y(n_723)
);

CKINVDCx14_ASAP7_75t_R g724 ( 
.A(n_662),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_637),
.B(n_590),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_R g726 ( 
.A(n_679),
.B(n_611),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_651),
.B(n_590),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_675),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_676),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_638),
.A2(n_590),
.B1(n_567),
.B2(n_518),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_677),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_641),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_651),
.B(n_623),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_644),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_674),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_694),
.A2(n_590),
.B1(n_567),
.B2(n_594),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_640),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_640),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_632),
.A2(n_583),
.B(n_574),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_677),
.A2(n_597),
.B1(n_594),
.B2(n_593),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_648),
.A2(n_593),
.B1(n_574),
.B2(n_588),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_633),
.A2(n_567),
.B1(n_590),
.B2(n_235),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_686),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_640),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_682),
.B(n_590),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_678),
.A2(n_598),
.B(n_588),
.C(n_429),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_682),
.B(n_567),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_668),
.A2(n_598),
.B(n_567),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_707),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_655),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_640),
.A2(n_231),
.B1(n_238),
.B2(n_239),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_649),
.B(n_336),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_631),
.B(n_567),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_649),
.B(n_567),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_SL g755 ( 
.A1(n_647),
.A2(n_341),
.B(n_345),
.C(n_444),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_658),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_660),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_661),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_631),
.B(n_429),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_L g760 ( 
.A1(n_656),
.A2(n_255),
.B(n_248),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_650),
.A2(n_245),
.B1(n_253),
.B2(n_252),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_SL g762 ( 
.A(n_672),
.B(n_256),
.C(n_251),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_SL g763 ( 
.A(n_659),
.B(n_243),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_704),
.B(n_626),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_706),
.A2(n_627),
.B(n_670),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_704),
.A2(n_444),
.B(n_443),
.C(n_431),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_SL g767 ( 
.A(n_621),
.B(n_700),
.C(n_671),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_626),
.B(n_431),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_650),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_666),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_650),
.B(n_443),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_650),
.B(n_692),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_697),
.B(n_440),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_698),
.A2(n_249),
.B(n_440),
.C(n_442),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_653),
.B(n_440),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_705),
.A2(n_442),
.B(n_421),
.C(n_395),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_692),
.B(n_442),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_628),
.B(n_6),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_700),
.B(n_437),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_722),
.A2(n_739),
.B(n_765),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_734),
.B(n_663),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_729),
.Y(n_783)
);

AND3x1_ASAP7_75t_L g784 ( 
.A(n_723),
.B(n_713),
.C(n_702),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_749),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_733),
.B(n_702),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_732),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_754),
.B(n_667),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_778),
.B(n_713),
.C(n_654),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_SL g790 ( 
.A1(n_774),
.A2(n_711),
.B(n_691),
.C(n_703),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_736),
.A2(n_692),
.B1(n_639),
.B2(n_669),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_735),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_720),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_767),
.A2(n_622),
.B(n_630),
.C(n_665),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_743),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_718),
.A2(n_634),
.A3(n_688),
.B(n_689),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_727),
.A2(n_625),
.B(n_696),
.C(n_709),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_745),
.A2(n_625),
.B(n_652),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_737),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_750),
.B(n_685),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_752),
.B(n_681),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_722),
.A2(n_699),
.B(n_709),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_747),
.A2(n_636),
.B(n_619),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_772),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_765),
.A2(n_629),
.B(n_692),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_772),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_763),
.B(n_710),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_SL g809 ( 
.A(n_726),
.B(n_690),
.C(n_673),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_773),
.Y(n_810)
);

AO31x2_ASAP7_75t_L g811 ( 
.A1(n_719),
.A2(n_680),
.A3(n_712),
.B(n_695),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_748),
.A2(n_642),
.B(n_645),
.Y(n_812)
);

AO31x2_ASAP7_75t_L g813 ( 
.A1(n_776),
.A2(n_684),
.A3(n_416),
.B(n_421),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_764),
.A2(n_683),
.B(n_693),
.C(n_708),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_742),
.A2(n_701),
.B1(n_437),
.B2(n_421),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_759),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_760),
.A2(n_416),
.B(n_437),
.C(n_267),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_716),
.A2(n_701),
.B(n_407),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_748),
.A2(n_437),
.B(n_420),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_762),
.A2(n_437),
.B1(n_420),
.B2(n_413),
.Y(n_820)
);

OA21x2_ASAP7_75t_L g821 ( 
.A1(n_716),
.A2(n_267),
.B(n_407),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_721),
.A2(n_267),
.B(n_407),
.Y(n_822)
);

AO31x2_ASAP7_75t_L g823 ( 
.A1(n_721),
.A2(n_267),
.A3(n_8),
.B(n_9),
.Y(n_823)
);

AO21x2_ASAP7_75t_L g824 ( 
.A1(n_715),
.A2(n_267),
.B(n_437),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_739),
.A2(n_78),
.B(n_166),
.Y(n_825)
);

AO31x2_ASAP7_75t_L g826 ( 
.A1(n_766),
.A2(n_741),
.A3(n_740),
.B(n_725),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_724),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_756),
.B(n_420),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_746),
.A2(n_420),
.B(n_413),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_769),
.B(n_7),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_772),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_755),
.A2(n_420),
.B(n_413),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_746),
.A2(n_77),
.B(n_165),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_730),
.A2(n_420),
.B(n_413),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_816),
.B(n_757),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_789),
.A2(n_808),
.B1(n_801),
.B2(n_786),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_786),
.A2(n_782),
.B1(n_779),
.B2(n_810),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_830),
.A2(n_775),
.B1(n_761),
.B2(n_770),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_788),
.A2(n_758),
.B1(n_753),
.B2(n_771),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_809),
.A2(n_751),
.B1(n_731),
.B2(n_768),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_780),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_783),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_833),
.A2(n_827),
.B1(n_807),
.B2(n_805),
.Y(n_843)
);

CKINVDCx11_ASAP7_75t_R g844 ( 
.A(n_802),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_785),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_800),
.B(n_717),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_787),
.A2(n_777),
.B1(n_771),
.B2(n_744),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_792),
.A2(n_777),
.B1(n_744),
.B2(n_738),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_795),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_831),
.A2(n_744),
.B1(n_738),
.B2(n_737),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_SL g851 ( 
.A1(n_805),
.A2(n_807),
.B1(n_788),
.B2(n_784),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_823),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_800),
.A2(n_738),
.B1(n_413),
.B2(n_411),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_793),
.A2(n_790),
.B1(n_791),
.B2(n_820),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_802),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_781),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_794),
.A2(n_791),
.B1(n_814),
.B2(n_828),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_828),
.B(n_7),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_823),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_802),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_799),
.Y(n_861)
);

CKINVDCx11_ASAP7_75t_R g862 ( 
.A(n_815),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_815),
.A2(n_413),
.B1(n_411),
.B2(n_408),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_823),
.Y(n_864)
);

CKINVDCx11_ASAP7_75t_R g865 ( 
.A(n_799),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_SL g866 ( 
.A1(n_825),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_806),
.B(n_11),
.Y(n_867)
);

BUFx2_ASAP7_75t_SL g868 ( 
.A(n_812),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_818),
.A2(n_411),
.B1(n_408),
.B2(n_398),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_824),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_824),
.Y(n_871)
);

CKINVDCx6p67_ASAP7_75t_R g872 ( 
.A(n_817),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_796),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_797),
.A2(n_411),
.B1(n_408),
.B2(n_398),
.Y(n_874)
);

BUFx8_ASAP7_75t_L g875 ( 
.A(n_796),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_796),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_811),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_818),
.A2(n_411),
.B1(n_408),
.B2(n_398),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_813),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_804),
.A2(n_411),
.B1(n_408),
.B2(n_398),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_829),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_829),
.A2(n_398),
.B1(n_389),
.B2(n_408),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_834),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_811),
.B(n_58),
.Y(n_884)
);

NAND2x1p5_ASAP7_75t_L g885 ( 
.A(n_803),
.B(n_389),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_822),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_398),
.B1(n_389),
.B2(n_14),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_819),
.Y(n_888)
);

INVx6_ASAP7_75t_L g889 ( 
.A(n_811),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_834),
.A2(n_389),
.B1(n_13),
.B2(n_14),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_798),
.A2(n_389),
.B1(n_13),
.B2(n_15),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_879),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_852),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_856),
.B(n_813),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_859),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_873),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_868),
.B(n_832),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_876),
.B(n_821),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_856),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_877),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_857),
.A2(n_826),
.B(n_79),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_870),
.B(n_826),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_871),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_877),
.B(n_826),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_877),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_877),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_889),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_889),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_885),
.A2(n_74),
.B(n_163),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_889),
.B(n_12),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_889),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_864),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_864),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_884),
.B(n_15),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_875),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_875),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_885),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_875),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_886),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_841),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_883),
.B(n_16),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_841),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_842),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_842),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_884),
.Y(n_926)
);

AO21x1_ASAP7_75t_SL g927 ( 
.A1(n_854),
.A2(n_17),
.B(n_18),
.Y(n_927)
);

OA21x2_ASAP7_75t_L g928 ( 
.A1(n_888),
.A2(n_17),
.B(n_18),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_924),
.B(n_851),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_901),
.A2(n_881),
.B(n_836),
.C(n_890),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_921),
.A2(n_881),
.B1(n_837),
.B2(n_891),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_924),
.B(n_867),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_922),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_922),
.B(n_849),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_921),
.B(n_858),
.Y(n_935)
);

AOI221xp5_ASAP7_75t_L g936 ( 
.A1(n_901),
.A2(n_866),
.B1(n_839),
.B2(n_835),
.C(n_838),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_910),
.B(n_884),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_910),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_922),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_910),
.B(n_861),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_912),
.B(n_845),
.Y(n_941)
);

CKINVDCx6p67_ASAP7_75t_R g942 ( 
.A(n_921),
.Y(n_942)
);

CKINVDCx10_ASAP7_75t_R g943 ( 
.A(n_927),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_921),
.A2(n_846),
.B1(n_860),
.B2(n_887),
.Y(n_944)
);

OA21x2_ASAP7_75t_L g945 ( 
.A1(n_901),
.A2(n_880),
.B(n_874),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_910),
.B(n_845),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_922),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_912),
.A2(n_862),
.B1(n_872),
.B2(n_843),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_922),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_912),
.B(n_860),
.Y(n_950)
);

NAND2x1_ASAP7_75t_L g951 ( 
.A(n_913),
.B(n_903),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_915),
.A2(n_862),
.B(n_872),
.C(n_844),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_925),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_913),
.A2(n_840),
.B(n_847),
.C(n_848),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_916),
.B(n_855),
.Y(n_955)
);

OA21x2_ASAP7_75t_L g956 ( 
.A1(n_893),
.A2(n_863),
.B(n_869),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_914),
.B(n_850),
.Y(n_957)
);

CKINVDCx6p67_ASAP7_75t_R g958 ( 
.A(n_914),
.Y(n_958)
);

AO32x2_ASAP7_75t_L g959 ( 
.A1(n_899),
.A2(n_878),
.A3(n_882),
.B1(n_865),
.B2(n_844),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_925),
.B(n_919),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_925),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_915),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_925),
.B(n_855),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_925),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_913),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_919),
.B(n_853),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_914),
.A2(n_865),
.B1(n_389),
.B2(n_22),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_920),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_964),
.B(n_904),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_968),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_960),
.B(n_903),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_904),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_933),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_939),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_947),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_949),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_953),
.B(n_902),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_961),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_934),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_963),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_938),
.B(n_904),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_935),
.B(n_903),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_938),
.B(n_904),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_963),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_951),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_938),
.B(n_892),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_946),
.B(n_892),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_965),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_965),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_942),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_930),
.A2(n_928),
.B1(n_914),
.B2(n_918),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_937),
.B(n_892),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_955),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_993),
.Y(n_994)
);

NAND2x1_ASAP7_75t_L g995 ( 
.A(n_985),
.B(n_955),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_975),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_975),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_982),
.Y(n_998)
);

INVx5_ASAP7_75t_SL g999 ( 
.A(n_989),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_975),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_980),
.B(n_932),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_980),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_973),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_985),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_991),
.A2(n_931),
.B1(n_930),
.B2(n_967),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_973),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_993),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_974),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_974),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_980),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_993),
.B(n_965),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_984),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_993),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_984),
.B(n_902),
.Y(n_1014)
);

AND3x2_ASAP7_75t_L g1015 ( 
.A(n_1007),
.B(n_918),
.C(n_950),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_1001),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1003),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_994),
.B(n_1007),
.Y(n_1018)
);

OAI31xp33_ASAP7_75t_L g1019 ( 
.A1(n_1013),
.A2(n_991),
.A3(n_990),
.B(n_931),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1013),
.B(n_986),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1003),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_994),
.B(n_986),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_994),
.B(n_986),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1003),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_998),
.B(n_990),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1022),
.B(n_994),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1016),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1022),
.B(n_999),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1017),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1017),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_L g1032 ( 
.A(n_1018),
.B(n_995),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1027),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1032),
.B(n_1018),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1028),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1028),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_SL g1037 ( 
.A1(n_1034),
.A2(n_1005),
.B(n_1019),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1033),
.A2(n_1005),
.B1(n_948),
.B2(n_1025),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1034),
.B(n_1033),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_SL g1040 ( 
.A1(n_1036),
.A2(n_1026),
.B1(n_1029),
.B2(n_935),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1035),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1035),
.B(n_1026),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

AOI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_1036),
.A2(n_1018),
.B(n_1030),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_1029),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1036),
.B(n_1023),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1035),
.Y(n_1047)
);

OAI31xp33_ASAP7_75t_L g1048 ( 
.A1(n_1037),
.A2(n_1027),
.A3(n_952),
.B(n_957),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1040),
.A2(n_995),
.B1(n_1027),
.B2(n_1022),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1038),
.A2(n_952),
.B(n_1031),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_1045),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1045),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1044),
.A2(n_1043),
.B(n_1039),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1039),
.A2(n_936),
.B(n_944),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1043),
.B(n_1022),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_1042),
.B(n_1046),
.C(n_1041),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_1047),
.A2(n_936),
.B(n_957),
.C(n_962),
.Y(n_1057)
);

NOR2x1_ASAP7_75t_L g1058 ( 
.A(n_1042),
.B(n_1021),
.Y(n_1058)
);

AOI211x1_ASAP7_75t_L g1059 ( 
.A1(n_1044),
.A2(n_1023),
.B(n_1020),
.C(n_982),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1045),
.B(n_1020),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1045),
.B(n_1021),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1041),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1045),
.B(n_1015),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1052),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1054),
.A2(n_958),
.B1(n_1004),
.B2(n_955),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1051),
.B(n_1052),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1057),
.A2(n_1050),
.B(n_1048),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1056),
.B(n_1063),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1060),
.B(n_1024),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1062),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1055),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1060),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1053),
.B(n_1024),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1057),
.A2(n_929),
.B(n_1011),
.C(n_950),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1049),
.A2(n_1011),
.B(n_916),
.C(n_944),
.Y(n_1075)
);

AOI32xp33_ASAP7_75t_L g1076 ( 
.A1(n_1058),
.A2(n_1011),
.A3(n_943),
.B1(n_1000),
.B2(n_996),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1061),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1061),
.A2(n_954),
.B(n_1001),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1059),
.A2(n_927),
.B1(n_916),
.B2(n_928),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1054),
.A2(n_916),
.B1(n_1000),
.B2(n_996),
.Y(n_1080)
);

AOI222xp33_ASAP7_75t_L g1081 ( 
.A1(n_1054),
.A2(n_954),
.B1(n_1011),
.B2(n_940),
.C1(n_999),
.C2(n_997),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1052),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1072),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1067),
.A2(n_928),
.B(n_941),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1071),
.B(n_999),
.Y(n_1085)
);

NAND4xp25_ASAP7_75t_SL g1086 ( 
.A(n_1076),
.B(n_988),
.C(n_997),
.D(n_989),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1068),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_1066),
.B(n_989),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1082),
.B(n_1002),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1064),
.B(n_1006),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1070),
.A2(n_928),
.B(n_1006),
.Y(n_1091)
);

OAI211xp5_ASAP7_75t_SL g1092 ( 
.A1(n_1081),
.A2(n_988),
.B(n_984),
.C(n_1008),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1077),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1073),
.B(n_979),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1080),
.B(n_999),
.Y(n_1095)
);

AND3x1_ASAP7_75t_L g1096 ( 
.A(n_1074),
.B(n_1009),
.C(n_1008),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1073),
.B(n_1069),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1078),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1065),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_1086),
.B(n_1079),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_L g1101 ( 
.A(n_1098),
.B(n_1097),
.Y(n_1101)
);

OAI211xp5_ASAP7_75t_L g1102 ( 
.A1(n_1087),
.A2(n_1075),
.B(n_928),
.C(n_24),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1083),
.Y(n_1103)
);

NAND4xp25_ASAP7_75t_L g1104 ( 
.A(n_1097),
.B(n_916),
.C(n_966),
.D(n_983),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1093),
.B(n_1085),
.Y(n_1105)
);

AOI211xp5_ASAP7_75t_L g1106 ( 
.A1(n_1095),
.A2(n_19),
.B(n_20),
.C(n_25),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1090),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_SL g1108 ( 
.A1(n_1089),
.A2(n_1009),
.B(n_1012),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_1096),
.A2(n_1010),
.B1(n_979),
.B2(n_970),
.C(n_971),
.Y(n_1109)
);

CKINVDCx16_ASAP7_75t_R g1110 ( 
.A(n_1099),
.Y(n_1110)
);

AOI322xp5_ASAP7_75t_L g1111 ( 
.A1(n_1088),
.A2(n_983),
.A3(n_981),
.B1(n_992),
.B2(n_927),
.C1(n_972),
.C2(n_969),
.Y(n_1111)
);

AOI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1092),
.A2(n_20),
.B(n_25),
.C(n_26),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_1084),
.B(n_1094),
.C(n_1090),
.Y(n_1113)
);

OAI31xp33_ASAP7_75t_L g1114 ( 
.A1(n_1091),
.A2(n_927),
.A3(n_928),
.B(n_29),
.Y(n_1114)
);

OAI211xp5_ASAP7_75t_L g1115 ( 
.A1(n_1087),
.A2(n_928),
.B(n_28),
.C(n_30),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1087),
.A2(n_909),
.B(n_1014),
.C(n_970),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1087),
.A2(n_928),
.B(n_971),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1087),
.A2(n_976),
.B1(n_978),
.B2(n_926),
.C(n_34),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1085),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1097),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_1087),
.B(n_909),
.C(n_926),
.Y(n_1121)
);

AOI322xp5_ASAP7_75t_L g1122 ( 
.A1(n_1087),
.A2(n_981),
.A3(n_983),
.B1(n_992),
.B2(n_969),
.C1(n_972),
.C2(n_987),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1085),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1110),
.A2(n_1113),
.B(n_1105),
.Y(n_1124)
);

AO22x2_ASAP7_75t_L g1125 ( 
.A1(n_1120),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_1125)
);

AOI221xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1112),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_1126)
);

OAI31xp33_ASAP7_75t_L g1127 ( 
.A1(n_1102),
.A2(n_35),
.A3(n_40),
.B(n_41),
.Y(n_1127)
);

AOI211xp5_ASAP7_75t_L g1128 ( 
.A1(n_1123),
.A2(n_42),
.B(n_43),
.C(n_46),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1106),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1100),
.A2(n_999),
.B1(n_945),
.B2(n_926),
.Y(n_1130)
);

XNOR2x1_ASAP7_75t_L g1131 ( 
.A(n_1101),
.B(n_47),
.Y(n_1131)
);

NAND5xp2_ASAP7_75t_L g1132 ( 
.A(n_1107),
.B(n_981),
.C(n_50),
.D(n_51),
.E(n_52),
.Y(n_1132)
);

OAI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1119),
.A2(n_945),
.B1(n_1014),
.B2(n_976),
.C(n_897),
.Y(n_1133)
);

AOI211xp5_ASAP7_75t_L g1134 ( 
.A1(n_1115),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1103),
.B(n_49),
.C(n_52),
.Y(n_1135)
);

AOI211xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1118),
.A2(n_53),
.B(n_56),
.C(n_977),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1104),
.A2(n_1108),
.B1(n_1114),
.B2(n_1117),
.C(n_1121),
.Y(n_1137)
);

XNOR2xp5_ASAP7_75t_L g1138 ( 
.A(n_1109),
.B(n_53),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1114),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_1111),
.Y(n_1140)
);

OAI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1116),
.A2(n_56),
.B(n_909),
.C(n_978),
.Y(n_1141)
);

OAI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1122),
.A2(n_897),
.B1(n_920),
.B2(n_923),
.C(n_919),
.Y(n_1142)
);

OAI211xp5_ASAP7_75t_L g1143 ( 
.A1(n_1106),
.A2(n_909),
.B(n_992),
.C(n_920),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1110),
.A2(n_923),
.B(n_893),
.Y(n_1144)
);

NAND4xp25_ASAP7_75t_L g1145 ( 
.A(n_1123),
.B(n_987),
.C(n_972),
.D(n_969),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_SL g1146 ( 
.A(n_1106),
.B(n_987),
.C(n_923),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1102),
.A2(n_893),
.B1(n_908),
.B2(n_906),
.C(n_895),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_1131),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1132),
.B(n_61),
.Y(n_1149)
);

NAND4xp75_ASAP7_75t_L g1150 ( 
.A(n_1124),
.B(n_956),
.C(n_896),
.D(n_906),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1125),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1140),
.A2(n_908),
.B1(n_906),
.B2(n_900),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1125),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1139),
.Y(n_1154)
);

NAND4xp75_ASAP7_75t_L g1155 ( 
.A(n_1127),
.B(n_956),
.C(n_896),
.D(n_908),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1135),
.B(n_977),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1136),
.B(n_977),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1146),
.A2(n_900),
.B1(n_911),
.B2(n_907),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1126),
.A2(n_900),
.B1(n_911),
.B2(n_907),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1129),
.B(n_62),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_SL g1161 ( 
.A(n_1141),
.B(n_63),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1128),
.B(n_959),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1138),
.B(n_1143),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1134),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1144),
.B(n_65),
.Y(n_1165)
);

XOR2xp5_ASAP7_75t_L g1166 ( 
.A(n_1130),
.B(n_67),
.Y(n_1166)
);

XNOR2xp5_ASAP7_75t_L g1167 ( 
.A(n_1137),
.B(n_68),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1147),
.B(n_900),
.C(n_902),
.Y(n_1168)
);

NAND4xp25_ASAP7_75t_L g1169 ( 
.A(n_1145),
.B(n_902),
.C(n_900),
.D(n_907),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1142),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1151),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_L g1172 ( 
.A(n_1153),
.B(n_1133),
.Y(n_1172)
);

OR3x1_ASAP7_75t_L g1173 ( 
.A(n_1154),
.B(n_896),
.C(n_71),
.Y(n_1173)
);

NAND4xp25_ASAP7_75t_L g1174 ( 
.A(n_1152),
.B(n_900),
.C(n_907),
.D(n_905),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1148),
.A2(n_900),
.B1(n_911),
.B2(n_907),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1167),
.B(n_895),
.C(n_897),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1156),
.Y(n_1177)
);

OAI322xp33_ASAP7_75t_L g1178 ( 
.A1(n_1170),
.A2(n_917),
.A3(n_892),
.B1(n_899),
.B2(n_905),
.C1(n_911),
.C2(n_959),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1149),
.B(n_892),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1156),
.B(n_911),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1164),
.B(n_905),
.Y(n_1181)
);

AOI322xp5_ASAP7_75t_L g1182 ( 
.A1(n_1163),
.A2(n_959),
.A3(n_905),
.B1(n_917),
.B2(n_899),
.C1(n_894),
.C2(n_898),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_L g1183 ( 
.A(n_1160),
.B(n_70),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1165),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_1166),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1171),
.B(n_1157),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1185),
.A2(n_1162),
.B1(n_1161),
.B2(n_1155),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1177),
.A2(n_1158),
.B1(n_1159),
.B2(n_1150),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1184),
.B(n_1168),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_L g1190 ( 
.A(n_1183),
.B(n_1172),
.C(n_1179),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1173),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1181),
.Y(n_1192)
);

XNOR2xp5_ASAP7_75t_L g1193 ( 
.A(n_1176),
.B(n_1169),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1180),
.Y(n_1194)
);

NAND4xp75_ASAP7_75t_L g1195 ( 
.A(n_1175),
.B(n_72),
.C(n_80),
.D(n_81),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1178),
.A2(n_905),
.B1(n_897),
.B2(n_917),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1174),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1182),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_SL g1199 ( 
.A1(n_1173),
.A2(n_897),
.B1(n_959),
.B2(n_917),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1184),
.A2(n_897),
.B(n_894),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1186),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1190),
.A2(n_917),
.B1(n_897),
.B2(n_894),
.Y(n_1202)
);

AO22x2_ASAP7_75t_L g1203 ( 
.A1(n_1192),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_1203)
);

OAI22x1_ASAP7_75t_L g1204 ( 
.A1(n_1187),
.A2(n_899),
.B1(n_894),
.B2(n_91),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_1191),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1198),
.A2(n_897),
.B1(n_90),
.B2(n_92),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1195),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1188),
.A2(n_897),
.B1(n_894),
.B2(n_898),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1189),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1194),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1210),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1201),
.B(n_1197),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1205),
.Y(n_1213)
);

XNOR2xp5_ASAP7_75t_L g1214 ( 
.A(n_1206),
.B(n_1193),
.Y(n_1214)
);

XNOR2xp5_ASAP7_75t_L g1215 ( 
.A(n_1209),
.B(n_1199),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1208),
.A2(n_1196),
.B1(n_1200),
.B2(n_894),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1213),
.A2(n_1207),
.B1(n_1204),
.B2(n_1203),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1211),
.A2(n_1202),
.B1(n_1203),
.B2(n_894),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1214),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1212),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1217),
.A2(n_1215),
.B1(n_1216),
.B2(n_898),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1221),
.A2(n_1220),
.B1(n_1219),
.B2(n_1218),
.Y(n_1222)
);

OAI22x1_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_87),
.B1(n_95),
.B2(n_96),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1223),
.Y(n_1224)
);

OAI221xp5_ASAP7_75t_R g1225 ( 
.A1(n_1224),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.C(n_107),
.Y(n_1225)
);

AOI211xp5_ASAP7_75t_L g1226 ( 
.A1(n_1225),
.A2(n_108),
.B(n_109),
.C(n_111),
.Y(n_1226)
);


endmodule