module fake_jpeg_23456_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_39),
.B1(n_27),
.B2(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_51),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_33),
.C(n_24),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_26),
.B1(n_21),
.B2(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_21),
.B1(n_26),
.B2(n_17),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_31),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_38),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_34),
.B1(n_39),
.B2(n_38),
.Y(n_75)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_29),
.B1(n_16),
.B2(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_30),
.B1(n_39),
.B2(n_38),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_75),
.B1(n_85),
.B2(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_69),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

NAND2x1p5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_41),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_41),
.B(n_35),
.C(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_0),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_27),
.B1(n_25),
.B2(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_2),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_62),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_92),
.A2(n_114),
.B1(n_78),
.B2(n_80),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_49),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_99),
.C(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_103),
.B1(n_108),
.B2(n_84),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_102),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_13),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_115),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_60),
.B1(n_51),
.B2(n_61),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_10),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_35),
.B(n_41),
.C(n_10),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_41),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_83),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_42),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_45),
.B1(n_44),
.B2(n_42),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_2),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_119),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_R g118 ( 
.A(n_102),
.B(n_73),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_130),
.B(n_114),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_129),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_63),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_63),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_70),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_72),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_133),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_86),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_95),
.B1(n_108),
.B2(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_138),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_85),
.B1(n_78),
.B2(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_41),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_148),
.B(n_154),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_96),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_169),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_106),
.B(n_97),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_166),
.B1(n_137),
.B2(n_68),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_106),
.B(n_97),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_167),
.B1(n_109),
.B2(n_76),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_172),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_76),
.B1(n_68),
.B2(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_41),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_130),
.C(n_127),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_177),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_128),
.B1(n_130),
.B2(n_122),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_178),
.B1(n_154),
.B2(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_118),
.B(n_127),
.C(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_127),
.B(n_142),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_194),
.B(n_148),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_113),
.C(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_185),
.B1(n_189),
.B2(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_74),
.B(n_104),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_124),
.B1(n_74),
.B2(n_66),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_156),
.B1(n_144),
.B2(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_150),
.C(n_167),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_211),
.C(n_41),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_155),
.B1(n_160),
.B2(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_210),
.B1(n_214),
.B2(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_213),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_157),
.B1(n_168),
.B2(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_173),
.B(n_180),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_150),
.B1(n_158),
.B2(n_170),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_147),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_91),
.B1(n_66),
.B2(n_41),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_175),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_41),
.B(n_3),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_5),
.B(n_6),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_41),
.B1(n_3),
.B2(n_4),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_182),
.B1(n_192),
.B2(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_183),
.C(n_191),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_235),
.B(n_202),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_234),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_236),
.B(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_200),
.C(n_204),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_231),
.Y(n_241)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_244),
.C(n_248),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_209),
.C(n_217),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_211),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_222),
.Y(n_254)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_221),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_210),
.C(n_202),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_216),
.B(n_218),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_219),
.B(n_7),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_231),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_14),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_258),
.B(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_229),
.C(n_225),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_256),
.C(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_224),
.C(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_236),
.C(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_239),
.C(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_6),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_264),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_246),
.CI(n_243),
.CON(n_264),
.SN(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_250),
.A2(n_241),
.B1(n_246),
.B2(n_9),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_268),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_267),
.C(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_268),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_7),
.C(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_8),
.C(n_9),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_262),
.B(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_278),
.C(n_279),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_273),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_10),
.C(n_11),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_281),
.B(n_12),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_283),
.Y(n_284)
);


endmodule