module fake_jpeg_29788_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_62),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_53),
.Y(n_152)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_16),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_56),
.B(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_60),
.Y(n_136)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_72),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_16),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g167 ( 
.A(n_76),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_14),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_101),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_90),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_38),
.B(n_41),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_14),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_104),
.Y(n_141)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_56),
.A2(n_102),
.B1(n_100),
.B2(n_94),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_142),
.B1(n_36),
.B2(n_28),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_41),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_112),
.B(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_64),
.B(n_38),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_117),
.B(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_51),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_51),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_165),
.Y(n_172)
);

INVx2_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g227 ( 
.A(n_128),
.B(n_145),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_57),
.A2(n_36),
.B1(n_28),
.B2(n_24),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_25),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_151),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_84),
.A2(n_50),
.B(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_42),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_91),
.B(n_42),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_153),
.B(n_163),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_59),
.B(n_48),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_75),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_65),
.B(n_27),
.Y(n_165)
);

BUFx4f_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_166),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_108),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_170),
.B(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_48),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_173),
.B(n_175),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_130),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_176),
.A2(n_177),
.B1(n_214),
.B2(n_21),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_82),
.B1(n_78),
.B2(n_77),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_114),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_180),
.B(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_50),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_186),
.Y(n_249)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_26),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_187),
.Y(n_279)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_111),
.B(n_26),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_191),
.B(n_198),
.Y(n_259)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_194),
.B(n_196),
.Y(n_277)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_141),
.B(n_46),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_136),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_44),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_200),
.B(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_27),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_114),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_124),
.B(n_37),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_208),
.B(n_3),
.C(n_4),
.Y(n_280)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_150),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_136),
.B(n_157),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_215),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_135),
.A2(n_73),
.B1(n_36),
.B2(n_28),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_132),
.B(n_32),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_223),
.B1(n_225),
.B2(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_219),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_132),
.B(n_29),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_220),
.B(n_221),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_157),
.B(n_29),
.Y(n_221)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

BUFx4f_ASAP7_75t_SL g267 ( 
.A(n_222),
.Y(n_267)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_140),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_120),
.B(n_29),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_226),
.A2(n_167),
.B(n_37),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_147),
.A2(n_37),
.B1(n_30),
.B2(n_21),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_107),
.B1(n_149),
.B2(n_37),
.Y(n_257)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_176),
.A2(n_161),
.B1(n_140),
.B2(n_131),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_230),
.A2(n_232),
.B1(n_183),
.B2(n_222),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_131),
.B1(n_134),
.B2(n_164),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_150),
.B(n_139),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_236),
.A2(n_248),
.B(n_258),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_123),
.B1(n_164),
.B2(n_134),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_238),
.A2(n_183),
.B1(n_178),
.B2(n_211),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g244 ( 
.A1(n_195),
.A2(n_166),
.B1(n_126),
.B2(n_149),
.Y(n_244)
);

AO22x2_ASAP7_75t_L g320 ( 
.A1(n_244),
.A2(n_266),
.B1(n_4),
.B2(n_6),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_186),
.A2(n_29),
.B(n_152),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_253),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_265),
.B1(n_168),
.B2(n_225),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_200),
.A2(n_29),
.B(n_152),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_197),
.A2(n_107),
.B(n_21),
.C(n_2),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_210),
.B(n_216),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_214),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_184),
.B(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_270),
.Y(n_313)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_196),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_275),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_196),
.A2(n_13),
.B1(n_12),
.B2(n_5),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_208),
.B(n_6),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_212),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_288),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_249),
.B(n_172),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_284),
.B(n_299),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_287),
.A2(n_310),
.B(n_320),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_193),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_203),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_302),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_174),
.C(n_207),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_311),
.Y(n_334)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_247),
.B1(n_279),
.B2(n_239),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_251),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_295),
.B(n_296),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_179),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_297),
.A2(n_306),
.B1(n_328),
.B2(n_233),
.Y(n_345)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_234),
.B(n_169),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_202),
.B1(n_185),
.B2(n_217),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_261),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_301),
.B(n_308),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_194),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_188),
.B1(n_223),
.B2(n_189),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_317),
.B1(n_247),
.B2(n_279),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_230),
.A2(n_194),
.B1(n_208),
.B2(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_260),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_236),
.B(n_206),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_229),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_314),
.Y(n_335)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_190),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_209),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_315),
.B(n_319),
.Y(n_363)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_4),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_321),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_268),
.B(n_6),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_6),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_322),
.B(n_324),
.Y(n_368)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_246),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_280),
.B(n_7),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_10),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_266),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_329),
.A2(n_10),
.B(n_11),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_10),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_287),
.A2(n_233),
.B(n_255),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_336),
.A2(n_349),
.B(n_353),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_282),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_340),
.C(n_362),
.Y(n_396)
);

OAI22x1_ASAP7_75t_SL g339 ( 
.A1(n_311),
.A2(n_266),
.B1(n_262),
.B2(n_244),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_339),
.A2(n_346),
.B1(n_355),
.B2(n_361),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_250),
.C(n_241),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_341),
.B(n_301),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_345),
.A2(n_351),
.B1(n_293),
.B2(n_326),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_292),
.A2(n_282),
.B(n_250),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_306),
.A2(n_244),
.B1(n_239),
.B2(n_241),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_243),
.B(n_267),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_290),
.A2(n_286),
.B1(n_297),
.B2(n_328),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_289),
.B(n_244),
.CI(n_267),
.CON(n_360),
.SN(n_360)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_360),
.B(n_327),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_245),
.B1(n_254),
.B2(n_256),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_283),
.B(n_267),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_310),
.A2(n_313),
.B(n_318),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_329),
.B(n_320),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_314),
.A2(n_254),
.B1(n_240),
.B2(n_243),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_369),
.A2(n_303),
.B1(n_298),
.B2(n_285),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_371),
.B(n_358),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_288),
.B(n_256),
.C(n_313),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_337),
.C(n_366),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_321),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_375),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_284),
.Y(n_374)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_320),
.Y(n_375)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_378),
.A2(n_381),
.B(n_392),
.Y(n_428)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_380),
.B(n_382),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_342),
.A2(n_317),
.B(n_324),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_383),
.A2(n_387),
.B(n_391),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_384),
.Y(n_413)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_312),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_389),
.B(n_408),
.Y(n_437)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_316),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_349),
.A2(n_307),
.B(n_320),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_325),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_402),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_394),
.A2(n_397),
.B1(n_369),
.B2(n_351),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_395),
.A2(n_406),
.B1(n_358),
.B2(n_370),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_345),
.A2(n_285),
.B1(n_304),
.B2(n_323),
.Y(n_397)
);

INVx8_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_398),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_347),
.A2(n_339),
.B1(n_342),
.B2(n_346),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_399),
.A2(n_356),
.B1(n_368),
.B2(n_367),
.Y(n_414)
);

BUFx24_ASAP7_75t_SL g400 ( 
.A(n_338),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_400),
.B(n_380),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_353),
.A2(n_344),
.B(n_340),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_381),
.B(n_402),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_362),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_350),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_403),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_367),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_404),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_388),
.Y(n_438)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_407),
.Y(n_431)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_357),
.Y(n_408)
);

AO21x2_ASAP7_75t_L g409 ( 
.A1(n_385),
.A2(n_392),
.B(n_401),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_409),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_372),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_410),
.B(n_421),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_412),
.A2(n_423),
.B1(n_398),
.B2(n_407),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_414),
.A2(n_417),
.B1(n_377),
.B2(n_379),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_370),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_395),
.B(n_397),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_405),
.B(n_341),
.Y(n_421)
);

NOR4xp25_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_371),
.C(n_332),
.D(n_331),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_429),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_394),
.A2(n_352),
.B1(n_331),
.B2(n_332),
.Y(n_423)
);

OAI22x1_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_383),
.B1(n_385),
.B2(n_406),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_376),
.B1(n_398),
.B2(n_415),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_432),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_396),
.B(n_403),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_435),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_404),
.B(n_393),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g436 ( 
.A(n_373),
.B(n_375),
.CI(n_378),
.CON(n_436),
.SN(n_436)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_376),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_387),
.C(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_413),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_451),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_456),
.B1(n_458),
.B2(n_415),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_446),
.A2(n_459),
.B1(n_463),
.B2(n_419),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_428),
.Y(n_473)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_391),
.B(n_386),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_390),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_454),
.Y(n_475)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_457),
.Y(n_484)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_425),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_462),
.B1(n_464),
.B2(n_467),
.Y(n_479)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_427),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_409),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_438),
.C(n_421),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_428),
.C(n_437),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_430),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_432),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_478),
.C(n_481),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_477),
.Y(n_506)
);

INVx6_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_476),
.A2(n_446),
.B1(n_457),
.B2(n_445),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_409),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_409),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_487),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_439),
.C(n_414),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_486),
.C(n_488),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_485),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_439),
.C(n_419),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_444),
.A2(n_412),
.B1(n_416),
.B2(n_436),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_435),
.C(n_431),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_430),
.C(n_411),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_445),
.C(n_461),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_484),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_499),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_492),
.A2(n_504),
.B1(n_503),
.B2(n_502),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_471),
.A2(n_445),
.B(n_451),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_493),
.A2(n_505),
.B(n_470),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_496),
.B(n_507),
.Y(n_508)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_498),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_479),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_454),
.B1(n_456),
.B2(n_443),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_503),
.Y(n_517)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_502),
.Y(n_509)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_478),
.A2(n_459),
.B(n_476),
.C(n_481),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_504),
.A2(n_496),
.B(n_499),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_483),
.B(n_486),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_510),
.A2(n_521),
.B(n_508),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_497),
.B(n_477),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_515),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_491),
.B(n_504),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_473),
.B(n_488),
.Y(n_514)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_514),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_501),
.B(n_469),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_501),
.A2(n_475),
.B1(n_490),
.B2(n_505),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_519),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_494),
.B(n_498),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_497),
.B(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_520),
.B(n_521),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_491),
.C(n_494),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_495),
.C(n_507),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_513),
.B(n_495),
.Y(n_523)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_523),
.Y(n_537)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_524),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_526),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_527),
.B(n_529),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_509),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_531),
.B(n_533),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_510),
.C(n_512),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_514),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_538),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_518),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_539),
.B(n_529),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_541),
.B(n_542),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_527),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_537),
.B(n_530),
.Y(n_543)
);

NOR2x1_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_540),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_546),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_547),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_548),
.A2(n_536),
.B(n_545),
.Y(n_549)
);

OAI221xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_534),
.B1(n_544),
.B2(n_528),
.C(n_509),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_534),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_532),
.Y(n_552)
);


endmodule