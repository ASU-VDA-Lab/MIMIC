module fake_jpeg_21192_n_135 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_19),
.Y(n_45)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_41),
.B1(n_15),
.B2(n_17),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.C(n_31),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_26),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_33),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_14),
.B(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_1),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_35),
.B1(n_24),
.B2(n_29),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_35),
.B1(n_36),
.B2(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_64),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_9),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_31),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_75),
.CI(n_1),
.CON(n_83),
.SN(n_83)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

AOI21x1_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_2),
.B(n_3),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_28),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_52),
.B(n_45),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_89),
.B(n_2),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_43),
.C(n_48),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_7),
.C(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_91),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_69),
.B1(n_72),
.B2(n_60),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_5),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_71),
.A3(n_59),
.B1(n_62),
.B2(n_72),
.C1(n_65),
.C2(n_74),
.Y(n_95)
);

OA21x2_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_82),
.B(n_83),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_64),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_85),
.C(n_84),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_103),
.B1(n_78),
.B2(n_90),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_69),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_80),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_54),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_92),
.B1(n_112),
.B2(n_104),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_109),
.C(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_86),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_102),
.B(n_99),
.C(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_94),
.B1(n_96),
.B2(n_92),
.C(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_109),
.C(n_108),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_87),
.C(n_89),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_103),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_124),
.C(n_115),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_106),
.C(n_9),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_7),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_127),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_79),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_113),
.C(n_67),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_122),
.B(n_12),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_10),
.C(n_12),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_56),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_129),
.Y(n_135)
);


endmodule