module fake_jpeg_18258_n_209 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_17),
.B1(n_21),
.B2(n_16),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_17),
.B1(n_15),
.B2(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_32),
.B1(n_34),
.B2(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_36),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_66),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_32),
.B1(n_38),
.B2(n_37),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_43),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_58),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_60),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_14),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_14),
.B1(n_19),
.B2(n_18),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_38),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_74),
.B1(n_22),
.B2(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_87),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_35),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_62),
.B(n_57),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_22),
.C(n_19),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_69),
.C(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_97),
.B1(n_96),
.B2(n_95),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_110),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_74),
.B1(n_56),
.B2(n_70),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_77),
.B(n_83),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_106),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_66),
.B1(n_72),
.B2(n_58),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_109),
.B1(n_77),
.B2(n_94),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_72),
.B1(n_53),
.B2(n_63),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_114),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_68),
.B1(n_73),
.B2(n_61),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_81),
.B1(n_82),
.B2(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_61),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_77),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_116),
.B1(n_104),
.B2(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_57),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_117),
.B1(n_112),
.B2(n_108),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_132),
.B1(n_135),
.B2(n_139),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_84),
.C(n_94),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_115),
.C(n_106),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_92),
.B1(n_87),
.B2(n_89),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_79),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_81),
.B1(n_78),
.B2(n_5),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_98),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_98),
.B1(n_106),
.B2(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_151),
.B1(n_158),
.B2(n_130),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_138),
.C(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_121),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_156),
.B1(n_139),
.B2(n_78),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_125),
.C(n_140),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_129),
.C(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_127),
.C(n_132),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_171),
.B1(n_157),
.B2(n_155),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_122),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_145),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_172),
.B(n_178),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_142),
.B1(n_144),
.B2(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_158),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_6),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_8),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_166),
.B1(n_165),
.B2(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_184),
.B1(n_180),
.B2(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_162),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_6),
.B(n_7),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_9),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_8),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_179),
.C(n_173),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_188),
.B(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_187),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_13),
.B(n_10),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g202 ( 
.A(n_200),
.B(n_192),
.Y(n_202)
);

OAI21x1_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_194),
.B(n_10),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_205),
.B(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_9),
.C(n_11),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_207),
.A2(n_12),
.B(n_13),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_12),
.Y(n_209)
);


endmodule