module fake_jpeg_11348_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_23),
.B(n_10),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_1),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_48),
.B1(n_40),
.B2(n_43),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_7),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_36),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_24),
.C(n_34),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_76),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_73),
.B1(n_74),
.B2(n_58),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_57),
.B1(n_41),
.B2(n_64),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_8),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AO21x2_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_25),
.B(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_94),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_71),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_18),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_9),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_11),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_14),
.C(n_17),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_99),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_20),
.C(n_22),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_91),
.B1(n_95),
.B2(n_83),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_101),
.B(n_88),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_98),
.A3(n_89),
.B1(n_101),
.B2(n_92),
.C1(n_30),
.C2(n_31),
.Y(n_105)
);

OAI322xp33_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.A3(n_103),
.B1(n_102),
.B2(n_28),
.C1(n_29),
.C2(n_32),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_26),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_27),
.B(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_82),
.Y(n_111)
);


endmodule