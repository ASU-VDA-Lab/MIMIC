module fake_netlist_6_119_n_133 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_61, n_39, n_63, n_60, n_59, n_32, n_4, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_133);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_133;

wire n_91;
wire n_119;
wire n_88;
wire n_98;
wire n_113;
wire n_73;
wire n_68;
wire n_83;
wire n_101;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_75;
wire n_109;
wire n_122;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_112;
wire n_81;
wire n_76;
wire n_124;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_116;
wire n_117;
wire n_118;
wire n_65;
wire n_93;
wire n_80;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_115;
wire n_69;
wire n_128;
wire n_79;

INVx5_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AOI22x1_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_61),
.B1(n_48),
.B2(n_52),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_9),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_37),
.A2(n_13),
.B1(n_6),
.B2(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_11),
.Y(n_82)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_57),
.B(n_19),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_60),
.B(n_8),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_18),
.B(n_15),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_2),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_5),
.B(n_10),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_12),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_17),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_23),
.Y(n_98)
);

NOR2xp67_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_62),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_82),
.B1(n_86),
.B2(n_78),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_69),
.B(n_74),
.C(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_87),
.B(n_84),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_76),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_100),
.B(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_67),
.B1(n_83),
.B2(n_68),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_93),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_24),
.B(n_25),
.Y(n_109)
);

OAI21x1_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_26),
.B(n_28),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_32),
.B(n_36),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_106),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_105),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_118),
.B1(n_124),
.B2(n_122),
.Y(n_127)
);

NAND4xp75_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_125),
.C(n_109),
.D(n_117),
.Y(n_128)
);

NAND2x1p5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_114),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_123),
.B1(n_111),
.B2(n_42),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_59),
.B1(n_40),
.B2(n_44),
.Y(n_131)
);

AOI221x1_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_38),
.B1(n_45),
.B2(n_47),
.C(n_49),
.Y(n_132)
);

OR2x6_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_51),
.Y(n_133)
);


endmodule