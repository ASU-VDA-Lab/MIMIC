module real_jpeg_21163_n_11 (n_5, n_4, n_8, n_0, n_256, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_256;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_0),
.A2(n_2),
.B1(n_17),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_0),
.A2(n_6),
.B1(n_23),
.B2(n_27),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_5),
.B1(n_27),
.B2(n_52),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_0),
.A2(n_4),
.B1(n_27),
.B2(n_46),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_1),
.A2(n_2),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_6),
.B1(n_16),
.B2(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_4),
.B1(n_16),
.B2(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_5),
.B1(n_16),
.B2(n_52),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_10),
.B1(n_17),
.B2(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_20),
.B(n_39),
.C(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_4),
.A2(n_7),
.B1(n_44),
.B2(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_4),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_4),
.A2(n_9),
.B1(n_46),
.B2(n_53),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_10),
.B1(n_39),
.B2(n_46),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_4),
.A2(n_39),
.B(n_53),
.C(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_9),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_5),
.B(n_85),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_10),
.B1(n_39),
.B2(n_52),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_5),
.A2(n_9),
.B(n_10),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_8),
.B1(n_20),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_6),
.A2(n_7),
.B1(n_23),
.B2(n_44),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_10),
.B1(n_23),
.B2(n_39),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_10),
.B(n_98),
.Y(n_97)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_10),
.B(n_23),
.C(n_143),
.Y(n_142)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_10),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_45),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_32),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_30),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_24),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_18),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_25),
.B(n_34),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_62),
.B(n_254),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_57),
.C(n_58),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_35),
.A2(n_36),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.C(n_48),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_37),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_37),
.A2(n_74),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_37),
.A2(n_76),
.B(n_94),
.C(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_37),
.A2(n_74),
.B1(n_194),
.B2(n_195),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_37),
.A2(n_74),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_37),
.A2(n_195),
.B(n_214),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_37),
.A2(n_74),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_37),
.A2(n_74),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_39),
.B(n_51),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_39),
.B(n_88),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_39),
.A2(n_44),
.B(n_46),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_40),
.A2(n_48),
.B1(n_224),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_40),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_48),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_48),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_56),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_51),
.A2(n_54),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OA22x2_ASAP7_75t_SL g210 ( 
.A1(n_51),
.A2(n_54),
.B1(n_56),
.B2(n_199),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_52),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_57),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_247),
.B(n_253),
.Y(n_62)
);

OAI321xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_219),
.A3(n_239),
.B1(n_245),
.B2(n_246),
.C(n_256),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_204),
.B(n_218),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_186),
.B(n_203),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_113),
.B(n_168),
.C(n_185),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_102),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_68),
.B(n_102),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_91),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_81),
.B2(n_82),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_70),
.B(n_82),
.C(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI211xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_74),
.B(n_75),
.C(n_80),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_79),
.B1(n_83),
.B2(n_90),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_79),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_79),
.B1(n_120),
.B2(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_99),
.C(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_72),
.A2(n_79),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_72),
.B(n_151),
.C(n_157),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_72),
.A2(n_79),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_72),
.B(n_83),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_72),
.B(n_175),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_74),
.B(n_77),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_74),
.B(n_224),
.C(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_74),
.B(n_233),
.C(n_238),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_75),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_76),
.A2(n_79),
.B(n_145),
.C(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_76),
.A2(n_77),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_76),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_76),
.B(n_210),
.Y(n_211)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_99),
.C(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_80),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_84),
.A2(n_88),
.B1(n_89),
.B2(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_101),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_92),
.A2(n_93),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_92),
.A2(n_93),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_109),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_109),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_99),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_154)
);

NAND2x1_ASAP7_75t_SL g158 ( 
.A(n_99),
.B(n_142),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_110),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_104),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_106),
.B1(n_141),
.B2(n_145),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_110),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_167),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_160),
.B(n_166),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_147),
.B(n_159),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_138),
.B(n_146),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_127),
.B(n_137),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_122),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_170),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_182),
.B2(n_184),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_181),
.C(n_184),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_178),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_183),
.B(n_202),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_191),
.B(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_188),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_205),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.CI(n_201),
.CON(n_189),
.SN(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_191),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_200),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_197),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_197),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_216),
.B2(n_217),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_213),
.C(n_217),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_211),
.A2(n_221),
.B1(n_228),
.B2(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_216),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_231),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_231),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.C(n_229),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_230),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_250),
.Y(n_252)
);


endmodule