module fake_jpeg_31672_n_445 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_48),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_54),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_77),
.Y(n_101)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_16),
.B(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_86),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_87),
.Y(n_124)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_92),
.Y(n_133)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_90),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_18),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_43),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_23),
.B1(n_44),
.B2(n_19),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_76),
.B1(n_43),
.B2(n_71),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_46),
.B1(n_41),
.B2(n_23),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_96),
.A2(n_98),
.B1(n_121),
.B2(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_97),
.B(n_128),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_41),
.B1(n_23),
.B2(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_44),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_20),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_32),
.B1(n_22),
.B2(n_39),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_104),
.A2(n_145),
.B1(n_20),
.B2(n_60),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_32),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_122),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_65),
.A2(n_18),
.B1(n_37),
.B2(n_24),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_29),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_135),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_29),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_27),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_143),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_73),
.A2(n_18),
.B1(n_37),
.B2(n_33),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_18),
.B1(n_37),
.B2(n_33),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_147),
.B1(n_76),
.B2(n_68),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_58),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_39),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_5),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_59),
.A2(n_40),
.B1(n_24),
.B2(n_43),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_86),
.A2(n_37),
.B1(n_40),
.B2(n_27),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_150),
.Y(n_213)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_152),
.A2(n_110),
.B(n_11),
.C(n_12),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_99),
.A2(n_62),
.B(n_37),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_154),
.A2(n_190),
.B(n_11),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_156),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_162),
.B1(n_156),
.B2(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_100),
.A2(n_83),
.B1(n_81),
.B2(n_78),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_192),
.B1(n_195),
.B2(n_110),
.Y(n_219)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_53),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_161),
.B(n_163),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_95),
.A2(n_43),
.B1(n_50),
.B2(n_93),
.Y(n_162)
);

OA22x2_ASAP7_75t_SL g218 ( 
.A1(n_162),
.A2(n_145),
.B1(n_136),
.B2(n_129),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_43),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_142),
.B1(n_105),
.B2(n_118),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_176),
.B1(n_188),
.B2(n_114),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_2),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_104),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_101),
.B(n_3),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_94),
.C(n_116),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_178),
.B(n_8),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_180),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_118),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_6),
.B(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_113),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_140),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_218),
.B1(n_155),
.B2(n_195),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_223),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_200),
.A2(n_206),
.B1(n_222),
.B2(n_146),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_205),
.B(n_184),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_134),
.B1(n_111),
.B2(n_123),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_233),
.C(n_175),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_219),
.A2(n_226),
.B1(n_126),
.B2(n_134),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_159),
.B1(n_163),
.B2(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_182),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_110),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_215),
.B(n_190),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_236),
.A2(n_265),
.B1(n_270),
.B2(n_211),
.Y(n_288)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_238),
.A2(n_260),
.B(n_151),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_239),
.A2(n_244),
.B1(n_246),
.B2(n_253),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_243),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_172),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_164),
.B1(n_113),
.B2(n_140),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_256),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_136),
.B1(n_129),
.B2(n_146),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_148),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_233),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_254),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_218),
.B1(n_235),
.B2(n_219),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_148),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_222),
.B1(n_221),
.B2(n_225),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_160),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_165),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_257),
.B(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_204),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_259),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_149),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_168),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_198),
.A2(n_126),
.B1(n_186),
.B2(n_112),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_268),
.B1(n_211),
.B2(n_177),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_198),
.A2(n_183),
.B1(n_167),
.B2(n_193),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_263),
.A2(n_230),
.B1(n_217),
.B2(n_227),
.Y(n_297)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_222),
.A2(n_208),
.B1(n_107),
.B2(n_120),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_203),
.B(n_170),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_230),
.B(n_185),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_222),
.A2(n_174),
.B1(n_150),
.B2(n_187),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_207),
.C(n_225),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_290),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_274),
.A2(n_286),
.B1(n_293),
.B2(n_300),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_203),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_239),
.A2(n_213),
.B1(n_212),
.B2(n_211),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_297),
.B1(n_266),
.B2(n_267),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_289),
.B1(n_298),
.B2(n_246),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_236),
.A2(n_265),
.B1(n_251),
.B2(n_256),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_217),
.C(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_253),
.A2(n_213),
.B1(n_177),
.B2(n_123),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_238),
.A2(n_220),
.B1(n_202),
.B2(n_228),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_244),
.A2(n_202),
.B1(n_228),
.B2(n_111),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_262),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_303),
.A2(n_307),
.B1(n_300),
.B2(n_275),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_304),
.A2(n_316),
.B1(n_324),
.B2(n_280),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_279),
.B(n_240),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_305),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_260),
.B1(n_268),
.B2(n_240),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_325),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_276),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_310),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_282),
.A2(n_284),
.B(n_301),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_321),
.B(n_299),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_282),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_314),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_270),
.B1(n_254),
.B2(n_269),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_323),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_241),
.Y(n_322)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_292),
.B(n_259),
.Y(n_323)
);

AOI22x1_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_283),
.B1(n_291),
.B2(n_286),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_258),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_284),
.B(n_264),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_327),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_281),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_242),
.B(n_250),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_277),
.C(n_275),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_339),
.C(n_340),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_336),
.A2(n_344),
.B1(n_313),
.B2(n_316),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_272),
.C(n_290),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_296),
.C(n_285),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_285),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_351),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_281),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_346),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_280),
.B1(n_299),
.B2(n_271),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_345),
.A2(n_317),
.B(n_327),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_271),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_349),
.A2(n_317),
.B1(n_324),
.B2(n_328),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_248),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_250),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_355),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_11),
.C(n_13),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_327),
.C(n_330),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_324),
.B1(n_353),
.B2(n_351),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_350),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_360),
.B(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_332),
.B(n_305),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_365),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_333),
.A2(n_322),
.B1(n_313),
.B2(n_321),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_355),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_367),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_334),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_368),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_338),
.A2(n_307),
.B1(n_320),
.B2(n_315),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_369),
.A2(n_377),
.B1(n_344),
.B2(n_309),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_315),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_370),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_310),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_375),
.Y(n_390)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_339),
.C(n_346),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g379 ( 
.A(n_358),
.B(n_341),
.CI(n_343),
.CON(n_379),
.SN(n_379)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_387),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_357),
.A2(n_345),
.B1(n_336),
.B2(n_352),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_383),
.A2(n_386),
.B1(n_377),
.B2(n_359),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_368),
.A2(n_304),
.B(n_342),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_392),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_391),
.A2(n_359),
.B1(n_365),
.B2(n_353),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_382),
.B(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_395),
.B(n_396),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_380),
.A2(n_369),
.B(n_375),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_390),
.A2(n_371),
.B(n_367),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_404),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g400 ( 
.A(n_381),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_402),
.Y(n_410)
);

OAI21x1_ASAP7_75t_SL g401 ( 
.A1(n_381),
.A2(n_384),
.B(n_388),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_389),
.B1(n_388),
.B2(n_394),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g402 ( 
.A(n_394),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_407),
.Y(n_411)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_371),
.C(n_392),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_414),
.C(n_416),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_378),
.C(n_383),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_391),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_386),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_378),
.C(n_366),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_418),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_366),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_419),
.B(n_363),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_425),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_422),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_347),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_409),
.Y(n_425)
);

NOR3xp33_ASAP7_75t_SL g426 ( 
.A(n_417),
.B(n_408),
.C(n_379),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_427),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_376),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_428),
.A2(n_393),
.B1(n_415),
.B2(n_414),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_429),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_413),
.B(n_393),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_423),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_335),
.C(n_379),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_420),
.C(n_411),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_435),
.A2(n_436),
.B(n_438),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_432),
.B(n_423),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_437),
.A2(n_433),
.B(n_430),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_439),
.C(n_411),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_441),
.A2(n_426),
.B(n_331),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_329),
.B(n_356),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_443),
.B(n_363),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_13),
.Y(n_445)
);


endmodule