module fake_ariane_693_n_2375 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2375);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2375;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_2370;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_1083;
wire n_337;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_307;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_261;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_348;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2275;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_133),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_154),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_112),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_98),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_155),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_71),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_4),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_66),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_89),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_27),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_59),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_83),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_191),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_87),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_164),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_15),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_22),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_138),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_66),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_11),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_69),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_27),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_73),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_121),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_38),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_189),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_177),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_65),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_152),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_102),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_68),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_127),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_74),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_209),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_62),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_59),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_173),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_25),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_117),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_130),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_111),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_162),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_113),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_44),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_158),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_11),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_149),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_187),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_13),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_166),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_201),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_174),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_9),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_219),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_90),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_95),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_142),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_23),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_94),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_69),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_157),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_50),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_143),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_35),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_19),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

BUFx2_ASAP7_75t_SL g305 ( 
.A(n_84),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_192),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_190),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_183),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_1),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_58),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_118),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_205),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_67),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_73),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_67),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_49),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_35),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_109),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_193),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_68),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_9),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_175),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_56),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_58),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_184),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_26),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_103),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_197),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_144),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_128),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_171),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_79),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_82),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_60),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_159),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_141),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_120),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_179),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_224),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_217),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_202),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_38),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_84),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_39),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_213),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_136),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_0),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_126),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_115),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_71),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_153),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_186),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_148),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_195),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_29),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_226),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_196),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_167),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_91),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_122),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_82),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_72),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_63),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_52),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_119),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_150),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_145),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_131),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_165),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_199),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_214),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_194),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_6),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_53),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_227),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_110),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_23),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_163),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_124),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_108),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_54),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_40),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_40),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_181),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_180),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_30),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_43),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_147),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_74),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_8),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_106),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_33),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_225),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_77),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_8),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_114),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_207),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_107),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_146),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_18),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_42),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_96),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_137),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_7),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_57),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_42),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_80),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_139),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_156),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_161),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_49),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_3),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_25),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_34),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_34),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_75),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_16),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_46),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_99),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_132),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_218),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_216),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_21),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_47),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_92),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_19),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_140),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_104),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_72),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_206),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_52),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_77),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_211),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_37),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_172),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_198),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_22),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_56),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_93),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_30),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_3),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_86),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_21),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_51),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_76),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_6),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_16),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_134),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_48),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_290),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_413),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_275),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_279),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_234),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_353),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_413),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_326),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_365),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_234),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_353),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_232),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_232),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_235),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_235),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_287),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_280),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_273),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_273),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_277),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_281),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_281),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_282),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_276),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_350),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_287),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_282),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_285),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_433),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_285),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_371),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_377),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_288),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_288),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_294),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_237),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_294),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_305),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_304),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_242),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_298),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_276),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_299),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_299),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_246),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_403),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_280),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_304),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_236),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_230),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_298),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_300),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_300),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_247),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_249),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_250),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_257),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_270),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_308),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_308),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_319),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_319),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_433),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_322),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_252),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_420),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_329),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_433),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_329),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_280),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_348),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_348),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_356),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_253),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_280),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_356),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_360),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_443),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_360),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_236),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_367),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_448),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_254),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_260),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_240),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_431),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_449),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_267),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_374),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_268),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_367),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_370),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_286),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_374),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_327),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_370),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_373),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_345),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_373),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_289),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_295),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_386),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_289),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_386),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_301),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_303),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_313),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_387),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_387),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_399),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_315),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_452),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_457),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_526),
.B(n_369),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_559),
.B(n_270),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_470),
.A2(n_427),
.B(n_399),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_470),
.B(n_437),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_472),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_511),
.B(n_431),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_461),
.B(n_238),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_552),
.A2(n_346),
.B1(n_363),
.B2(n_241),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_464),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_510),
.B(n_475),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_471),
.B(n_427),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_453),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_558),
.A2(n_388),
.B1(n_408),
.B2(n_309),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_471),
.B(n_432),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_472),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_492),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_454),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_472),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_512),
.A2(n_255),
.B1(n_263),
.B2(n_240),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_504),
.B(n_431),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_473),
.A2(n_441),
.B(n_432),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_497),
.B(n_501),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_504),
.B(n_431),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_456),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_455),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_555),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_519),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_467),
.Y(n_611)
);

OA21x2_ASAP7_75t_L g612 ( 
.A1(n_473),
.A2(n_444),
.B(n_441),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_486),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_527),
.A2(n_263),
.B1(n_265),
.B2(n_255),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_455),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_458),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_458),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_529),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_459),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_459),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_559),
.B(n_309),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_505),
.B(n_265),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_555),
.Y(n_625)
);

BUFx8_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_493),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_475),
.B(n_444),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_474),
.B(n_408),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_474),
.B(n_477),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_506),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_469),
.B(n_476),
.Y(n_632)
);

BUFx6f_ASAP7_75t_SL g633 ( 
.A(n_487),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_555),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_477),
.B(n_451),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_462),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_462),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_483),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_465),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_483),
.Y(n_641)
);

NOR2x1_ASAP7_75t_L g642 ( 
.A(n_478),
.B(n_327),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_478),
.B(n_451),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_490),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_345),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_465),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_503),
.B(n_415),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_522),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_522),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_575),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_479),
.B(n_450),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_531),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_468),
.A2(n_463),
.B1(n_466),
.B2(n_460),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_487),
.B(n_450),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_479),
.B(n_238),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_531),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_480),
.B(n_229),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_509),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_480),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_481),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_481),
.B(n_415),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_482),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_520),
.B(n_289),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_482),
.B(n_229),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_516),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_500),
.B(n_289),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_484),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_484),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_488),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_488),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_588),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_663),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_588),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_588),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_586),
.B(n_508),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_585),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_631),
.B(n_517),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_635),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_577),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_588),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_630),
.B(n_500),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_602),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_630),
.B(n_489),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_586),
.A2(n_491),
.B1(n_494),
.B2(n_489),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_602),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_663),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_663),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_586),
.B(n_518),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_602),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_602),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_611),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_651),
.B(n_528),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_663),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_663),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_611),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_668),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_585),
.A2(n_494),
.B1(n_495),
.B2(n_491),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_663),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_630),
.B(n_495),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_611),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_610),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_611),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_651),
.B(n_537),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_617),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_664),
.B(n_546),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_576),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_654),
.A2(n_498),
.B1(n_502),
.B2(n_496),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_668),
.B(n_533),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_617),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_667),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_617),
.Y(n_712)
);

BUFx6f_ASAP7_75t_SL g713 ( 
.A(n_579),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_600),
.A2(n_567),
.B1(n_564),
.B2(n_538),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_617),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_664),
.B(n_547),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_630),
.B(n_551),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_661),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_600),
.A2(n_549),
.B1(n_541),
.B2(n_545),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_667),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_633),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_662),
.B(n_543),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_592),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_661),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_576),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_580),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_661),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_614),
.A2(n_550),
.B1(n_557),
.B2(n_553),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_671),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_R g731 ( 
.A(n_597),
.B(n_565),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_654),
.A2(n_498),
.B1(n_502),
.B2(n_496),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_668),
.B(n_513),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_671),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_601),
.B(n_569),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_644),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_644),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_671),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_601),
.B(n_570),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_583),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_592),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_598),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_660),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_606),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_660),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_581),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_598),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_668),
.B(n_669),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_608),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_669),
.B(n_513),
.Y(n_751)
);

NOR2x1p5_ASAP7_75t_L g752 ( 
.A(n_623),
.B(n_548),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_624),
.B(n_623),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_608),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_615),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_629),
.A2(n_515),
.B1(n_521),
.B2(n_514),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_670),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_670),
.B(n_514),
.Y(n_758)
);

AOI21x1_ASAP7_75t_L g759 ( 
.A1(n_615),
.A2(n_521),
.B(n_515),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_578),
.B(n_571),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_606),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_616),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_624),
.B(n_499),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_662),
.B(n_523),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_616),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_582),
.B(n_666),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_618),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_618),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_629),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_662),
.B(n_523),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_620),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_620),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_582),
.B(n_524),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_621),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_621),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_629),
.B(n_524),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_637),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_629),
.B(n_525),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_636),
.B(n_525),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_638),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_638),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_640),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_640),
.B(n_530),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_647),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_590),
.B(n_507),
.Y(n_786)
);

XOR2xp5_ASAP7_75t_L g787 ( 
.A(n_619),
.B(n_317),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_579),
.B(n_530),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_581),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_578),
.B(n_532),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_647),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_636),
.B(n_643),
.Y(n_792)
);

NOR2x1p5_ASAP7_75t_L g793 ( 
.A(n_626),
.B(n_278),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_639),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_639),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_644),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_636),
.B(n_532),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_581),
.Y(n_798)
);

NOR2x1p5_ASAP7_75t_L g799 ( 
.A(n_626),
.B(n_278),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_581),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_644),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_581),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_639),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_603),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_603),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_641),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_SL g807 ( 
.A(n_587),
.B(n_320),
.C(n_318),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_614),
.B(n_305),
.Y(n_808)
);

AOI21x1_ASAP7_75t_L g809 ( 
.A1(n_603),
.A2(n_535),
.B(n_534),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_659),
.Y(n_810)
);

INVx5_ASAP7_75t_L g811 ( 
.A(n_635),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_603),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_641),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_641),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_646),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_595),
.A2(n_652),
.B(n_658),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_636),
.A2(n_535),
.B1(n_536),
.B2(n_534),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_646),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_643),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_603),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_594),
.A2(n_376),
.B1(n_328),
.B2(n_334),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_646),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_584),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_612),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_612),
.Y(n_825)
);

CKINVDCx6p67_ASAP7_75t_R g826 ( 
.A(n_633),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_644),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_584),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_662),
.B(n_536),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_612),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_633),
.B(n_539),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_612),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_644),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_SL g834 ( 
.A(n_680),
.B(n_632),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_790),
.B(n_648),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_707),
.B(n_658),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_725),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_760),
.B(n_677),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_721),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_723),
.B(n_648),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_721),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_807),
.A2(n_752),
.B1(n_808),
.B2(n_769),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_725),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_744),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_742),
.B(n_769),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_676),
.B(n_632),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_808),
.A2(n_587),
.B1(n_665),
.B2(n_594),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_697),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_707),
.B(n_665),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_725),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_689),
.B(n_593),
.Y(n_851)
);

BUFx6f_ASAP7_75t_SL g852 ( 
.A(n_721),
.Y(n_852)
);

BUFx5_ASAP7_75t_L g853 ( 
.A(n_798),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_753),
.B(n_645),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_766),
.B(n_706),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_819),
.B(n_628),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_707),
.B(n_747),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_744),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_726),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_726),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_726),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_746),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_731),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_819),
.B(n_655),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_716),
.B(n_633),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_753),
.B(n_607),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_752),
.A2(n_808),
.B1(n_816),
.B2(n_821),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_786),
.B(n_745),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_747),
.B(n_643),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_831),
.B(n_643),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_792),
.A2(n_652),
.B1(n_595),
.B2(n_336),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_786),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_685),
.B(n_604),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_579),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_711),
.B(n_579),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_746),
.Y(n_876)
);

BUFx5_ASAP7_75t_L g877 ( 
.A(n_798),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_720),
.B(n_622),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_747),
.B(n_626),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_747),
.B(n_626),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_757),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_789),
.B(n_622),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_709),
.B(n_613),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_720),
.A2(n_622),
.B1(n_642),
.B2(n_659),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_736),
.B(n_740),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_816),
.B(n_622),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_749),
.A2(n_612),
.B(n_589),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_728),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_697),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_693),
.B(n_627),
.C(n_302),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_721),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_757),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_697),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_697),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_765),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_702),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_745),
.B(n_659),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_765),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_728),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_704),
.B(n_302),
.C(n_297),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_816),
.B(n_645),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_698),
.B(n_642),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_684),
.B(n_700),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_728),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_764),
.B(n_539),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_771),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_734),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_773),
.A2(n_310),
.B(n_314),
.C(n_297),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_764),
.B(n_540),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_771),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_734),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_787),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_761),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_761),
.B(n_562),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_787),
.B(n_682),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_713),
.A2(n_656),
.B1(n_361),
.B2(n_262),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_770),
.B(n_540),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_734),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_770),
.B(n_542),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_775),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_775),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_808),
.A2(n_656),
.B1(n_544),
.B2(n_554),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_829),
.B(n_542),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_741),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_717),
.B(n_763),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_829),
.B(n_544),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_756),
.B(n_554),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_817),
.B(n_556),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_810),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_741),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_776),
.B(n_556),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_808),
.B(n_562),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_741),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_779),
.B(n_780),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_743),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_789),
.B(n_560),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_801),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_743),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_777),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_777),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_797),
.B(n_560),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_722),
.B(n_561),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_678),
.B(n_325),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_801),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_722),
.B(n_561),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_713),
.A2(n_656),
.B1(n_262),
.B2(n_311),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_793),
.B(n_563),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_782),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_782),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_708),
.B(n_562),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_743),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_732),
.B(n_563),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_826),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_785),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_713),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_748),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_733),
.B(n_566),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_748),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_810),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_748),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_785),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_789),
.B(n_566),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_791),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_791),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_789),
.B(n_824),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_751),
.B(n_568),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_824),
.B(n_750),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_713),
.A2(n_656),
.B1(n_572),
.B2(n_573),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_701),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_824),
.B(n_568),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_758),
.B(n_572),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_810),
.B(n_344),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_793),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_788),
.B(n_573),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_701),
.B(n_574),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_784),
.B(n_729),
.C(n_712),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_705),
.B(n_574),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_705),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_824),
.B(n_243),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_750),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_750),
.B(n_243),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_712),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_799),
.B(n_754),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_697),
.A2(n_656),
.B1(n_400),
.B2(n_311),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_799),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_754),
.B(n_400),
.Y(n_986)
);

AOI22x1_ASAP7_75t_L g987 ( 
.A1(n_754),
.A2(n_314),
.B1(n_316),
.B2(n_310),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_L g988 ( 
.A(n_800),
.B(n_656),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_715),
.B(n_364),
.C(n_357),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_755),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_800),
.B(n_656),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_714),
.B(n_316),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_826),
.B(n_366),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_719),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_718),
.B(n_323),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_755),
.B(n_274),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_715),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_672),
.B(n_656),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_672),
.B(n_231),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_755),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_L g1001 ( 
.A(n_802),
.B(n_379),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_672),
.B(n_674),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_801),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_762),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_762),
.B(n_274),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_762),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_718),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_674),
.B(n_272),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_802),
.B(n_383),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_937),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_838),
.B(n_687),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_L g1012 ( 
.A(n_863),
.B(n_724),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_837),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_863),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_854),
.B(n_724),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_947),
.B(n_767),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_853),
.B(n_767),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_SL g1018 ( 
.A(n_883),
.B(n_385),
.C(n_384),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_953),
.B(n_727),
.Y(n_1019)
);

INVx8_ASAP7_75t_L g1020 ( 
.A(n_852),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_835),
.B(n_767),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_847),
.A2(n_772),
.B1(n_774),
.B2(n_768),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_896),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_953),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_844),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_L g1026 ( 
.A(n_866),
.B(n_727),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_846),
.B(n_687),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_840),
.B(n_768),
.Y(n_1028)
);

AND2x6_ASAP7_75t_L g1029 ( 
.A(n_983),
.B(n_804),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_937),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_856),
.B(n_768),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_858),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_947),
.B(n_772),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_872),
.B(n_730),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_853),
.B(n_772),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_862),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_889),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_852),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_845),
.A2(n_778),
.B1(n_781),
.B2(n_774),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_876),
.Y(n_1040)
);

AND2x6_ASAP7_75t_SL g1041 ( 
.A(n_943),
.B(n_323),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_864),
.B(n_774),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_929),
.B(n_687),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_932),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_881),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_942),
.B(n_945),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_852),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_868),
.B(n_730),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_873),
.B(n_687),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_905),
.B(n_778),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_892),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_895),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_947),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_898),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_965),
.A2(n_781),
.B(n_778),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_837),
.Y(n_1056)
);

AO22x1_ASAP7_75t_L g1057 ( 
.A1(n_994),
.A2(n_391),
.B1(n_396),
.B2(n_389),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_992),
.A2(n_783),
.B1(n_781),
.B2(n_739),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_909),
.B(n_783),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_SL g1060 ( 
.A1(n_994),
.A2(n_402),
.B1(n_406),
.B2(n_397),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_917),
.B(n_783),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_973),
.B(n_674),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_929),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_843),
.Y(n_1064)
);

AND2x4_ASAP7_75t_SL g1065 ( 
.A(n_955),
.B(n_292),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_937),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_919),
.B(n_735),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_914),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_906),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_891),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_843),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_912),
.A2(n_409),
.B1(n_414),
.B2(n_407),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_850),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_903),
.A2(n_920),
.B1(n_921),
.B2(n_910),
.Y(n_1075)
);

CKINVDCx8_ASAP7_75t_R g1076 ( 
.A(n_993),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_939),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_940),
.A2(n_739),
.B(n_735),
.C(n_804),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_867),
.A2(n_812),
.B1(n_820),
.B2(n_805),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_897),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_937),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_923),
.B(n_675),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_944),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_889),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_842),
.A2(n_447),
.B1(n_442),
.B2(n_440),
.C(n_439),
.Y(n_1085)
);

AND2x6_ASAP7_75t_SL g1086 ( 
.A(n_885),
.B(n_335),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_948),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_850),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_949),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_954),
.A2(n_694),
.B(n_675),
.C(n_683),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_926),
.B(n_675),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_961),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_934),
.B(n_681),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_891),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_834),
.B(n_809),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_859),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_963),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_915),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_944),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_950),
.B(n_681),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_944),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_965),
.A2(n_688),
.B(n_673),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_944),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_964),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_913),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_925),
.B(n_694),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_969),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_952),
.B(n_681),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_855),
.A2(n_694),
.B1(n_688),
.B2(n_673),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_966),
.B(n_683),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_978),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_890),
.B(n_900),
.C(n_851),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_874),
.B(n_809),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1003),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_972),
.B(n_425),
.C(n_418),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_976),
.A2(n_812),
.B(n_820),
.C(n_805),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_853),
.B(n_877),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_989),
.B(n_436),
.C(n_426),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_882),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_859),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1003),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_901),
.B(n_694),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_875),
.B(n_683),
.Y(n_1123)
);

INVxp33_ASAP7_75t_L g1124 ( 
.A(n_865),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_971),
.B(n_931),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_853),
.B(n_686),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_983),
.B(n_686),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_990),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_990),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_982),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1003),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_985),
.B(n_686),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_853),
.B(n_690),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_997),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_878),
.B(n_690),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1007),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_860),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_983),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_902),
.A2(n_335),
.B1(n_352),
.B2(n_349),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_870),
.B(n_690),
.Y(n_1140)
);

AND2x6_ASAP7_75t_SL g1141 ( 
.A(n_995),
.B(n_349),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_975),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_941),
.B(n_691),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_839),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_886),
.A2(n_830),
.B1(n_832),
.B2(n_825),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_839),
.B(n_691),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_977),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_860),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_841),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_861),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_927),
.B(n_691),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_928),
.B(n_692),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_861),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_888),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_SL g1155 ( 
.A1(n_922),
.A2(n_375),
.B1(n_392),
.B2(n_352),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_841),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_888),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_879),
.A2(n_695),
.B1(n_699),
.B2(n_825),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_899),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_899),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_904),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1000),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_853),
.B(n_692),
.Y(n_1163)
);

XOR2x2_ASAP7_75t_L g1164 ( 
.A(n_879),
.B(n_375),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_957),
.B(n_692),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_904),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_880),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_907),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_853),
.B(n_696),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_999),
.Y(n_1170)
);

BUFx4_ASAP7_75t_L g1171 ( 
.A(n_1008),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_877),
.B(n_696),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_907),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_911),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_974),
.B(n_696),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_911),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_918),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_918),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_877),
.B(n_703),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1000),
.B(n_703),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1006),
.B(n_703),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1009),
.A2(n_434),
.B1(n_445),
.B2(n_446),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_880),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_924),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_848),
.Y(n_1185)
);

BUFx4f_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

INVx8_ASAP7_75t_L g1187 ( 
.A(n_882),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_924),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_848),
.B(n_710),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_893),
.B(n_710),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_877),
.B(n_710),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_930),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_871),
.B(n_830),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_877),
.B(n_695),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_930),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_869),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_893),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_933),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_877),
.B(n_699),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1001),
.A2(n_832),
.B1(n_818),
.B2(n_794),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_933),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_884),
.B(n_869),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_987),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_894),
.B(n_737),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1025),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1018),
.A2(n_849),
.B(n_836),
.C(n_1001),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1064),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1046),
.B(n_935),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1023),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1117),
.A2(n_967),
.B(n_988),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1171),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1117),
.A2(n_967),
.B(n_988),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1125),
.B(n_935),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1080),
.A2(n_849),
.B(n_836),
.C(n_1009),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_R g1215 ( 
.A(n_1024),
.B(n_759),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1017),
.A2(n_991),
.B(n_894),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1020),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_L g1218 ( 
.A(n_1112),
.B(n_394),
.C(n_392),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1026),
.A2(n_991),
.B1(n_959),
.B2(n_857),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_1023),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1014),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1186),
.B(n_877),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1017),
.A2(n_979),
.B(n_857),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_SL g1224 ( 
.A(n_1071),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1142),
.B(n_938),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1035),
.A2(n_1021),
.B(n_1031),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1060),
.A2(n_908),
.B1(n_445),
.B2(n_434),
.C(n_428),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_1030),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_L g1229 ( 
.A(n_1071),
.B(n_1094),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1098),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1032),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1030),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1076),
.B(n_292),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1105),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1147),
.B(n_938),
.Y(n_1235)
);

BUFx8_ASAP7_75t_SL g1236 ( 
.A(n_1038),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1080),
.B(n_951),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1044),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1035),
.A2(n_979),
.B(n_887),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1057),
.A2(n_416),
.B1(n_417),
.B2(n_394),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1011),
.B(n_951),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1124),
.B(n_936),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1053),
.A2(n_936),
.B1(n_970),
.B2(n_962),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1044),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1075),
.A2(n_1059),
.B1(n_1061),
.B2(n_1050),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1124),
.B(n_962),
.Y(n_1246)
);

NAND2xp33_ASAP7_75t_SL g1247 ( 
.A(n_1118),
.B(n_970),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1016),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1042),
.A2(n_1002),
.B(n_958),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1115),
.A2(n_986),
.B(n_981),
.C(n_417),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1028),
.A2(n_958),
.B(n_956),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1010),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1036),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1040),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1045),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1011),
.A2(n_986),
.B(n_981),
.C(n_419),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1027),
.B(n_956),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1027),
.B(n_960),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1182),
.B(n_419),
.C(n_416),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1106),
.B(n_960),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1093),
.A2(n_1004),
.B(n_980),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1051),
.Y(n_1262)
);

INVx3_ASAP7_75t_SL g1263 ( 
.A(n_1047),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1030),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1049),
.A2(n_1004),
.B(n_980),
.Y(n_1265)
);

OAI221xp5_ASAP7_75t_L g1266 ( 
.A1(n_1085),
.A2(n_916),
.B1(n_984),
.B2(n_428),
.C(n_446),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1016),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1106),
.B(n_968),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1052),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1094),
.B(n_292),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1186),
.B(n_946),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1194),
.A2(n_998),
.B(n_996),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1170),
.B(n_737),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1064),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_SL g1275 ( 
.A(n_1182),
.B(n_1118),
.C(n_1167),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1015),
.B(n_996),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1020),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1029),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1054),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1034),
.B(n_1005),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1194),
.A2(n_1005),
.B(n_738),
.Y(n_1281)
);

AO32x2_ASAP7_75t_L g1282 ( 
.A1(n_1155),
.A2(n_759),
.A3(n_803),
.B1(n_794),
.B2(n_795),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1073),
.B(n_233),
.C(n_228),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1199),
.A2(n_1133),
.B(n_1126),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1048),
.B(n_292),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1065),
.A2(n_393),
.B1(n_395),
.B2(n_296),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1033),
.B(n_801),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1067),
.A2(n_796),
.B1(n_738),
.B2(n_827),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1199),
.A2(n_796),
.B(n_738),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1041),
.B(n_738),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1088),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1088),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1068),
.B(n_827),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1010),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1086),
.B(n_801),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1070),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1122),
.B(n_794),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1141),
.B(n_833),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1020),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1149),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1019),
.B(n_393),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1133),
.A2(n_833),
.B(n_828),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1058),
.B(n_1128),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1029),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1058),
.B(n_795),
.Y(n_1305)
);

INVx3_ASAP7_75t_SL g1306 ( 
.A(n_1065),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1055),
.A2(n_828),
.B(n_823),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1128),
.B(n_795),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1164),
.B(n_393),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_1022),
.B(n_833),
.C(n_381),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1149),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1029),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1129),
.B(n_803),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1132),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1166),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1140),
.A2(n_828),
.B(n_823),
.C(n_284),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1029),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1012),
.B(n_833),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1140),
.A2(n_284),
.B(n_381),
.C(n_818),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1022),
.A2(n_803),
.B1(n_822),
.B2(n_818),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1129),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1138),
.B(n_833),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1119),
.A2(n_833),
.B1(n_412),
.B2(n_372),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1077),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_R g1325 ( 
.A(n_1144),
.B(n_239),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1087),
.B(n_393),
.Y(n_1326)
);

INVx3_ASAP7_75t_SL g1327 ( 
.A(n_1144),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1089),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1144),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1166),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1144),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1119),
.A2(n_822),
.B(n_815),
.C(n_814),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1013),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1163),
.A2(n_813),
.B(n_806),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1156),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1158),
.A2(n_813),
.B(n_806),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1162),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1163),
.A2(n_813),
.B(n_806),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1162),
.B(n_814),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1156),
.B(n_244),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1092),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1196),
.A2(n_822),
.B(n_815),
.C(n_814),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1097),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1104),
.B(n_815),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1010),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1169),
.A2(n_811),
.B(n_679),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1145),
.B(n_679),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_SL g1348 ( 
.A1(n_1107),
.A2(n_609),
.B(n_589),
.C(n_591),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_1156),
.B(n_245),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1111),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_SL g1351 ( 
.A(n_1183),
.B(n_339),
.C(n_251),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1156),
.B(n_248),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1132),
.B(n_256),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1145),
.B(n_679),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1062),
.B(n_679),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1169),
.A2(n_811),
.B(n_679),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1062),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1063),
.B(n_679),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1010),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1066),
.Y(n_1360)
);

AO32x1_ASAP7_75t_L g1361 ( 
.A1(n_1203),
.A2(n_653),
.A3(n_649),
.B1(n_591),
.B2(n_596),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1196),
.B(n_258),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1202),
.A2(n_1136),
.B1(n_1193),
.B2(n_1134),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1095),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1100),
.B(n_811),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1081),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1029),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_SL g1368 ( 
.A1(n_1172),
.A2(n_584),
.B(n_589),
.C(n_591),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1245),
.A2(n_1241),
.B(n_1257),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1238),
.B(n_1130),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1333),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1304),
.B(n_1081),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1244),
.B(n_1127),
.Y(n_1373)
);

AO32x2_ASAP7_75t_L g1374 ( 
.A1(n_1363),
.A2(n_1039),
.A3(n_1185),
.B1(n_1090),
.B2(n_1139),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1327),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1245),
.A2(n_1159),
.B(n_1116),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1209),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1241),
.A2(n_1179),
.B(n_1172),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1307),
.A2(n_1102),
.B(n_1179),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_SL g1380 ( 
.A1(n_1214),
.A2(n_1109),
.B(n_1185),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1257),
.A2(n_1191),
.B(n_1165),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1363),
.A2(n_1213),
.B1(n_1208),
.B2(n_1242),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_SL g1383 ( 
.A(n_1233),
.B(n_261),
.C(n_259),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1258),
.A2(n_1191),
.B(n_1078),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1239),
.A2(n_1200),
.B(n_1108),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1220),
.B(n_1127),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1205),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1218),
.B(n_1078),
.C(n_1082),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1206),
.A2(n_1187),
.B(n_1110),
.C(n_1091),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1226),
.A2(n_1113),
.B(n_1116),
.Y(n_1390)
);

AO32x2_ASAP7_75t_L g1391 ( 
.A1(n_1288),
.A2(n_1320),
.A3(n_1282),
.B1(n_1357),
.B2(n_1361),
.Y(n_1391)
);

AO32x2_ASAP7_75t_L g1392 ( 
.A1(n_1288),
.A2(n_1320),
.A3(n_1282),
.B1(n_1361),
.B2(n_1228),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_R g1393 ( 
.A(n_1311),
.B(n_1081),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1309),
.A2(n_1139),
.B(n_1200),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1304),
.B(n_1081),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1231),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1228),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1277),
.B(n_1099),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1321),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1284),
.A2(n_1152),
.B(n_1151),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1210),
.A2(n_1181),
.B(n_1180),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1236),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1237),
.A2(n_1143),
.B(n_1135),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1258),
.A2(n_1090),
.B(n_1069),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1260),
.A2(n_1123),
.B(n_1175),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1232),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1337),
.B(n_1079),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1300),
.B(n_1099),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1253),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1212),
.A2(n_1153),
.B(n_1148),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1297),
.A2(n_1178),
.A3(n_1201),
.B(n_1198),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1246),
.A2(n_1187),
.B(n_1159),
.C(n_1146),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1223),
.A2(n_1161),
.B(n_1157),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1207),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1260),
.A2(n_1069),
.B(n_1037),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1232),
.Y(n_1416)
);

O2A1O1Ixp5_ASAP7_75t_SL g1417 ( 
.A1(n_1318),
.A2(n_649),
.B(n_653),
.C(n_1340),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1254),
.Y(n_1418)
);

AOI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1268),
.A2(n_1187),
.B(n_1079),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1248),
.B(n_1174),
.Y(n_1420)
);

OAI22x1_ASAP7_75t_L g1421 ( 
.A1(n_1298),
.A2(n_1177),
.B1(n_1192),
.B2(n_1188),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1221),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1275),
.A2(n_1043),
.B(n_1204),
.C(n_1037),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1213),
.A2(n_1101),
.B(n_1083),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1285),
.B(n_1056),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1302),
.A2(n_1272),
.B(n_1261),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1314),
.B(n_1072),
.Y(n_1427)
);

NAND3x1_ASAP7_75t_L g1428 ( 
.A(n_1290),
.B(n_1084),
.C(n_0),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1255),
.Y(n_1429)
);

AO31x2_ASAP7_75t_L g1430 ( 
.A1(n_1297),
.A2(n_1074),
.A3(n_1096),
.B(n_1195),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_SL g1431 ( 
.A1(n_1276),
.A2(n_1137),
.B(n_1120),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1208),
.A2(n_1268),
.B1(n_1303),
.B2(n_1269),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1325),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1216),
.A2(n_1222),
.B(n_1249),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1252),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1265),
.A2(n_1190),
.B(n_1189),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1240),
.B(n_1326),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_SL g1438 ( 
.A(n_1304),
.B(n_1114),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1234),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1229),
.B(n_1083),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1334),
.A2(n_1154),
.B(n_1150),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1251),
.A2(n_1103),
.B(n_1066),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1230),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1338),
.A2(n_1168),
.B(n_1160),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1306),
.B(n_1146),
.Y(n_1445)
);

AO31x2_ASAP7_75t_L g1446 ( 
.A1(n_1319),
.A2(n_1173),
.A3(n_1176),
.B(n_1184),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1247),
.A2(n_1227),
.B(n_1250),
.C(n_1256),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1281),
.A2(n_1043),
.B(n_599),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1262),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1346),
.A2(n_599),
.B(n_596),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1362),
.B(n_1197),
.Y(n_1451)
);

NAND2xp33_ASAP7_75t_L g1452 ( 
.A(n_1215),
.B(n_1114),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1303),
.A2(n_1197),
.B1(n_1204),
.B2(n_1103),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_SL g1454 ( 
.A(n_1286),
.B(n_266),
.C(n_264),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1267),
.B(n_1101),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1273),
.B(n_1189),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1279),
.B(n_1190),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1263),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1225),
.B(n_1103),
.Y(n_1459)
);

AO31x2_ASAP7_75t_L g1460 ( 
.A1(n_1347),
.A2(n_625),
.A3(n_634),
.B(n_609),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1224),
.Y(n_1461)
);

BUFx10_ASAP7_75t_L g1462 ( 
.A(n_1224),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1266),
.A2(n_1197),
.B(n_1131),
.C(n_1121),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1310),
.A2(n_1295),
.B(n_1219),
.C(n_1259),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1274),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1356),
.A2(n_1121),
.B(n_1114),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1349),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1217),
.Y(n_1468)
);

AOI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1347),
.A2(n_609),
.B(n_605),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1289),
.A2(n_1365),
.B(n_1354),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1225),
.A2(n_1131),
.B(n_1121),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1264),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1354),
.A2(n_625),
.B(n_605),
.Y(n_1473)
);

AOI31xp67_ASAP7_75t_L g1474 ( 
.A1(n_1243),
.A2(n_634),
.A3(n_605),
.B(n_625),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1353),
.B(n_1296),
.Y(n_1475)
);

AO32x2_ASAP7_75t_L g1476 ( 
.A1(n_1282),
.A2(n_1361),
.A3(n_1264),
.B1(n_1366),
.B2(n_1299),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1305),
.A2(n_634),
.B(n_1197),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1351),
.A2(n_1),
.B(n_2),
.Y(n_1478)
);

BUFx10_ASAP7_75t_L g1479 ( 
.A(n_1331),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1235),
.B(n_1131),
.Y(n_1480)
);

BUFx4_ASAP7_75t_SL g1481 ( 
.A(n_1329),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1324),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1211),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1278),
.B(n_1131),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1335),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1235),
.B(n_650),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1291),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1316),
.A2(n_811),
.B(n_395),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1304),
.B(n_269),
.Y(n_1489)
);

OAI22x1_ASAP7_75t_L g1490 ( 
.A1(n_1328),
.A2(n_340),
.B1(n_338),
.B2(n_337),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1305),
.A2(n_811),
.B(n_657),
.Y(n_1491)
);

AO32x2_ASAP7_75t_L g1492 ( 
.A1(n_1366),
.A2(n_650),
.A3(n_657),
.B1(n_5),
.B2(n_10),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1292),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1341),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1342),
.A2(n_811),
.B(n_657),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1355),
.B(n_1312),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1308),
.A2(n_429),
.B(n_430),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1332),
.A2(n_657),
.B(n_650),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1308),
.A2(n_657),
.B(n_650),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1343),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1301),
.B(n_271),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1315),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1331),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1313),
.A2(n_429),
.B(n_430),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1283),
.B(n_657),
.C(n_650),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1276),
.A2(n_362),
.B(n_291),
.Y(n_1506)
);

AO31x2_ASAP7_75t_L g1507 ( 
.A1(n_1330),
.A2(n_650),
.A3(n_430),
.B(n_429),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1350),
.B(n_1364),
.Y(n_1508)
);

OAI21xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1313),
.A2(n_10),
.B(n_12),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1270),
.B(n_13),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1344),
.A2(n_358),
.B(n_438),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1339),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1252),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1339),
.A2(n_635),
.B(n_169),
.Y(n_1514)
);

NAND2x1_ASAP7_75t_L g1515 ( 
.A(n_1331),
.B(n_635),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1280),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1368),
.A2(n_430),
.B(n_435),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1352),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1293),
.B(n_14),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1355),
.B(n_14),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1323),
.B(n_15),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1252),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1271),
.A2(n_355),
.B(n_424),
.C(n_423),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1287),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1294),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1336),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1348),
.A2(n_430),
.B(n_422),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1294),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1294),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1322),
.A2(n_347),
.B(n_411),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1317),
.A2(n_421),
.B(n_410),
.C(n_405),
.Y(n_1531)
);

AO32x2_ASAP7_75t_L g1532 ( 
.A1(n_1336),
.A2(n_17),
.A3(n_20),
.B1(n_24),
.B2(n_26),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1367),
.B(n_17),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1358),
.B(n_1345),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1345),
.B(n_20),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1345),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1358),
.A2(n_404),
.B(n_401),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1359),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1359),
.A2(n_1360),
.B1(n_398),
.B2(n_390),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1359),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_R g1541 ( 
.A(n_1360),
.B(n_283),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1360),
.B(n_28),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1245),
.A2(n_382),
.B(n_380),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1220),
.B(n_31),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1205),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1363),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1304),
.B(n_88),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1370),
.B(n_32),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1473),
.A2(n_125),
.B(n_222),
.Y(n_1549)
);

AOI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1469),
.A2(n_378),
.B(n_368),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1394),
.A2(n_359),
.B1(n_354),
.B2(n_351),
.C(n_343),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1387),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1396),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_36),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_101),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1433),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1478),
.A2(n_342),
.B1(n_341),
.B2(n_333),
.C(n_332),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1409),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1418),
.Y(n_1559)
);

NAND2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1372),
.B(n_221),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1534),
.B(n_1496),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1394),
.A2(n_331),
.B(n_330),
.C(n_324),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1429),
.Y(n_1563)
);

CKINVDCx8_ASAP7_75t_R g1564 ( 
.A(n_1375),
.Y(n_1564)
);

CKINVDCx11_ASAP7_75t_R g1565 ( 
.A(n_1402),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1526),
.A2(n_1477),
.B(n_1431),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1426),
.A2(n_321),
.B(n_312),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1377),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1458),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1475),
.B(n_36),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1447),
.A2(n_307),
.B(n_306),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1499),
.A2(n_215),
.B(n_212),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1424),
.B(n_210),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1437),
.B(n_37),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1471),
.B(n_208),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1399),
.B(n_39),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1449),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1543),
.A2(n_293),
.B(n_43),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1451),
.B(n_41),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1375),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1513),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1496),
.B(n_204),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1481),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1513),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1462),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1491),
.A2(n_203),
.B(n_200),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1372),
.B(n_188),
.Y(n_1587)
);

NAND2x1p5_ASAP7_75t_L g1588 ( 
.A(n_1513),
.B(n_182),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1484),
.B(n_176),
.Y(n_1589)
);

AO21x2_ASAP7_75t_L g1590 ( 
.A1(n_1390),
.A2(n_151),
.B(n_135),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1508),
.B(n_41),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1546),
.A2(n_1478),
.B1(n_1500),
.B2(n_1538),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1470),
.A2(n_129),
.B(n_123),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1484),
.B(n_116),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1369),
.A2(n_105),
.B(n_100),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1373),
.B(n_45),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1390),
.A2(n_45),
.B(n_46),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1482),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1494),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1479),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1389),
.A2(n_48),
.B(n_50),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1479),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1382),
.B(n_51),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1546),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1388),
.A2(n_55),
.B(n_57),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1545),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1404),
.A2(n_60),
.B(n_61),
.Y(n_1607)
);

AO21x2_ASAP7_75t_L g1608 ( 
.A1(n_1403),
.A2(n_61),
.B(n_63),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1434),
.A2(n_1379),
.B(n_1514),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1460),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1484),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1385),
.A2(n_64),
.B(n_65),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1400),
.A2(n_64),
.B(n_70),
.Y(n_1613)
);

BUFx8_ASAP7_75t_L g1614 ( 
.A(n_1467),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1510),
.B(n_70),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1388),
.A2(n_75),
.B(n_76),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1414),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1407),
.B(n_78),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_SL g1619 ( 
.A1(n_1380),
.A2(n_78),
.B(n_79),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1461),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1420),
.B(n_80),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1384),
.A2(n_81),
.B(n_83),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1386),
.B(n_81),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1411),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1382),
.B(n_85),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1498),
.A2(n_85),
.B(n_1442),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1401),
.A2(n_1413),
.B(n_1410),
.Y(n_1627)
);

OR2x6_ASAP7_75t_L g1628 ( 
.A(n_1376),
.B(n_1453),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1453),
.B(n_1436),
.Y(n_1629)
);

AOI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1497),
.A2(n_1504),
.B(n_1466),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1411),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1465),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1487),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1452),
.A2(n_1381),
.B(n_1415),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1493),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_SL g1636 ( 
.A1(n_1500),
.A2(n_1538),
.B(n_1463),
.C(n_1464),
.Y(n_1636)
);

AOI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1421),
.A2(n_1506),
.B(n_1501),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1450),
.A2(n_1495),
.B(n_1448),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1393),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1439),
.B(n_1512),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1502),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1460),
.Y(n_1642)
);

CKINVDCx6p67_ASAP7_75t_R g1643 ( 
.A(n_1468),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1371),
.Y(n_1644)
);

NAND2xp33_ASAP7_75t_R g1645 ( 
.A(n_1506),
.B(n_1537),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1519),
.A2(n_1544),
.B1(n_1521),
.B2(n_1511),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1540),
.B(n_1435),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1457),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1511),
.A2(n_1530),
.B(n_1505),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1422),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1441),
.A2(n_1444),
.B(n_1378),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1435),
.B(n_1528),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1411),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1459),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1533),
.B(n_1485),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1459),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1432),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_1518),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1425),
.B(n_1432),
.Y(n_1659)
);

NAND2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1472),
.B(n_1398),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1509),
.A2(n_1490),
.B1(n_1454),
.B2(n_1383),
.C(n_1419),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1445),
.B(n_1456),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1520),
.B(n_1427),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1524),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1455),
.B(n_1398),
.Y(n_1665)
);

AOI31xp67_ASAP7_75t_L g1666 ( 
.A1(n_1486),
.A2(n_1480),
.A3(n_1489),
.B(n_1535),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1462),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1443),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1460),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1480),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1419),
.B(n_1542),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1509),
.A2(n_1483),
.B1(n_1405),
.B2(n_1537),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1412),
.B(n_1530),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1446),
.Y(n_1674)
);

OAI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1417),
.A2(n_1436),
.B(n_1517),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1405),
.A2(n_1541),
.B1(n_1505),
.B2(n_1488),
.Y(n_1676)
);

O2A1O1Ixp33_ASAP7_75t_SL g1677 ( 
.A1(n_1423),
.A2(n_1523),
.B(n_1531),
.C(n_1515),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1488),
.A2(n_1527),
.B(n_1547),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1428),
.A2(n_1539),
.B1(n_1416),
.B2(n_1406),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1529),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1539),
.A2(n_1406),
.B1(n_1416),
.B2(n_1397),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1446),
.Y(n_1682)
);

OA21x2_ASAP7_75t_L g1683 ( 
.A1(n_1474),
.A2(n_1374),
.B(n_1476),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1532),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1446),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1547),
.B(n_1408),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1397),
.A2(n_1507),
.B(n_1374),
.Y(n_1687)
);

AO31x2_ASAP7_75t_L g1688 ( 
.A1(n_1374),
.A2(n_1391),
.A3(n_1476),
.B(n_1392),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1507),
.A2(n_1395),
.B(n_1392),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1507),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1503),
.A2(n_1395),
.B(n_1440),
.C(n_1492),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1476),
.A2(n_1392),
.B(n_1391),
.Y(n_1692)
);

INVx6_ASAP7_75t_L g1693 ( 
.A(n_1472),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1438),
.A2(n_1391),
.B(n_1532),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1528),
.B(n_1536),
.Y(n_1695)
);

OA21x2_ASAP7_75t_L g1696 ( 
.A1(n_1532),
.A2(n_1492),
.B(n_1440),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1492),
.A2(n_1472),
.B(n_1522),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1528),
.A2(n_1536),
.B(n_1522),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1536),
.Y(n_1699)
);

AOI221x1_ASAP7_75t_L g1700 ( 
.A1(n_1525),
.A2(n_1546),
.B1(n_1538),
.B2(n_1500),
.C(n_1247),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1525),
.A2(n_1473),
.B(n_1469),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1387),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1513),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1546),
.A2(n_1309),
.B1(n_614),
.B2(n_600),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1478),
.B(n_883),
.C(n_1546),
.Y(n_1706)
);

INVxp67_ASAP7_75t_SL g1707 ( 
.A(n_1526),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1534),
.B(n_1496),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1394),
.A2(n_838),
.B(n_1478),
.C(n_1447),
.Y(n_1709)
);

AO31x2_ASAP7_75t_L g1710 ( 
.A1(n_1526),
.A2(n_1432),
.A3(n_1421),
.B(n_1369),
.Y(n_1710)
);

AO31x2_ASAP7_75t_L g1711 ( 
.A1(n_1526),
.A2(n_1432),
.A3(n_1421),
.B(n_1369),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1516),
.B(n_1377),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1394),
.B(n_883),
.Y(n_1713)
);

OAI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1394),
.A2(n_834),
.B1(n_1309),
.B2(n_883),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1430),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1394),
.A2(n_808),
.B1(n_1546),
.B2(n_1478),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1387),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1387),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1369),
.A2(n_1245),
.B(n_1117),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1447),
.A2(n_838),
.B1(n_1080),
.B2(n_1394),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1370),
.B(n_1238),
.Y(n_1724)
);

AO21x2_ASAP7_75t_L g1725 ( 
.A1(n_1526),
.A2(n_1469),
.B(n_1477),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1726)
);

OAI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1387),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1370),
.B(n_1238),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1730)
);

BUFx8_ASAP7_75t_L g1731 ( 
.A(n_1375),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_L g1732 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1430),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1387),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1426),
.A2(n_1473),
.B(n_1470),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1394),
.A2(n_838),
.B(n_1478),
.C(n_1447),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1458),
.Y(n_1737)
);

CKINVDCx11_ASAP7_75t_R g1738 ( 
.A(n_1402),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1513),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1481),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1513),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1473),
.A2(n_1469),
.B(n_1426),
.Y(n_1742)
);

OAI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1447),
.A2(n_838),
.B(n_883),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1426),
.A2(n_1473),
.B(n_1470),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1722),
.A2(n_1657),
.B(n_1713),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1657),
.A2(n_1713),
.B(n_1743),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1709),
.A2(n_1736),
.B(n_1723),
.C(n_1625),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1639),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1724),
.B(n_1729),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1712),
.B(n_1568),
.Y(n_1750)
);

OA21x2_ASAP7_75t_L g1751 ( 
.A1(n_1689),
.A2(n_1714),
.B(n_1703),
.Y(n_1751)
);

O2A1O1Ixp5_ASAP7_75t_L g1752 ( 
.A1(n_1625),
.A2(n_1718),
.B(n_1592),
.C(n_1601),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1717),
.A2(n_1726),
.B(n_1720),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1705),
.A2(n_1706),
.B1(n_1709),
.B2(n_1736),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1718),
.Y(n_1755)
);

AND2x4_ASAP7_75t_SL g1756 ( 
.A(n_1584),
.B(n_1561),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1562),
.A2(n_1575),
.B(n_1573),
.Y(n_1757)
);

OA21x2_ASAP7_75t_L g1758 ( 
.A1(n_1727),
.A2(n_1732),
.B(n_1730),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1562),
.A2(n_1673),
.B(n_1705),
.C(n_1578),
.Y(n_1759)
);

A2O1A1Ixp33_ASAP7_75t_SL g1760 ( 
.A1(n_1605),
.A2(n_1616),
.B(n_1603),
.C(n_1649),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1655),
.B(n_1615),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1640),
.B(n_1568),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1610),
.Y(n_1764)
);

BUFx4f_ASAP7_75t_SL g1765 ( 
.A(n_1731),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1731),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_L g1768 ( 
.A(n_1585),
.B(n_1600),
.Y(n_1768)
);

O2A1O1Ixp5_ASAP7_75t_L g1769 ( 
.A1(n_1592),
.A2(n_1604),
.B(n_1673),
.C(n_1646),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1731),
.Y(n_1770)
);

AOI21x1_ASAP7_75t_SL g1771 ( 
.A1(n_1576),
.A2(n_1548),
.B(n_1570),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1691),
.A2(n_1579),
.B(n_1671),
.C(n_1676),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1575),
.A2(n_1573),
.B(n_1589),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1552),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1575),
.A2(n_1573),
.B(n_1589),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1663),
.B(n_1659),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1579),
.B(n_1561),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1648),
.B(n_1670),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1610),
.Y(n_1779)
);

AOI21x1_ASAP7_75t_SL g1780 ( 
.A1(n_1591),
.A2(n_1596),
.B(n_1652),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1604),
.A2(n_1636),
.B(n_1557),
.C(n_1571),
.Y(n_1781)
);

NOR2xp67_ASAP7_75t_L g1782 ( 
.A(n_1600),
.B(n_1602),
.Y(n_1782)
);

AOI21x1_ASAP7_75t_SL g1783 ( 
.A1(n_1652),
.A2(n_1647),
.B(n_1594),
.Y(n_1783)
);

OA21x2_ASAP7_75t_L g1784 ( 
.A1(n_1742),
.A2(n_1609),
.B(n_1627),
.Y(n_1784)
);

O2A1O1Ixp5_ASAP7_75t_L g1785 ( 
.A1(n_1679),
.A2(n_1637),
.B(n_1671),
.C(n_1681),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1580),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1676),
.A2(n_1551),
.B1(n_1628),
.B2(n_1661),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1708),
.B(n_1665),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1662),
.B(n_1654),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1589),
.A2(n_1594),
.B(n_1582),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1656),
.B(n_1618),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1658),
.A2(n_1583),
.B1(n_1740),
.B2(n_1650),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_R g1793 ( 
.A(n_1564),
.B(n_1658),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1594),
.A2(n_1582),
.B(n_1597),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1553),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1558),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1559),
.B(n_1563),
.Y(n_1797)
);

AOI21x1_ASAP7_75t_SL g1798 ( 
.A1(n_1647),
.A2(n_1582),
.B(n_1555),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1634),
.A2(n_1636),
.B(n_1628),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1577),
.B(n_1598),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1599),
.B(n_1606),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1702),
.B(n_1719),
.Y(n_1802)
);

OA21x2_ASAP7_75t_L g1803 ( 
.A1(n_1651),
.A2(n_1687),
.B(n_1694),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1556),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1721),
.B(n_1728),
.Y(n_1805)
);

O2A1O1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1619),
.A2(n_1677),
.B(n_1554),
.C(n_1621),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_SL g1807 ( 
.A1(n_1597),
.A2(n_1700),
.B(n_1595),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1734),
.B(n_1664),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1629),
.B(n_1680),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1647),
.B(n_1699),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1672),
.B(n_1617),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1672),
.B(n_1632),
.Y(n_1812)
);

AOI21x1_ASAP7_75t_SL g1813 ( 
.A1(n_1555),
.A2(n_1643),
.B(n_1642),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1695),
.B(n_1698),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1698),
.B(n_1696),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1597),
.A2(n_1645),
.B1(n_1622),
.B2(n_1677),
.C(n_1595),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1633),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1611),
.B(n_1697),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1698),
.Y(n_1819)
);

AOI21x1_ASAP7_75t_SL g1820 ( 
.A1(n_1555),
.A2(n_1642),
.B(n_1669),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1614),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1614),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1635),
.Y(n_1823)
);

AOI21x1_ASAP7_75t_SL g1824 ( 
.A1(n_1669),
.A2(n_1607),
.B(n_1738),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1684),
.A2(n_1612),
.B(n_1678),
.C(n_1675),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1696),
.B(n_1644),
.Y(n_1826)
);

AOI21x1_ASAP7_75t_SL g1827 ( 
.A1(n_1607),
.A2(n_1738),
.B(n_1565),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1608),
.A2(n_1622),
.B(n_1595),
.C(n_1590),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1696),
.B(n_1611),
.Y(n_1829)
);

CKINVDCx16_ASAP7_75t_R g1830 ( 
.A(n_1668),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1611),
.B(n_1602),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1641),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1667),
.A2(n_1668),
.B1(n_1622),
.B2(n_1650),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1692),
.B(n_1688),
.Y(n_1834)
);

BUFx4f_ASAP7_75t_SL g1835 ( 
.A(n_1614),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1584),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1588),
.A2(n_1686),
.B(n_1560),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1667),
.A2(n_1692),
.B1(n_1620),
.B2(n_1737),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1584),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1581),
.B(n_1704),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1710),
.B(n_1711),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1624),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1588),
.A2(n_1686),
.B(n_1560),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1692),
.B(n_1688),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1688),
.B(n_1704),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1688),
.B(n_1739),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1581),
.B(n_1739),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1565),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1710),
.B(n_1711),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1741),
.B(n_1608),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1741),
.B(n_1660),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1569),
.Y(n_1852)
);

NOR2xp67_ASAP7_75t_L g1853 ( 
.A(n_1624),
.B(n_1631),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1660),
.B(n_1711),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1612),
.A2(n_1593),
.B(n_1653),
.C(n_1631),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1710),
.B(n_1711),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1710),
.B(n_1653),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1683),
.B(n_1716),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1569),
.Y(n_1859)
);

AOI21x1_ASAP7_75t_SL g1860 ( 
.A1(n_1620),
.A2(n_1567),
.B(n_1645),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1613),
.B(n_1693),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1613),
.B(n_1683),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1613),
.Y(n_1863)
);

OA21x2_ASAP7_75t_L g1864 ( 
.A1(n_1690),
.A2(n_1701),
.B(n_1682),
.Y(n_1864)
);

O2A1O1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1567),
.A2(n_1587),
.B(n_1683),
.C(n_1674),
.Y(n_1865)
);

A2O1A1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1586),
.A2(n_1626),
.B(n_1572),
.C(n_1549),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1707),
.B(n_1587),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1674),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1682),
.A2(n_1685),
.B(n_1733),
.C(n_1690),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1566),
.B(n_1685),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1550),
.A2(n_1744),
.B1(n_1735),
.B2(n_1630),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1638),
.A2(n_1707),
.B(n_1566),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1725),
.A2(n_1722),
.B(n_1657),
.Y(n_1873)
);

BUFx4f_ASAP7_75t_L g1874 ( 
.A(n_1666),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1725),
.Y(n_1875)
);

AOI21x1_ASAP7_75t_SL g1876 ( 
.A1(n_1603),
.A2(n_1576),
.B(n_1544),
.Y(n_1876)
);

BUFx4_ASAP7_75t_R g1877 ( 
.A(n_1628),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1724),
.B(n_1729),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1552),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_SL g1881 ( 
.A1(n_1709),
.A2(n_1736),
.B(n_1713),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1611),
.B(n_1561),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1698),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1722),
.A2(n_1657),
.B(n_1713),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1709),
.A2(n_1736),
.B(n_1713),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1724),
.B(n_1729),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1610),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1552),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1713),
.A2(n_1705),
.B1(n_1706),
.B2(n_1709),
.Y(n_1890)
);

A2O1A1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1713),
.A2(n_1709),
.B(n_1736),
.C(n_1743),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1713),
.A2(n_1705),
.B1(n_1706),
.B2(n_1709),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1713),
.A2(n_1705),
.B1(n_1706),
.B2(n_1709),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1724),
.B(n_1729),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1552),
.Y(n_1896)
);

A2O1A1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1713),
.A2(n_1709),
.B(n_1736),
.C(n_1743),
.Y(n_1897)
);

OA21x2_ASAP7_75t_L g1898 ( 
.A1(n_1689),
.A2(n_1714),
.B(n_1703),
.Y(n_1898)
);

OA22x2_ASAP7_75t_L g1899 ( 
.A1(n_1715),
.A2(n_1394),
.B1(n_1478),
.B2(n_1743),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1900)
);

AOI21x1_ASAP7_75t_SL g1901 ( 
.A1(n_1603),
.A2(n_1576),
.B(n_1544),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1709),
.A2(n_1736),
.B(n_1713),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1552),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1713),
.A2(n_1705),
.B1(n_1706),
.B2(n_1709),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1552),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1689),
.A2(n_1714),
.B(n_1703),
.Y(n_1909)
);

O2A1O1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1743),
.A2(n_1713),
.B(n_1736),
.C(n_1709),
.Y(n_1910)
);

OR2x6_ASAP7_75t_L g1911 ( 
.A(n_1794),
.B(n_1790),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1826),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1861),
.Y(n_1913)
);

AO21x2_ASAP7_75t_L g1914 ( 
.A1(n_1816),
.A2(n_1828),
.B(n_1807),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1845),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1846),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1776),
.B(n_1763),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1759),
.A2(n_1892),
.B1(n_1893),
.B2(n_1907),
.C(n_1890),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1803),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1774),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1767),
.B(n_1886),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1749),
.B(n_1878),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1829),
.B(n_1815),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1887),
.B(n_1894),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1750),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1834),
.B(n_1844),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1795),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1764),
.B(n_1779),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1767),
.B(n_1886),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1796),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1899),
.A2(n_1755),
.B1(n_1754),
.B2(n_1787),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1814),
.B(n_1800),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1855),
.A2(n_1871),
.B(n_1856),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1879),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1899),
.A2(n_1755),
.B1(n_1746),
.B2(n_1811),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1889),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1789),
.B(n_1791),
.Y(n_1937)
);

OA21x2_ASAP7_75t_L g1938 ( 
.A1(n_1873),
.A2(n_1825),
.B(n_1799),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1803),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1896),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1808),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1801),
.B(n_1802),
.Y(n_1942)
);

AO21x1_ASAP7_75t_SL g1943 ( 
.A1(n_1877),
.A2(n_1862),
.B(n_1854),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1759),
.B(n_1772),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1767),
.B(n_1886),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1904),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1903),
.B(n_1908),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1769),
.A2(n_1897),
.B(n_1891),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1797),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1764),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1772),
.A2(n_1910),
.B1(n_1885),
.B2(n_1902),
.C(n_1881),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1805),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1817),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1903),
.B(n_1745),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1823),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1884),
.B(n_1809),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1872),
.A2(n_1863),
.B(n_1860),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1803),
.B(n_1779),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1832),
.Y(n_1959)
);

OR2x6_ASAP7_75t_L g1960 ( 
.A(n_1773),
.B(n_1775),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1858),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1778),
.Y(n_1962)
);

AOI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1875),
.A2(n_1833),
.B(n_1784),
.Y(n_1963)
);

CKINVDCx8_ASAP7_75t_R g1964 ( 
.A(n_1830),
.Y(n_1964)
);

AO21x2_ASAP7_75t_L g1965 ( 
.A1(n_1855),
.A2(n_1825),
.B(n_1865),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1888),
.B(n_1850),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1812),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1888),
.B(n_1838),
.Y(n_1968)
);

BUFx2_ASAP7_75t_L g1969 ( 
.A(n_1819),
.Y(n_1969)
);

NOR2x1_ASAP7_75t_SL g1970 ( 
.A(n_1877),
.B(n_1786),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1842),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1819),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1883),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1891),
.A2(n_1897),
.B(n_1752),
.Y(n_1974)
);

AOI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1875),
.A2(n_1784),
.B(n_1782),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1786),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1883),
.Y(n_1977)
);

AOI221x1_ASAP7_75t_L g1978 ( 
.A1(n_1757),
.A2(n_1843),
.B1(n_1837),
.B2(n_1867),
.C(n_1866),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1857),
.Y(n_1979)
);

AOI221xp5_ASAP7_75t_L g1980 ( 
.A1(n_1747),
.A2(n_1785),
.B1(n_1806),
.B2(n_1781),
.C(n_1760),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1804),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1751),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1841),
.Y(n_1983)
);

BUFx12f_ASAP7_75t_L g1984 ( 
.A(n_1848),
.Y(n_1984)
);

AO21x2_ASAP7_75t_L g1985 ( 
.A1(n_1869),
.A2(n_1866),
.B(n_1849),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1831),
.B(n_1788),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1818),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1847),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1777),
.B(n_1748),
.Y(n_1989)
);

AO21x2_ASAP7_75t_L g1990 ( 
.A1(n_1869),
.A2(n_1853),
.B(n_1760),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1751),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1868),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1762),
.B(n_1874),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1874),
.B(n_1906),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1840),
.B(n_1810),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1868),
.B(n_1905),
.Y(n_1996)
);

AOI21xp33_ASAP7_75t_L g1997 ( 
.A1(n_1870),
.A2(n_1851),
.B(n_1864),
.Y(n_1997)
);

INVx4_ASAP7_75t_L g1998 ( 
.A(n_1765),
.Y(n_1998)
);

AND2x2_ASAP7_75t_SL g1999 ( 
.A(n_1756),
.B(n_1820),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1768),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1864),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1852),
.B(n_1859),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1932),
.B(n_1751),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1932),
.B(n_1909),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1926),
.B(n_1895),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1926),
.B(n_1909),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1950),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1961),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1961),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1941),
.B(n_1909),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1912),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1966),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1923),
.B(n_1898),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1923),
.B(n_1898),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1917),
.B(n_1898),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1912),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1928),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1913),
.B(n_1880),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1928),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1911),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1913),
.B(n_1761),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1921),
.B(n_1766),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1915),
.B(n_1916),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1916),
.B(n_1900),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1996),
.B(n_1784),
.Y(n_2025)
);

NAND2x1p5_ASAP7_75t_SL g2026 ( 
.A(n_1944),
.B(n_1770),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1954),
.B(n_1753),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1925),
.B(n_1821),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_2001),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1954),
.B(n_1753),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1911),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1921),
.B(n_1766),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1951),
.B(n_1793),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1919),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1992),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1956),
.B(n_1753),
.Y(n_2036)
);

O2A1O1Ixp5_ASAP7_75t_L g2037 ( 
.A1(n_1974),
.A2(n_1836),
.B(n_1839),
.C(n_1824),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1956),
.B(n_1758),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1949),
.B(n_1758),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1918),
.A2(n_1835),
.B1(n_1765),
.B2(n_1822),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1931),
.A2(n_1882),
.B1(n_1793),
.B2(n_1792),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1992),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1919),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1921),
.B(n_1783),
.Y(n_2044)
);

AOI21xp33_ASAP7_75t_L g2045 ( 
.A1(n_1948),
.A2(n_1901),
.B(n_1876),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1919),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1960),
.Y(n_2047)
);

AOI31xp33_ASAP7_75t_L g2048 ( 
.A1(n_1935),
.A2(n_1980),
.A3(n_2000),
.B(n_1994),
.Y(n_2048)
);

NOR2x1_ASAP7_75t_L g2049 ( 
.A(n_1960),
.B(n_1827),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1920),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1952),
.B(n_1835),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1952),
.B(n_1771),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1919),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1967),
.B(n_1780),
.Y(n_2054)
);

AOI33xp33_ASAP7_75t_L g2055 ( 
.A1(n_1958),
.A2(n_1798),
.A3(n_1813),
.B1(n_1927),
.B2(n_1934),
.B3(n_1946),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1942),
.B(n_1988),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1929),
.B(n_1945),
.Y(n_2057)
);

BUFx2_ASAP7_75t_L g2058 ( 
.A(n_1969),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1939),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1963),
.A2(n_1957),
.B(n_1975),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2018),
.B(n_1994),
.Y(n_2061)
);

AOI222xp33_ASAP7_75t_L g2062 ( 
.A1(n_2052),
.A2(n_1967),
.B1(n_1983),
.B2(n_1937),
.C1(n_1958),
.C2(n_1979),
.Y(n_2062)
);

NAND4xp25_ASAP7_75t_L g2063 ( 
.A(n_2045),
.B(n_1968),
.C(n_1993),
.D(n_1939),
.Y(n_2063)
);

NAND3xp33_ASAP7_75t_L g2064 ( 
.A(n_2045),
.B(n_1938),
.C(n_1968),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2050),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_2022),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2052),
.B(n_1981),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2050),
.Y(n_2068)
);

AOI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_2048),
.A2(n_1914),
.B1(n_1962),
.B2(n_1965),
.C(n_1953),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2035),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_2057),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_2039),
.Y(n_2072)
);

OAI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2048),
.A2(n_1960),
.B1(n_1999),
.B2(n_1964),
.Y(n_2073)
);

OAI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_2054),
.A2(n_1962),
.B1(n_1983),
.B2(n_1993),
.C(n_1997),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_2049),
.A2(n_1970),
.B(n_1914),
.Y(n_2075)
);

AOI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2006),
.A2(n_1914),
.B1(n_1965),
.B2(n_1953),
.C(n_1959),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2039),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2033),
.A2(n_1965),
.B1(n_1990),
.B2(n_1985),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_2057),
.Y(n_2079)
);

AOI221xp5_ASAP7_75t_L g2080 ( 
.A1(n_2006),
.A2(n_1955),
.B1(n_1959),
.B2(n_1924),
.C(n_1922),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2041),
.A2(n_1990),
.B1(n_1985),
.B2(n_1938),
.Y(n_2081)
);

AOI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2015),
.A2(n_1955),
.B1(n_1920),
.B2(n_1940),
.C(n_1946),
.Y(n_2082)
);

OAI211xp5_ASAP7_75t_SL g2083 ( 
.A1(n_2051),
.A2(n_1964),
.B(n_1939),
.C(n_1989),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_2007),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_2005),
.B(n_1995),
.Y(n_2085)
);

NOR4xp25_ASAP7_75t_SL g2086 ( 
.A(n_2020),
.B(n_1970),
.C(n_1977),
.D(n_1972),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2021),
.B(n_1943),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_2028),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2023),
.B(n_1936),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2035),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2042),
.Y(n_2091)
);

AOI21x1_ASAP7_75t_L g2092 ( 
.A1(n_2049),
.A2(n_1963),
.B(n_1975),
.Y(n_2092)
);

AOI221xp5_ASAP7_75t_L g2093 ( 
.A1(n_2015),
.A2(n_1930),
.B1(n_1936),
.B2(n_1934),
.C(n_1940),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_2057),
.Y(n_2094)
);

AOI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_2010),
.A2(n_1927),
.B1(n_1930),
.B2(n_1939),
.C(n_1933),
.Y(n_2095)
);

AOI221xp5_ASAP7_75t_L g2096 ( 
.A1(n_2010),
.A2(n_1933),
.B1(n_1979),
.B2(n_1991),
.C(n_1982),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2042),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2011),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_2025),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_SL g2100 ( 
.A1(n_2040),
.A2(n_1977),
.B(n_1973),
.C(n_1972),
.Y(n_2100)
);

AOI221xp5_ASAP7_75t_L g2101 ( 
.A1(n_2036),
.A2(n_2038),
.B1(n_2026),
.B2(n_2003),
.C(n_2004),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2005),
.A2(n_1938),
.B1(n_1943),
.B2(n_1933),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2011),
.Y(n_2103)
);

AO31x2_ASAP7_75t_L g2104 ( 
.A1(n_2029),
.A2(n_1978),
.A3(n_1971),
.B(n_1987),
.Y(n_2104)
);

BUFx3_ASAP7_75t_L g2105 ( 
.A(n_2022),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2016),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2023),
.B(n_2017),
.Y(n_2107)
);

NAND4xp25_ASAP7_75t_SL g2108 ( 
.A(n_2055),
.B(n_2051),
.C(n_2028),
.D(n_2021),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2012),
.B(n_1976),
.Y(n_2109)
);

OAI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2024),
.A2(n_1978),
.B1(n_1986),
.B2(n_1947),
.Y(n_2110)
);

NAND4xp25_ASAP7_75t_L g2111 ( 
.A(n_2040),
.B(n_2037),
.C(n_2025),
.D(n_2058),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_2022),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_2024),
.A2(n_2008),
.B1(n_2009),
.B2(n_2047),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2056),
.A2(n_1999),
.B1(n_1945),
.B2(n_1929),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2070),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2075),
.B(n_2057),
.Y(n_2116)
);

INVx4_ASAP7_75t_SL g2117 ( 
.A(n_2104),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2104),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2090),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_2067),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2084),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2110),
.B(n_2022),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2104),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2087),
.B(n_2013),
.Y(n_2124)
);

OA21x2_ASAP7_75t_L g2125 ( 
.A1(n_2078),
.A2(n_2060),
.B(n_2076),
.Y(n_2125)
);

INVx4_ASAP7_75t_SL g2126 ( 
.A(n_2104),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2080),
.B(n_2082),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2091),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2110),
.B(n_2032),
.Y(n_2129)
);

OA21x2_ASAP7_75t_L g2130 ( 
.A1(n_2069),
.A2(n_2060),
.B(n_2053),
.Y(n_2130)
);

OA21x2_ASAP7_75t_L g2131 ( 
.A1(n_2096),
.A2(n_2046),
.B(n_2059),
.Y(n_2131)
);

CKINVDCx16_ASAP7_75t_R g2132 ( 
.A(n_2073),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2097),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2065),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_2105),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_2092),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_2105),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_2071),
.B(n_2044),
.Y(n_2138)
);

OAI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_2064),
.A2(n_2038),
.B(n_2026),
.Y(n_2139)
);

BUFx12f_ASAP7_75t_L g2140 ( 
.A(n_2066),
.Y(n_2140)
);

INVx4_ASAP7_75t_SL g2141 ( 
.A(n_2079),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_2112),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2068),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2098),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2103),
.Y(n_2145)
);

OR2x6_ASAP7_75t_L g2146 ( 
.A(n_2114),
.B(n_2047),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_2079),
.B(n_2044),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_2094),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2106),
.Y(n_2149)
);

OAI21x1_ASAP7_75t_L g2150 ( 
.A1(n_2102),
.A2(n_2034),
.B(n_2043),
.Y(n_2150)
);

OA21x2_ASAP7_75t_L g2151 ( 
.A1(n_2095),
.A2(n_2053),
.B(n_2046),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2094),
.B(n_2044),
.Y(n_2152)
);

NOR2x1_ASAP7_75t_L g2153 ( 
.A(n_2111),
.B(n_1998),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2099),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2108),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2093),
.B(n_2019),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2127),
.B(n_2156),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2115),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_2156),
.B(n_2127),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2115),
.Y(n_2160)
);

OAI221xp5_ASAP7_75t_L g2161 ( 
.A1(n_2139),
.A2(n_2102),
.B1(n_2081),
.B2(n_2101),
.C(n_2062),
.Y(n_2161)
);

NOR3xp33_ASAP7_75t_SL g2162 ( 
.A(n_2139),
.B(n_2132),
.C(n_2083),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2120),
.B(n_2121),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2153),
.B(n_2061),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2153),
.B(n_2027),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2151),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2119),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2140),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2155),
.B(n_2088),
.Y(n_2169)
);

BUFx3_ASAP7_75t_L g2170 ( 
.A(n_2140),
.Y(n_2170)
);

INVx4_ASAP7_75t_L g2171 ( 
.A(n_2136),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2141),
.B(n_2027),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_L g2173 ( 
.A(n_2125),
.B(n_2081),
.C(n_2063),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2141),
.B(n_2030),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_2119),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_2140),
.B(n_1984),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2128),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2142),
.Y(n_2178)
);

AND2x2_ASAP7_75t_SL g2179 ( 
.A(n_2132),
.B(n_2031),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2142),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_2141),
.B(n_2099),
.Y(n_2181)
);

INVx2_ASAP7_75t_SL g2182 ( 
.A(n_2138),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2151),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2141),
.B(n_2030),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2141),
.B(n_2100),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2138),
.B(n_2109),
.Y(n_2186)
);

BUFx2_ASAP7_75t_L g2187 ( 
.A(n_2136),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2125),
.B(n_2085),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2138),
.B(n_2014),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2154),
.B(n_2089),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2138),
.B(n_2014),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2125),
.B(n_2072),
.Y(n_2192)
);

INVx2_ASAP7_75t_SL g2193 ( 
.A(n_2147),
.Y(n_2193)
);

NAND2xp33_ASAP7_75t_SL g2194 ( 
.A(n_2135),
.B(n_2086),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2125),
.B(n_2072),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2147),
.B(n_2152),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2151),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_2136),
.B(n_2151),
.C(n_2131),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2154),
.B(n_2107),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2147),
.B(n_2003),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2128),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2133),
.Y(n_2202)
);

INVx1_ASAP7_75t_SL g2203 ( 
.A(n_2136),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2133),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2130),
.B(n_2077),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2134),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2130),
.B(n_2077),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_2136),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2154),
.B(n_2017),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2180),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_2168),
.B(n_1984),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2190),
.B(n_2134),
.Y(n_2212)
);

OAI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2173),
.A2(n_2131),
.B(n_2130),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2185),
.B(n_2147),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2185),
.B(n_2152),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2166),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2167),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_2168),
.B(n_2135),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2175),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2158),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2190),
.B(n_2143),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2158),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2180),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2166),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2196),
.B(n_2152),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2157),
.B(n_2143),
.Y(n_2226)
);

NOR3xp33_ASAP7_75t_L g2227 ( 
.A(n_2157),
.B(n_2129),
.C(n_2122),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2196),
.B(n_2152),
.Y(n_2228)
);

OR2x2_ASAP7_75t_L g2229 ( 
.A(n_2199),
.B(n_2144),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2164),
.B(n_2137),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2173),
.A2(n_2131),
.B1(n_2130),
.B2(n_2126),
.Y(n_2231)
);

OAI22xp33_ASAP7_75t_SL g2232 ( 
.A1(n_2159),
.A2(n_2146),
.B1(n_2074),
.B2(n_2118),
.Y(n_2232)
);

NAND2x1p5_ASAP7_75t_L g2233 ( 
.A(n_2179),
.B(n_2170),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2160),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_2170),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2164),
.B(n_2137),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2186),
.B(n_2124),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2199),
.B(n_2144),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2163),
.B(n_2145),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2160),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2159),
.B(n_2145),
.Y(n_2241)
);

AOI32xp33_ASAP7_75t_L g2242 ( 
.A1(n_2161),
.A2(n_2150),
.A3(n_2116),
.B1(n_2113),
.B2(n_2131),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2186),
.B(n_2124),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2209),
.B(n_2149),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2182),
.B(n_2193),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_2181),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2182),
.B(n_2148),
.Y(n_2247)
);

AOI21xp33_ASAP7_75t_L g2248 ( 
.A1(n_2198),
.A2(n_2136),
.B(n_2123),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2209),
.B(n_2149),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2177),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2241),
.B(n_2227),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2241),
.B(n_2178),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2235),
.B(n_2176),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2213),
.A2(n_2179),
.B1(n_2231),
.B2(n_2198),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2210),
.Y(n_2255)
);

INVxp67_ASAP7_75t_L g2256 ( 
.A(n_2223),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2226),
.B(n_2217),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2237),
.B(n_2170),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2219),
.B(n_2177),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_2246),
.B(n_2193),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_2233),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_2233),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2218),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2233),
.Y(n_2264)
);

INVx1_ASAP7_75t_SL g2265 ( 
.A(n_2235),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2216),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2237),
.B(n_2162),
.Y(n_2267)
);

INVx4_ASAP7_75t_L g2268 ( 
.A(n_2246),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2245),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2211),
.Y(n_2270)
);

HB1xp67_ASAP7_75t_L g2271 ( 
.A(n_2245),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2216),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2224),
.Y(n_2273)
);

NOR2xp67_ASAP7_75t_L g2274 ( 
.A(n_2246),
.B(n_2171),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_2224),
.Y(n_2275)
);

INVxp67_ASAP7_75t_L g2276 ( 
.A(n_2239),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_2248),
.A2(n_2179),
.B1(n_2183),
.B2(n_2166),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2220),
.B(n_2201),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2243),
.B(n_2165),
.Y(n_2279)
);

CKINVDCx16_ASAP7_75t_R g2280 ( 
.A(n_2230),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_SL g2281 ( 
.A1(n_2280),
.A2(n_2169),
.B1(n_2171),
.B2(n_2208),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2280),
.B(n_2230),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2255),
.Y(n_2283)
);

INVx2_ASAP7_75t_SL g2284 ( 
.A(n_2260),
.Y(n_2284)
);

A2O1A1Ixp33_ASAP7_75t_L g2285 ( 
.A1(n_2254),
.A2(n_2242),
.B(n_2183),
.C(n_2197),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2275),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2258),
.B(n_2236),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2265),
.B(n_2239),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2265),
.B(n_2243),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2251),
.A2(n_2232),
.B(n_2195),
.Y(n_2290)
);

O2A1O1Ixp33_ASAP7_75t_L g2291 ( 
.A1(n_2251),
.A2(n_2192),
.B(n_2207),
.C(n_2205),
.Y(n_2291)
);

A2O1A1Ixp33_ASAP7_75t_L g2292 ( 
.A1(n_2277),
.A2(n_2183),
.B(n_2197),
.C(n_2194),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2269),
.B(n_2236),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2275),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2275),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2272),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2258),
.B(n_2214),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2272),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2267),
.A2(n_2197),
.B1(n_2188),
.B2(n_2126),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2256),
.A2(n_2208),
.B(n_2187),
.Y(n_2300)
);

AOI321xp33_ASAP7_75t_SL g2301 ( 
.A1(n_2264),
.A2(n_2203),
.A3(n_2214),
.B1(n_2215),
.B2(n_2225),
.C(n_2228),
.Y(n_2301)
);

INVx1_ASAP7_75t_SL g2302 ( 
.A(n_2271),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2261),
.B(n_2171),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_2267),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2290),
.A2(n_2272),
.B1(n_2266),
.B2(n_2273),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2296),
.Y(n_2306)
);

AND2x4_ASAP7_75t_SL g2307 ( 
.A(n_2282),
.B(n_2253),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_2282),
.Y(n_2308)
);

INVxp67_ASAP7_75t_L g2309 ( 
.A(n_2284),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2297),
.B(n_2256),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2285),
.A2(n_2263),
.B1(n_2270),
.B2(n_2276),
.Y(n_2311)
);

INVx1_ASAP7_75t_SL g2312 ( 
.A(n_2287),
.Y(n_2312)
);

NAND2x1_ASAP7_75t_L g2313 ( 
.A(n_2297),
.B(n_2261),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2298),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2287),
.B(n_2264),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2304),
.B(n_2286),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2284),
.B(n_2279),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2286),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2295),
.A2(n_2273),
.B1(n_2266),
.B2(n_2262),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2295),
.B(n_2261),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2305),
.A2(n_2117),
.B1(n_2126),
.B2(n_2118),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2308),
.A2(n_2285),
.B1(n_2292),
.B2(n_2289),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2307),
.B(n_2261),
.Y(n_2323)
);

AOI222xp33_ASAP7_75t_L g2324 ( 
.A1(n_2305),
.A2(n_2292),
.B1(n_2294),
.B2(n_2288),
.C1(n_2126),
.C2(n_2117),
.Y(n_2324)
);

AOI221x1_ASAP7_75t_L g2325 ( 
.A1(n_2318),
.A2(n_2300),
.B1(n_2283),
.B2(n_2281),
.C(n_2268),
.Y(n_2325)
);

NAND3xp33_ASAP7_75t_L g2326 ( 
.A(n_2311),
.B(n_2291),
.C(n_2268),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2319),
.A2(n_2299),
.B1(n_2257),
.B2(n_2302),
.C(n_2262),
.Y(n_2327)
);

OAI21xp5_ASAP7_75t_SL g2328 ( 
.A1(n_2312),
.A2(n_2293),
.B(n_2252),
.Y(n_2328)
);

OAI221xp5_ASAP7_75t_L g2329 ( 
.A1(n_2319),
.A2(n_2257),
.B1(n_2203),
.B2(n_2274),
.C(n_2171),
.Y(n_2329)
);

O2A1O1Ixp33_ASAP7_75t_L g2330 ( 
.A1(n_2316),
.A2(n_2303),
.B(n_2259),
.C(n_2252),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2317),
.B(n_2279),
.Y(n_2331)
);

OAI321xp33_ASAP7_75t_L g2332 ( 
.A1(n_2315),
.A2(n_2301),
.A3(n_2303),
.B1(n_2259),
.B2(n_2187),
.C(n_2215),
.Y(n_2332)
);

AOI32xp33_ASAP7_75t_L g2333 ( 
.A1(n_2306),
.A2(n_2260),
.A3(n_2165),
.B1(n_2268),
.B2(n_2278),
.Y(n_2333)
);

AO221x1_ASAP7_75t_L g2334 ( 
.A1(n_2322),
.A2(n_2309),
.B1(n_2314),
.B2(n_2250),
.C(n_2240),
.Y(n_2334)
);

AOI322xp5_ASAP7_75t_L g2335 ( 
.A1(n_2327),
.A2(n_2310),
.A3(n_2320),
.B1(n_2313),
.B2(n_2278),
.C1(n_2123),
.C2(n_2118),
.Y(n_2335)
);

AOI21xp33_ASAP7_75t_SL g2336 ( 
.A1(n_2326),
.A2(n_2320),
.B(n_2260),
.Y(n_2336)
);

INVx1_ASAP7_75t_SL g2337 ( 
.A(n_2331),
.Y(n_2337)
);

O2A1O1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_2332),
.A2(n_2250),
.B(n_2274),
.C(n_2222),
.Y(n_2338)
);

OAI21xp33_ASAP7_75t_L g2339 ( 
.A1(n_2323),
.A2(n_2260),
.B(n_2234),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2328),
.B(n_2268),
.Y(n_2340)
);

O2A1O1Ixp33_ASAP7_75t_L g2341 ( 
.A1(n_2324),
.A2(n_2229),
.B(n_2238),
.C(n_2212),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2337),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2340),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2334),
.A2(n_2325),
.B(n_2330),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2341),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2338),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2339),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2336),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2335),
.Y(n_2349)
);

AND2x2_ASAP7_75t_SL g2350 ( 
.A(n_2342),
.B(n_2321),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_R g2351 ( 
.A(n_2347),
.B(n_2348),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2343),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2345),
.Y(n_2353)
);

OAI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2349),
.A2(n_2333),
.B1(n_2329),
.B2(n_2229),
.C(n_2238),
.Y(n_2354)
);

OAI221xp5_ASAP7_75t_L g2355 ( 
.A1(n_2344),
.A2(n_2212),
.B1(n_2221),
.B2(n_2244),
.C(n_2249),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2352),
.B(n_2344),
.Y(n_2356)
);

AOI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2353),
.A2(n_2346),
.B1(n_2228),
.B2(n_2225),
.Y(n_2357)
);

NOR2x1_ASAP7_75t_L g2358 ( 
.A(n_2355),
.B(n_2244),
.Y(n_2358)
);

NAND2x1_ASAP7_75t_L g2359 ( 
.A(n_2351),
.B(n_2247),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2358),
.B(n_2350),
.Y(n_2360)
);

BUFx2_ASAP7_75t_L g2361 ( 
.A(n_2359),
.Y(n_2361)
);

AOI222xp33_ASAP7_75t_L g2362 ( 
.A1(n_2360),
.A2(n_2356),
.B1(n_2354),
.B2(n_2126),
.C1(n_2117),
.C2(n_2357),
.Y(n_2362)
);

AOI31xp33_ASAP7_75t_L g2363 ( 
.A1(n_2360),
.A2(n_2002),
.A3(n_2247),
.B(n_2249),
.Y(n_2363)
);

OAI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2362),
.A2(n_2361),
.B(n_2221),
.Y(n_2364)
);

OR4x1_ASAP7_75t_L g2365 ( 
.A(n_2363),
.B(n_2206),
.C(n_2204),
.D(n_2201),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2365),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2364),
.B(n_2117),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2367),
.A2(n_2123),
.B1(n_2117),
.B2(n_2181),
.Y(n_2368)
);

INVx1_ASAP7_75t_SL g2369 ( 
.A(n_2366),
.Y(n_2369)
);

OAI22xp33_ASAP7_75t_L g2370 ( 
.A1(n_2369),
.A2(n_2206),
.B1(n_2204),
.B2(n_2202),
.Y(n_2370)
);

NAND4xp75_ASAP7_75t_L g2371 ( 
.A(n_2370),
.B(n_2368),
.C(n_2184),
.D(n_2172),
.Y(n_2371)
);

OAI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2371),
.A2(n_2181),
.B(n_2202),
.Y(n_2372)
);

NAND3xp33_ASAP7_75t_L g2373 ( 
.A(n_2372),
.B(n_2181),
.C(n_2172),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2373),
.A2(n_2184),
.B1(n_2174),
.B2(n_2189),
.Y(n_2374)
);

AOI211xp5_ASAP7_75t_L g2375 ( 
.A1(n_2374),
.A2(n_2174),
.B(n_2191),
.C(n_2200),
.Y(n_2375)
);


endmodule