module fake_jpeg_441_n_473 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_55),
.B(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_65),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_57),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_61),
.B(n_69),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_63),
.Y(n_160)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_68),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_10),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_70),
.B(n_79),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_11),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_81),
.B(n_94),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_19),
.B(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_88),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_35),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_93),
.B(n_106),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_95),
.B(n_99),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_0),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_28),
.Y(n_102)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_23),
.B(n_0),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_27),
.B(n_0),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_112),
.Y(n_136)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_27),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_51),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_2),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_31),
.B1(n_45),
.B2(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_138),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_54),
.B1(n_45),
.B2(n_34),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_53),
.Y(n_120)
);

NAND2x1p5_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_146),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_53),
.B1(n_54),
.B2(n_45),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_92),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_76),
.A2(n_86),
.B1(n_78),
.B2(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_134),
.A2(n_170),
.B1(n_142),
.B2(n_147),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_54),
.B1(n_34),
.B2(n_42),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_90),
.B(n_53),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_140),
.Y(n_199)
);

NAND2x1p5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_148),
.B(n_131),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_42),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_68),
.Y(n_201)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_57),
.Y(n_154)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_85),
.A2(n_50),
.B1(n_51),
.B2(n_46),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_122),
.B1(n_187),
.B2(n_138),
.Y(n_216)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_101),
.A2(n_25),
.B1(n_46),
.B2(n_41),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_182),
.B1(n_187),
.B2(n_110),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_98),
.A2(n_25),
.B1(n_41),
.B2(n_39),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_62),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_84),
.A2(n_37),
.B1(n_39),
.B2(n_4),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_189),
.B(n_196),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_191),
.Y(n_289)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_108),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_195),
.B(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_77),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_197),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_200),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_201),
.A2(n_210),
.B(n_214),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_2),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_2),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_211),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_3),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_204),
.B(n_209),
.Y(n_279)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_206),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_5),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_136),
.A2(n_67),
.B1(n_75),
.B2(n_113),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_5),
.Y(n_211)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_5),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_120),
.A2(n_83),
.B(n_37),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_215),
.A2(n_246),
.B(n_244),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_216),
.A2(n_247),
.B1(n_197),
.B2(n_198),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_117),
.A2(n_37),
.B1(n_39),
.B2(n_140),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_249),
.B1(n_215),
.B2(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_37),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_226),
.Y(n_265)
);

OR2x2_ASAP7_75t_SL g220 ( 
.A(n_136),
.B(n_39),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_170),
.C(n_201),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_158),
.A2(n_124),
.B(n_121),
.C(n_159),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_125),
.B(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_127),
.A2(n_141),
.B1(n_145),
.B2(n_118),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_173),
.A2(n_159),
.B1(n_139),
.B2(n_133),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_225),
.A2(n_238),
.B1(n_212),
.B2(n_200),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_164),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_153),
.Y(n_227)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_130),
.Y(n_231)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_232),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_129),
.B(n_135),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_139),
.Y(n_234)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_134),
.A2(n_174),
.B1(n_188),
.B2(n_144),
.Y(n_238)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_119),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_150),
.B(n_155),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_179),
.Y(n_243)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_157),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_150),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_155),
.A2(n_157),
.B(n_168),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_126),
.B(n_137),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_254),
.B(n_281),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_255),
.A2(n_264),
.B1(n_274),
.B2(n_277),
.Y(n_318)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_194),
.B1(n_249),
.B2(n_199),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_195),
.A2(n_202),
.B1(n_194),
.B2(n_218),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_190),
.B1(n_223),
.B2(n_236),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_194),
.A2(n_201),
.B(n_220),
.C(n_206),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_250),
.B(n_252),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_224),
.A2(n_241),
.B1(n_246),
.B2(n_226),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_203),
.B(n_221),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_287),
.C(n_290),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_192),
.B1(n_245),
.B2(n_224),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_211),
.B(n_242),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_213),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_213),
.B1(n_242),
.B2(n_237),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_239),
.B1(n_240),
.B2(n_207),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_282),
.B1(n_280),
.B2(n_289),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_297),
.A2(n_312),
.B1(n_325),
.B2(n_314),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_255),
.A2(n_207),
.B1(n_205),
.B2(n_219),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_298),
.A2(n_295),
.B1(n_267),
.B2(n_260),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_219),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_312),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_237),
.B1(n_190),
.B2(n_229),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_301),
.A2(n_306),
.B1(n_307),
.B2(n_315),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_302),
.B(n_321),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_303),
.B(n_304),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_248),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_264),
.A2(n_250),
.B1(n_261),
.B2(n_251),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_323),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_250),
.A2(n_252),
.B1(n_258),
.B2(n_265),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_275),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_316),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_285),
.B(n_271),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_317),
.A2(n_294),
.B(n_273),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_320),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_257),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_266),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_258),
.A2(n_277),
.B1(n_254),
.B2(n_284),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_324),
.A2(n_327),
.B1(n_331),
.B2(n_302),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_290),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_329),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_258),
.A2(n_279),
.B1(n_270),
.B2(n_268),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_253),
.B(n_268),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_286),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_330),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_269),
.A2(n_256),
.B1(n_294),
.B2(n_288),
.Y(n_331)
);

OA21x2_ASAP7_75t_SL g380 ( 
.A1(n_332),
.A2(n_348),
.B(n_297),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_260),
.C(n_267),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_342),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_356),
.B1(n_331),
.B2(n_306),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_291),
.C(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_291),
.C(n_309),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_299),
.C(n_326),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_351),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_296),
.A2(n_318),
.B1(n_325),
.B2(n_298),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_350),
.A2(n_313),
.B(n_311),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_308),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_353),
.A2(n_324),
.B1(n_315),
.B2(n_317),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_337),
.A2(n_325),
.B(n_310),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_376),
.B(n_335),
.Y(n_394)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_321),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_367),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_379),
.B1(n_332),
.B2(n_336),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_346),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_319),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_369),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_343),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_370),
.A2(n_357),
.B1(n_340),
.B2(n_353),
.Y(n_384)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_375),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_345),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_372),
.B(n_377),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_358),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_374),
.Y(n_403)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_337),
.A2(n_352),
.B(n_344),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_378),
.B(n_382),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_350),
.A2(n_305),
.B1(n_328),
.B2(n_320),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_380),
.B(n_348),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_381),
.A2(n_335),
.B(n_359),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_322),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_385),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_397),
.B1(n_379),
.B2(n_381),
.Y(n_409)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_344),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_388),
.A2(n_400),
.B1(n_361),
.B2(n_381),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_377),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_369),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_342),
.C(n_349),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_392),
.C(n_399),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_357),
.C(n_359),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_394),
.B(n_361),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_370),
.A2(n_333),
.B1(n_341),
.B2(n_364),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_333),
.C(n_341),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_360),
.B1(n_376),
.B2(n_365),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_374),
.B(n_368),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_407),
.B(n_417),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_373),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_411),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_410),
.A2(n_394),
.B(n_393),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_392),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_389),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_415),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_416),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_367),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_362),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_418),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_380),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_419),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_379),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_420),
.B(n_414),
.C(n_388),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_421),
.A2(n_400),
.B(n_415),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_384),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_425),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_403),
.Y(n_431)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_426),
.A2(n_412),
.B(n_414),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_434),
.A2(n_427),
.B1(n_424),
.B2(n_431),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_421),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_432),
.B(n_411),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_436),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_420),
.C(n_408),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_443),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_396),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_439),
.B(n_441),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_428),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_440),
.A2(n_430),
.B(n_425),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_397),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_433),
.C(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_447),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_438),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_449),
.B(n_452),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_437),
.B(n_430),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_440),
.C(n_442),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_433),
.C(n_429),
.Y(n_452)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_455),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_457),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_444),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_409),
.C(n_398),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_459),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_398),
.C(n_402),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_452),
.Y(n_461)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_461),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_450),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_375),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_460),
.A2(n_449),
.B(n_446),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_465),
.A2(n_463),
.B1(n_366),
.B2(n_378),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_464),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_468),
.B(n_469),
.Y(n_470)
);

OAI321xp33_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_371),
.A3(n_395),
.B1(n_463),
.B2(n_466),
.C(n_460),
.Y(n_471)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_471),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_395),
.Y(n_473)
);


endmodule