module fake_jpeg_17087_n_167 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx2_ASAP7_75t_SL g75 ( 
.A(n_72),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_50),
.B1(n_41),
.B2(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_45),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_61),
.B(n_43),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_63),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_47),
.B1(n_62),
.B2(n_55),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_59),
.B1(n_56),
.B2(n_49),
.Y(n_116)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_89),
.Y(n_98)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_58),
.Y(n_102)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_99),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_102),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_59),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_112),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_111),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_64),
.B1(n_60),
.B2(n_57),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_116),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_0),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_0),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_4),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_107),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_135),
.B(n_133),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_119),
.B1(n_101),
.B2(n_118),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_145),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_95),
.B1(n_117),
.B2(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_96),
.B1(n_108),
.B2(n_115),
.Y(n_149)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_140),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_141),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_153),
.B1(n_149),
.B2(n_120),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_146),
.B1(n_149),
.B2(n_124),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_128),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_98),
.C(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_98),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_94),
.C(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_7),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_14),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_20),
.B(n_23),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_24),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_26),
.C(n_27),
.Y(n_167)
);


endmodule