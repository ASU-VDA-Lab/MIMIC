module fake_jpeg_3084_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

AOI21xp33_ASAP7_75t_L g11 ( 
.A1(n_5),
.A2(n_2),
.B(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_21),
.B1(n_10),
.B2(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_6),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_15),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_23),
.B1(n_24),
.B2(n_20),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_32),
.B1(n_13),
.B2(n_17),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.C(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_22),
.B(n_19),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_29),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_13),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_30),
.C(n_26),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.C(n_40),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_33),
.C(n_9),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_0),
.C(n_5),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_38),
.B1(n_13),
.B2(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_51),
.B1(n_48),
.B2(n_47),
.Y(n_54)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_51),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_50),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_55),
.B(n_50),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_52),
.B(n_49),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_56),
.Y(n_59)
);


endmodule