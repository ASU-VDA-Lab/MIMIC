module fake_jpeg_31916_n_91 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx10_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_38),
.B1(n_32),
.B2(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_43),
.B1(n_33),
.B2(n_17),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_16),
.B1(n_28),
.B2(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_33),
.B(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_29),
.B1(n_13),
.B2(n_14),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_4),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_5),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_70),
.B1(n_15),
.B2(n_18),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_11),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_72),
.C(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_21),
.C(n_22),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_73),
.B(n_69),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_78),
.B1(n_76),
.B2(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_80),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_83),
.A3(n_64),
.B1(n_85),
.B2(n_63),
.C1(n_25),
.C2(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);


endmodule