module real_aes_5183_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g249 ( .A(n_0), .B(n_250), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_1), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_2), .A2(n_76), .B1(n_153), .B2(n_156), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_SL g334 ( .A1(n_3), .A2(n_265), .B(n_335), .C(n_336), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_4), .A2(n_61), .B1(n_254), .B2(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_5), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_6), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_7), .A2(n_53), .B1(n_239), .B2(n_257), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_8), .Y(n_364) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
INVxp67_ASAP7_75t_L g144 ( .A(n_9), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_9), .B(n_55), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_10), .A2(n_56), .B1(n_132), .B2(n_135), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_11), .A2(n_45), .B1(n_254), .B2(n_271), .Y(n_324) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_12), .A2(n_52), .B(n_227), .Y(n_226) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_12), .A2(n_52), .B(n_227), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_13), .B(n_93), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_14), .Y(n_286) );
BUFx3_ASAP7_75t_L g200 ( .A(n_15), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_16), .A2(n_258), .B(n_340), .C(n_341), .Y(n_339) );
OAI22xp33_ASAP7_75t_SL g253 ( .A1(n_17), .A2(n_30), .B1(n_233), .B2(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_18), .A2(n_23), .B1(n_233), .B2(n_235), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_19), .A2(n_68), .B1(n_178), .B2(n_180), .Y(n_177) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
O2A1O1Ixp5_ASAP7_75t_L g304 ( .A1(n_21), .A2(n_265), .B(n_305), .C(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g94 ( .A(n_22), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_22), .B(n_54), .Y(n_141) );
AOI221xp5_ASAP7_75t_L g159 ( .A1(n_24), .A2(n_41), .B1(n_160), .B2(n_163), .C(n_166), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_25), .A2(n_34), .B1(n_146), .B2(n_148), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_26), .B(n_243), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_27), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g87 ( .A1(n_28), .A2(n_42), .B1(n_88), .B2(n_111), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_29), .Y(n_82) );
INVx1_ASAP7_75t_L g227 ( .A(n_31), .Y(n_227) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_32), .Y(n_211) );
AND2x4_ASAP7_75t_L g228 ( .A(n_32), .B(n_209), .Y(n_228) );
AND2x4_ASAP7_75t_L g260 ( .A(n_32), .B(n_209), .Y(n_260) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_33), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_35), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_36), .A2(n_265), .B(n_290), .C(n_292), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_37), .Y(n_313) );
INVx2_ASAP7_75t_L g369 ( .A(n_38), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_39), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_40), .A2(n_69), .B1(n_116), .B2(n_121), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_43), .B(n_274), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_44), .A2(n_59), .B1(n_238), .B2(n_240), .Y(n_237) );
OA22x2_ASAP7_75t_L g98 ( .A1(n_46), .A2(n_55), .B1(n_93), .B2(n_97), .Y(n_98) );
INVx1_ASAP7_75t_L g128 ( .A(n_46), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_47), .Y(n_193) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_48), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_49), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g608 ( .A(n_50), .B(n_84), .Y(n_608) );
NAND2xp33_ASAP7_75t_R g328 ( .A(n_51), .B(n_226), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_51), .A2(n_75), .B1(n_243), .B2(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_54), .B(n_126), .Y(n_176) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_54), .Y(n_203) );
OAI21xp33_ASAP7_75t_L g129 ( .A1(n_55), .A2(n_60), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_57), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_58), .Y(n_365) );
INVx1_ASAP7_75t_L g96 ( .A(n_60), .Y(n_96) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_60), .B(n_72), .Y(n_174) );
INVx1_ASAP7_75t_L g167 ( .A(n_62), .Y(n_167) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_63), .Y(n_234) );
INVx1_ASAP7_75t_L g236 ( .A(n_63), .Y(n_236) );
BUFx5_ASAP7_75t_L g254 ( .A(n_63), .Y(n_254) );
INVx2_ASAP7_75t_L g345 ( .A(n_64), .Y(n_345) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_65), .Y(n_189) );
INVx2_ASAP7_75t_L g295 ( .A(n_66), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_67), .Y(n_342) );
INVx2_ASAP7_75t_SL g209 ( .A(n_70), .Y(n_209) );
INVx1_ASAP7_75t_L g311 ( .A(n_71), .Y(n_311) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_71), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_72), .B(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g317 ( .A(n_73), .Y(n_317) );
OAI21xp33_ASAP7_75t_SL g284 ( .A1(n_74), .A2(n_254), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_75), .B(n_243), .Y(n_359) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_75), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_195), .B1(n_212), .B2(n_595), .C(n_601), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_182), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_83), .B2(n_84), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_82), .B(n_337), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_83), .A2(n_84), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NOR2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_151), .Y(n_85) );
NAND4xp25_ASAP7_75t_L g86 ( .A(n_87), .B(n_115), .C(n_131), .D(n_145), .Y(n_86) );
BUFx4f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_99), .Y(n_89) );
AND2x4_ASAP7_75t_L g112 ( .A(n_90), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g132 ( .A(n_90), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g165 ( .A(n_90), .B(n_149), .Y(n_165) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_98), .Y(n_90) );
INVx1_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g91 ( .A(n_92), .B(n_95), .Y(n_91) );
NAND2xp33_ASAP7_75t_L g92 ( .A(n_93), .B(n_94), .Y(n_92) );
INVx2_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
INVx3_ASAP7_75t_L g102 ( .A(n_93), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g109 ( .A(n_93), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_94), .B(n_128), .Y(n_127) );
INVxp67_ASAP7_75t_L g204 ( .A(n_94), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_96), .A2(n_130), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g120 ( .A(n_98), .Y(n_120) );
AND2x2_ASAP7_75t_L g142 ( .A(n_98), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g147 ( .A(n_98), .B(n_119), .Y(n_147) );
AND2x4_ASAP7_75t_L g117 ( .A(n_99), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g123 ( .A(n_99), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_104), .Y(n_99) );
OR2x2_ASAP7_75t_L g114 ( .A(n_100), .B(n_105), .Y(n_114) );
AND2x4_ASAP7_75t_L g133 ( .A(n_100), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g138 ( .A(n_100), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_103), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_102), .B(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
NAND3xp33_ASAP7_75t_L g175 ( .A(n_103), .B(n_125), .C(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
BUFx12f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g154 ( .A(n_118), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g179 ( .A(n_118), .B(n_149), .Y(n_179) );
AND2x4_ASAP7_75t_L g181 ( .A(n_118), .B(n_133), .Y(n_181) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx2_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx8_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g148 ( .A(n_124), .B(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g158 ( .A(n_124), .B(n_155), .Y(n_158) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_128), .Y(n_205) );
AND2x4_ASAP7_75t_L g146 ( .A(n_133), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g149 ( .A(n_134), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx1_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_141), .Y(n_201) );
AND2x4_ASAP7_75t_L g162 ( .A(n_147), .B(n_149), .Y(n_162) );
NAND3xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_159), .C(n_177), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx6_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx12f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B1(n_193), .B2(n_194), .Y(n_182) );
CKINVDCx14_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B1(n_191), .B2(n_192), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_185), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_186), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_187), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_193), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_206), .Y(n_197) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g606 ( .A(n_199), .B(n_206), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .C(n_205), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_210), .Y(n_206) );
OR2x2_ASAP7_75t_L g610 ( .A(n_207), .B(n_211), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_207), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_207), .B(n_210), .Y(n_614) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_465), .Y(n_214) );
AND4x1_ASAP7_75t_L g215 ( .A(n_216), .B(n_413), .C(n_433), .D(n_445), .Y(n_215) );
AOI311xp33_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_296), .A3(n_329), .B(n_346), .C(n_383), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_276), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_246), .Y(n_219) );
INVx3_ASAP7_75t_L g382 ( .A(n_220), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_220), .B(n_406), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_220), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g535 ( .A(n_220), .B(n_519), .Y(n_535) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g424 ( .A(n_221), .B(n_350), .Y(n_424) );
INVx1_ASAP7_75t_L g487 ( .A(n_221), .Y(n_487) );
AND2x2_ASAP7_75t_L g529 ( .A(n_221), .B(n_261), .Y(n_529) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g505 ( .A(n_222), .Y(n_505) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_242), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_224), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
INVx1_ASAP7_75t_L g318 ( .A(n_226), .Y(n_318) );
INVx2_ASAP7_75t_L g378 ( .A(n_226), .Y(n_378) );
AND2x2_ASAP7_75t_L g281 ( .A(n_228), .B(n_282), .Y(n_281) );
INVx4_ASAP7_75t_L g314 ( .A(n_228), .Y(n_314) );
INVx1_ASAP7_75t_L g400 ( .A(n_229), .Y(n_400) );
OA22x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_232), .B1(n_237), .B2(n_241), .Y(n_229) );
INVx4_ASAP7_75t_L g599 ( .A(n_230), .Y(n_599) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g241 ( .A(n_231), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_231), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g258 ( .A(n_231), .Y(n_258) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_231), .Y(n_265) );
INVx4_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_231), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g240 ( .A(n_233), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g266 ( .A1(n_233), .A2(n_254), .B1(n_267), .B2(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_233), .A2(n_254), .B1(n_364), .B2(n_365), .Y(n_363) );
INVx6_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g257 ( .A(n_234), .Y(n_257) );
INVx2_ASAP7_75t_L g271 ( .A(n_234), .Y(n_271) );
INVx3_ASAP7_75t_L g291 ( .A(n_234), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_235), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_235), .B(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_235), .A2(n_271), .B1(n_368), .B2(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g239 ( .A(n_236), .Y(n_239) );
INVx1_ASAP7_75t_L g335 ( .A(n_238), .Y(n_335) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g403 ( .A(n_242), .Y(n_403) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g250 ( .A(n_244), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_244), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g344 ( .A(n_244), .B(n_345), .Y(n_344) );
INVx4_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g275 ( .A(n_245), .Y(n_275) );
BUFx3_ASAP7_75t_L g402 ( .A(n_245), .Y(n_402) );
AND2x2_ASAP7_75t_L g516 ( .A(n_246), .B(n_382), .Y(n_516) );
INVx1_ASAP7_75t_SL g540 ( .A(n_246), .Y(n_540) );
AND2x2_ASAP7_75t_L g553 ( .A(n_246), .B(n_504), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_246), .B(n_348), .Y(n_554) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_261), .Y(n_246) );
AND2x2_ASAP7_75t_L g437 ( .A(n_247), .B(n_279), .Y(n_437) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
NAND2xp33_ASAP7_75t_R g396 ( .A(n_248), .B(n_279), .Y(n_396) );
AND2x2_ASAP7_75t_L g406 ( .A(n_248), .B(n_261), .Y(n_406) );
INVx1_ASAP7_75t_L g477 ( .A(n_248), .Y(n_477) );
AND2x2_ASAP7_75t_L g519 ( .A(n_248), .B(n_279), .Y(n_519) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_248), .Y(n_546) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
INVx2_ASAP7_75t_L g263 ( .A(n_250), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g343 ( .A(n_250), .B(n_314), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_254), .A2(n_270), .B1(n_271), .B2(n_272), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_254), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_254), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_254), .B(n_313), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_258), .B(n_259), .Y(n_255) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_258), .A2(n_260), .B1(n_265), .B2(n_266), .C(n_269), .Y(n_264) );
INVx1_ASAP7_75t_L g327 ( .A(n_260), .Y(n_327) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_260), .Y(n_390) );
OR2x2_ASAP7_75t_L g398 ( .A(n_261), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g486 ( .A(n_261), .B(n_487), .Y(n_486) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_273), .Y(n_261) );
OA21x2_ASAP7_75t_L g352 ( .A1(n_262), .A2(n_264), .B(n_273), .Y(n_352) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g392 ( .A(n_263), .B(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_265), .A2(n_288), .B1(n_324), .B2(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g370 ( .A(n_265), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_265), .A2(n_288), .B1(n_363), .B2(n_367), .Y(n_391) );
INVx1_ASAP7_75t_L g340 ( .A(n_271), .Y(n_340) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_274), .B(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_275), .B(n_295), .Y(n_294) );
BUFx3_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
AND2x2_ASAP7_75t_L g549 ( .A(n_276), .B(n_530), .Y(n_549) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g558 ( .A(n_277), .B(n_496), .Y(n_558) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g405 ( .A(n_278), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g499 ( .A(n_278), .Y(n_499) );
AND2x2_ASAP7_75t_L g504 ( .A(n_278), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx2_ASAP7_75t_L g348 ( .A(n_279), .Y(n_348) );
INVx2_ASAP7_75t_L g419 ( .A(n_279), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_279), .B(n_352), .Y(n_422) );
INVx1_ASAP7_75t_L g449 ( .A(n_279), .Y(n_449) );
OR2x2_ASAP7_75t_L g456 ( .A(n_279), .B(n_350), .Y(n_456) );
AND2x2_ASAP7_75t_L g490 ( .A(n_279), .B(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B(n_294), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_289), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_287), .A2(n_314), .B1(n_362), .B2(n_366), .C(n_370), .Y(n_361) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_288), .A2(n_309), .B1(n_310), .B2(n_312), .Y(n_308) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g305 ( .A(n_291), .Y(n_305) );
INVx1_ASAP7_75t_L g309 ( .A(n_291), .Y(n_309) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_298), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g473 ( .A(n_299), .B(n_410), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_319), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_300), .B(n_358), .Y(n_581) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g460 ( .A(n_301), .B(n_321), .Y(n_460) );
AND2x2_ASAP7_75t_L g481 ( .A(n_301), .B(n_374), .Y(n_481) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_R g355 ( .A(n_302), .Y(n_355) );
INVx2_ASAP7_75t_L g412 ( .A(n_302), .Y(n_412) );
AND2x2_ASAP7_75t_L g462 ( .A(n_302), .B(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_302), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_302), .B(n_332), .Y(n_510) );
AND2x2_ASAP7_75t_L g515 ( .A(n_302), .B(n_431), .Y(n_515) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_315), .B(n_316), .Y(n_302) );
NOR3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_308), .C(n_314), .Y(n_303) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_307), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_315), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g411 ( .A(n_320), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g584 ( .A(n_320), .B(n_431), .Y(n_584) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g387 ( .A(n_321), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_321), .Y(n_428) );
INVx1_ASAP7_75t_L g463 ( .A(n_321), .Y(n_463) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_328), .Y(n_321) );
AND2x2_ASAP7_75t_L g375 ( .A(n_322), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_SL g480 ( .A(n_331), .Y(n_480) );
INVx1_ASAP7_75t_L g502 ( .A(n_331), .Y(n_502) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g357 ( .A(n_332), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_332), .Y(n_379) );
INVx1_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_332), .Y(n_410) );
AND2x4_ASAP7_75t_L g415 ( .A(n_332), .B(n_388), .Y(n_415) );
INVx2_ASAP7_75t_L g431 ( .A(n_332), .Y(n_431) );
AND2x2_ASAP7_75t_L g441 ( .A(n_332), .B(n_358), .Y(n_441) );
AO31x2_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_338), .A3(n_343), .B(n_344), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_340), .Y(n_600) );
OAI22xp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_353), .B1(n_371), .B2(n_380), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g381 ( .A(n_349), .B(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_349), .A2(n_434), .B1(n_438), .B2(n_444), .Y(n_433) );
AND2x4_ASAP7_75t_L g530 ( .A(n_349), .B(n_531), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_349), .B(n_498), .Y(n_575) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x4_ASAP7_75t_L g496 ( .A(n_351), .B(n_399), .Y(n_496) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g491 ( .A(n_352), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g565 ( .A(n_356), .B(n_462), .Y(n_565) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g469 ( .A(n_357), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_358), .B(n_412), .Y(n_432) );
AND2x2_ASAP7_75t_L g464 ( .A(n_358), .B(n_386), .Y(n_464) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g374 ( .A(n_360), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g588 ( .A1(n_371), .A2(n_589), .B(n_592), .Y(n_588) );
HB1xp67_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_379), .Y(n_372) );
OR2x2_ASAP7_75t_L g551 ( .A(n_373), .B(n_386), .Y(n_551) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g572 ( .A(n_374), .Y(n_572) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g446 ( .A(n_382), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g523 ( .A(n_382), .B(n_406), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_394), .B1(n_404), .B2(n_407), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x4_ASAP7_75t_L g508 ( .A(n_387), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g514 ( .A(n_387), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g452 ( .A(n_388), .Y(n_452) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_392), .Y(n_388) );
AND2x2_ASAP7_75t_L g596 ( .A(n_390), .B(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_397), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g593 ( .A(n_397), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g457 ( .A(n_398), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_403), .Y(n_399) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_404), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVxp67_ASAP7_75t_L g525 ( .A(n_409), .Y(n_525) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g414 ( .A(n_411), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g440 ( .A(n_411), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g447 ( .A(n_411), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g521 ( .A(n_411), .B(n_480), .Y(n_521) );
OAI31xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .A3(n_418), .B(n_420), .Y(n_413) );
INVx2_ASAP7_75t_L g425 ( .A(n_414), .Y(n_425) );
INVx2_ASAP7_75t_SL g443 ( .A(n_415), .Y(n_443) );
AND2x2_ASAP7_75t_L g459 ( .A(n_415), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g556 ( .A(n_415), .B(n_470), .Y(n_556) );
AND2x4_ASAP7_75t_L g576 ( .A(n_415), .B(n_462), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_415), .B(n_427), .Y(n_591) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_425), .C(n_426), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_422), .B(n_477), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_423), .A2(n_454), .B1(n_458), .B2(n_461), .Y(n_453) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
OR2x2_ASAP7_75t_L g442 ( .A(n_427), .B(n_443), .Y(n_442) );
AOI322xp5_ASAP7_75t_L g526 ( .A1(n_427), .A2(n_450), .A3(n_527), .B1(n_530), .B2(n_532), .C1(n_533), .C2(n_536), .Y(n_526) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g587 ( .A(n_429), .Y(n_587) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g563 ( .A(n_430), .Y(n_563) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g585 ( .A(n_432), .Y(n_585) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g536 ( .A(n_441), .B(n_462), .Y(n_536) );
INVx2_ASAP7_75t_L g542 ( .A(n_442), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_450), .B(n_453), .Y(n_445) );
INVx1_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
INVx1_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_449), .B(n_491), .Y(n_569) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_451), .B(n_493), .Y(n_532) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g594 ( .A(n_456), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_457), .A2(n_583), .B1(n_586), .B2(n_587), .Y(n_582) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g562 ( .A(n_460), .B(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_461), .A2(n_479), .B1(n_482), .B2(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx2_ASAP7_75t_SL g493 ( .A(n_462), .Y(n_493) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_466), .B(n_547), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_506), .C(n_526), .D(n_537), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .C(n_492), .Y(n_467) );
AOI21xp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_472), .B(n_474), .Y(n_468) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
NAND2x1p5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g500 ( .A(n_481), .Y(n_500) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_481), .Y(n_559) );
INVxp33_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI322xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .A3(n_495), .B1(n_497), .B2(n_500), .C1(n_501), .C2(n_503), .Y(n_492) );
OR2x2_ASAP7_75t_L g524 ( .A(n_493), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g507 ( .A(n_495), .Y(n_507) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_496), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g541 ( .A(n_498), .Y(n_541) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_502), .A2(n_512), .B(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g531 ( .A(n_505), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_505), .B(n_546), .Y(n_545) );
AOI221x1_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_511), .B2(n_516), .C(n_517), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g571 ( .A(n_510), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_514), .A2(n_549), .B(n_550), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .B1(n_522), .B2(n_524), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_519), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_521), .A2(n_538), .B1(n_542), .B2(n_543), .Y(n_537) );
OAI221xp5_ASAP7_75t_SL g577 ( .A1(n_522), .A2(n_571), .B1(n_578), .B2(n_579), .C(n_582), .Y(n_577) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_540), .B(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g544 ( .A(n_541), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_545), .Y(n_578) );
INVxp67_ASAP7_75t_L g568 ( .A(n_546), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_557), .C(n_573), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_554), .B2(n_555), .Y(n_550) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_560), .B2(n_566), .C(n_570), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g586 ( .A(n_569), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_577), .C(n_588), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
BUFx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OA21x2_ASAP7_75t_L g612 ( .A1(n_597), .A2(n_613), .B(n_614), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI222xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_607), .B2(n_609), .C1(n_611), .C2(n_615), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_616), .Y(n_615) );
endmodule