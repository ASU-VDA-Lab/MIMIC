module fake_ibex_235_n_93 (n_7, n_20, n_17, n_25, n_18, n_3, n_22, n_28, n_32, n_4, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_14, n_0, n_9, n_12, n_15, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_93);

input n_7;
input n_20;
input n_17;
input n_25;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_4;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_14;
input n_0;
input n_9;
input n_12;
input n_15;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_93;

wire n_85;
wire n_84;
wire n_64;
wire n_73;
wire n_65;
wire n_55;
wire n_63;
wire n_76;
wire n_67;
wire n_38;
wire n_37;
wire n_47;
wire n_82;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_75;
wire n_69;
wire n_48;
wire n_57;
wire n_59;
wire n_39;
wire n_62;
wire n_71;
wire n_61;
wire n_42;
wire n_77;
wire n_88;
wire n_44;
wire n_51;
wire n_46;
wire n_80;
wire n_49;
wire n_40;
wire n_66;
wire n_74;
wire n_90;
wire n_58;
wire n_43;
wire n_33;
wire n_72;
wire n_34;
wire n_52;
wire n_36;
wire n_41;
wire n_45;
wire n_89;
wire n_83;
wire n_53;
wire n_50;
wire n_92;
wire n_68;
wire n_79;
wire n_81;
wire n_35;
wire n_56;
wire n_91;
wire n_54;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_11),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_30),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_13),
.A2(n_16),
.B1(n_19),
.B2(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_49),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_55),
.B1(n_38),
.B2(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_44),
.Y(n_67)
);

NOR2x1p5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_44),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_48),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_54),
.B(n_42),
.C(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_65),
.B1(n_58),
.B2(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_76),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_69),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_72),
.C(n_84),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

AOI22x1_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_85),
.B1(n_68),
.B2(n_52),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_67),
.Y(n_93)
);


endmodule