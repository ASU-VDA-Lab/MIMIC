module fake_aes_4330_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_9), .B(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
OAI22xp5_ASAP7_75t_SL g15 ( .A1(n_0), .A2(n_3), .B1(n_8), .B2(n_2), .Y(n_15) );
AOI22xp33_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
AOI211xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_1), .B(n_3), .C(n_10), .Y(n_18) );
OAI21xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_11), .B(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NAND2x1_ASAP7_75t_L g24 ( .A(n_22), .B(n_12), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
INVxp67_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
AOI221xp5_ASAP7_75t_SL g28 ( .A1(n_26), .A2(n_19), .B1(n_21), .B2(n_16), .C(n_18), .Y(n_28) );
NAND4xp75_ASAP7_75t_L g29 ( .A(n_28), .B(n_12), .C(n_22), .D(n_27), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_28), .B(n_22), .Y(n_30) );
INVx1_ASAP7_75t_SL g31 ( .A(n_30), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OAI22xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_12), .B1(n_22), .B2(n_31), .Y(n_33) );
NAND2x1p5_ASAP7_75t_L g34 ( .A(n_33), .B(n_12), .Y(n_34) );
endmodule