module fake_jpeg_10327_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx6_ASAP7_75t_SL g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NAND3xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_15),
.C(n_16),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_0),
.C(n_1),
.Y(n_14)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_17),
.B(n_18),
.C(n_3),
.D(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_5),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_7),
.B1(n_10),
.B2(n_6),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_18),
.B(n_6),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_7),
.Y(n_26)
);

OA21x2_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_23),
.B(n_10),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_25),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_10),
.B1(n_13),
.B2(n_5),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_10),
.B(n_3),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_33),
.B(n_34),
.C(n_4),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_3),
.Y(n_34)
);

OAI31xp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_31),
.A3(n_32),
.B(n_29),
.Y(n_36)
);


endmodule