module fake_jpeg_30541_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_22),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_50),
.B1(n_42),
.B2(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_19),
.B1(n_31),
.B2(n_30),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_34),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_3),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_59),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_35),
.B(n_44),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_63),
.B(n_5),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_33),
.B1(n_43),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_70),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_77),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_76),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_79),
.B(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_89),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_24),
.C(n_25),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_92),
.C(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_81),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_83),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_65),
.B1(n_80),
.B2(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_92),
.C(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_98),
.B1(n_86),
.B2(n_85),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_105),
.Y(n_106)
);

NAND4xp25_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_98),
.C(n_94),
.D(n_103),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_100),
.Y(n_108)
);


endmodule