module real_jpeg_26638_n_23 (n_17, n_8, n_116, n_0, n_21, n_2, n_10, n_114, n_9, n_12, n_6, n_121, n_11, n_14, n_120, n_7, n_22, n_18, n_3, n_117, n_119, n_5, n_4, n_115, n_122, n_1, n_20, n_19, n_118, n_16, n_15, n_13, n_113, n_23);

input n_17;
input n_8;
input n_116;
input n_0;
input n_21;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_14;
input n_120;
input n_7;
input n_22;
input n_18;
input n_3;
input n_117;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_20;
input n_19;
input n_118;
input n_16;
input n_15;
input n_13;
input n_113;

output n_23;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_0),
.Y(n_109)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_2),
.B(n_35),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.C(n_104),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_4),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_6),
.B(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_7),
.B(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_8),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_9),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_11),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_11),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_12),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_12),
.B(n_74),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_16),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_16),
.B(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_17),
.B(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_18),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_19),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_20),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_43),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_86),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_28),
.B(n_97),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_28),
.B(n_109),
.Y(n_108)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_107),
.B(n_111),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B(n_106),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_100),
.B(n_103),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_95),
.B(n_99),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_90),
.C(n_94),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_89),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_88),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_83),
.B(n_87),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_82),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_77),
.B(n_81),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_73),
.B(n_76),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_72),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_66),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_75),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_79),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_110),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_113),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_114),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_115),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_116),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_117),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_118),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_119),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_120),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_121),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_122),
.Y(n_93)
);


endmodule