module real_aes_17062_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_0), .A2(n_70), .B1(n_563), .B2(n_691), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_0), .A2(n_257), .B1(n_429), .B2(n_432), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_1), .A2(n_214), .B1(n_432), .B2(n_958), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_1), .A2(n_59), .B1(n_354), .B2(n_985), .Y(n_1138) );
INVx1_ASAP7_75t_L g1033 ( .A(n_2), .Y(n_1033) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_3), .A2(n_654), .B(n_656), .C(n_669), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_3), .B(n_314), .Y(n_685) );
INVx1_ASAP7_75t_L g974 ( .A(n_4), .Y(n_974) );
AOI22xp5_ASAP7_75t_SL g1227 ( .A1(n_5), .A2(n_264), .B1(n_1210), .B2(n_1218), .Y(n_1227) );
INVx1_ASAP7_75t_L g1129 ( .A(n_6), .Y(n_1129) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_6), .A2(n_62), .B1(n_705), .B2(n_837), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_7), .A2(n_73), .B1(n_691), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_7), .A2(n_45), .B1(n_889), .B2(n_890), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g1424 ( .A1(n_8), .A2(n_145), .B1(n_365), .B2(n_1425), .Y(n_1424) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_8), .Y(n_1447) );
INVx1_ASAP7_75t_L g737 ( .A(n_9), .Y(n_737) );
AO22x1_ASAP7_75t_L g763 ( .A1(n_9), .A2(n_142), .B1(n_417), .B2(n_665), .Y(n_763) );
INVx1_ASAP7_75t_L g295 ( .A(n_10), .Y(n_295) );
AND2x2_ASAP7_75t_L g346 ( .A(n_10), .B(n_235), .Y(n_346) );
AND2x2_ASAP7_75t_L g407 ( .A(n_10), .B(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_10), .B(n_305), .Y(n_522) );
INVx1_ASAP7_75t_L g747 ( .A(n_11), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_11), .A2(n_100), .B1(n_422), .B2(n_661), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_12), .A2(n_144), .B1(n_553), .B2(n_1024), .C(n_1028), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_12), .A2(n_53), .B1(n_432), .B2(n_806), .Y(n_1040) );
INVx1_ASAP7_75t_L g924 ( .A(n_13), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g943 ( .A1(n_13), .A2(n_157), .B1(n_944), .B2(n_945), .C(n_946), .Y(n_943) );
INVx2_ASAP7_75t_L g1205 ( .A(n_14), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_14), .B(n_1206), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_14), .B(n_105), .Y(n_1213) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_15), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_16), .Y(n_1167) );
AOI22xp5_ASAP7_75t_SL g1241 ( .A1(n_17), .A2(n_132), .B1(n_1210), .B2(n_1218), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_18), .A2(n_41), .B1(n_380), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_18), .A2(n_278), .B1(n_889), .B2(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1172 ( .A(n_19), .Y(n_1172) );
AOI22xp5_ASAP7_75t_SL g1236 ( .A1(n_20), .A2(n_253), .B1(n_1207), .B2(n_1212), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_21), .A2(n_154), .B1(n_369), .B2(n_374), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_21), .A2(n_233), .B1(n_440), .B2(n_444), .C(n_448), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g670 ( .A1(n_22), .A2(n_671), .B(n_673), .C(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g716 ( .A(n_22), .Y(n_716) );
INVx1_ASAP7_75t_L g972 ( .A(n_23), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_23), .A2(n_138), .B1(n_945), .B2(n_998), .C(n_999), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_24), .A2(n_98), .B1(n_314), .B2(n_1043), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1489 ( .A1(n_25), .A2(n_115), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1498 ( .A1(n_25), .A2(n_279), .B1(n_1499), .B2(n_1502), .Y(n_1498) );
AOI22xp33_ASAP7_75t_SL g978 ( .A1(n_26), .A2(n_278), .B1(n_979), .B2(n_980), .Y(n_978) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_26), .A2(n_41), .B1(n_661), .B2(n_663), .C(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_27), .A2(n_90), .B1(n_388), .B2(n_827), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_27), .A2(n_165), .B1(n_426), .B2(n_440), .C(n_885), .Y(n_959) );
NAND2xp5_ASAP7_75t_SL g807 ( .A(n_28), .B(n_421), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_28), .A2(n_159), .B1(n_388), .B2(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1484 ( .A(n_29), .Y(n_1484) );
INVx1_ASAP7_75t_L g409 ( .A(n_30), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_31), .A2(n_159), .B1(n_417), .B2(n_658), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_31), .A2(n_251), .B1(n_388), .B2(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g1114 ( .A(n_32), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1201 ( .A1(n_33), .A2(n_180), .B1(n_1202), .B2(n_1207), .Y(n_1201) );
XOR2x2_ASAP7_75t_L g1046 ( .A(n_34), .B(n_1047), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_34), .A2(n_95), .B1(n_1210), .B2(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g594 ( .A(n_35), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g1209 ( .A1(n_36), .A2(n_183), .B1(n_1210), .B2(n_1212), .Y(n_1209) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_37), .A2(n_87), .B1(n_1202), .B2(n_1210), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_38), .A2(n_233), .B1(n_369), .B2(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_38), .A2(n_154), .B1(n_429), .B2(n_431), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_39), .A2(n_60), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_39), .A2(n_274), .B1(n_365), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_40), .A2(n_128), .B1(n_869), .B2(n_870), .Y(n_868) );
INVxp67_ASAP7_75t_SL g907 ( .A(n_40), .Y(n_907) );
INVx1_ASAP7_75t_L g321 ( .A(n_42), .Y(n_321) );
INVx1_ASAP7_75t_L g338 ( .A(n_42), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_43), .A2(n_123), .B1(n_365), .B2(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_43), .A2(n_68), .B1(n_421), .B2(n_424), .C(n_426), .Y(n_420) );
INVx1_ASAP7_75t_L g792 ( .A(n_44), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_45), .A2(n_133), .B1(n_691), .B2(n_865), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_46), .A2(n_272), .B1(n_1202), .B2(n_1207), .Y(n_1221) );
INVx1_ASAP7_75t_L g1483 ( .A(n_47), .Y(n_1483) );
INVx1_ASAP7_75t_L g975 ( .A(n_48), .Y(n_975) );
INVx1_ASAP7_75t_L g288 ( .A(n_49), .Y(n_288) );
INVx2_ASAP7_75t_L g324 ( .A(n_50), .Y(n_324) );
INVx1_ASAP7_75t_L g782 ( .A(n_51), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g967 ( .A(n_52), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_53), .A2(n_67), .B1(n_367), .B2(n_1024), .C(n_1025), .Y(n_1023) );
INVx1_ASAP7_75t_L g874 ( .A(n_54), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_55), .A2(n_120), .B1(n_887), .B2(n_1053), .C(n_1055), .Y(n_1052) );
INVx1_ASAP7_75t_L g1098 ( .A(n_55), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1237 ( .A1(n_56), .A2(n_63), .B1(n_1202), .B2(n_1210), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_57), .A2(n_215), .B1(n_440), .B2(n_958), .Y(n_1532) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_57), .A2(n_89), .B1(n_374), .B2(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1017 ( .A(n_58), .Y(n_1017) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_59), .A2(n_202), .B1(n_426), .B2(n_1037), .C(n_1123), .Y(n_1122) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_60), .A2(n_99), .B1(n_365), .B2(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g1016 ( .A(n_61), .Y(n_1016) );
INVx1_ASAP7_75t_L g1128 ( .A(n_62), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1428 ( .A1(n_64), .A2(n_66), .B1(n_365), .B2(n_367), .Y(n_1428) );
AOI221xp5_ASAP7_75t_L g1436 ( .A1(n_64), .A2(n_145), .B1(n_424), .B2(n_887), .C(n_1437), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_65), .A2(n_126), .B1(n_429), .B2(n_1057), .Y(n_1061) );
INVx1_ASAP7_75t_L g1085 ( .A(n_65), .Y(n_1085) );
INVxp67_ASAP7_75t_SL g1449 ( .A(n_66), .Y(n_1449) );
AOI221xp5_ASAP7_75t_L g1036 ( .A1(n_67), .A2(n_144), .B1(n_446), .B2(n_668), .C(n_1037), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_68), .A2(n_227), .B1(n_365), .B2(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g835 ( .A(n_69), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_70), .A2(n_77), .B1(n_446), .B2(n_628), .C(n_953), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g1160 ( .A1(n_71), .A2(n_188), .B1(n_388), .B2(n_860), .Y(n_1160) );
AOI22xp33_ASAP7_75t_SL g1188 ( .A1(n_71), .A2(n_243), .B1(n_429), .B2(n_995), .Y(n_1188) );
AOI22xp33_ASAP7_75t_SL g1426 ( .A1(n_72), .A2(n_191), .B1(n_865), .B2(n_930), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_72), .A2(n_129), .B1(n_429), .B2(n_431), .Y(n_1439) );
INVx1_ASAP7_75t_L g902 ( .A(n_73), .Y(n_902) );
INVx1_ASAP7_75t_L g620 ( .A(n_74), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_74), .A2(n_124), .B1(n_425), .B2(n_628), .C(n_635), .Y(n_634) );
AOI21xp33_ASAP7_75t_L g1117 ( .A1(n_75), .A2(n_448), .B(n_1063), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_75), .A2(n_176), .B1(n_563), .B2(n_707), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_76), .A2(n_221), .B1(n_460), .B2(n_779), .Y(n_968) );
OAI211xp5_ASAP7_75t_L g987 ( .A1(n_76), .A2(n_955), .B(n_988), .C(n_996), .Y(n_987) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_77), .A2(n_257), .B1(n_563), .B2(n_691), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1429 ( .A1(n_78), .A2(n_267), .B1(n_837), .B2(n_937), .Y(n_1429) );
INVx1_ASAP7_75t_L g1442 ( .A(n_78), .Y(n_1442) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_79), .A2(n_179), .B1(n_380), .B2(n_557), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_79), .A2(n_88), .B1(n_890), .B2(n_958), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g1217 ( .A1(n_80), .A2(n_190), .B1(n_1207), .B2(n_1218), .Y(n_1217) );
OAI222xp33_ASAP7_75t_L g753 ( .A1(n_81), .A2(n_216), .B1(n_575), .B2(n_577), .C1(n_754), .C2(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g766 ( .A(n_81), .Y(n_766) );
OAI211xp5_ASAP7_75t_L g1112 ( .A1(n_82), .A2(n_998), .B(n_1113), .C(n_1115), .Y(n_1112) );
INVx1_ASAP7_75t_L g1136 ( .A(n_82), .Y(n_1136) );
INVx1_ASAP7_75t_L g853 ( .A(n_83), .Y(n_853) );
OAI222xp33_ASAP7_75t_L g893 ( .A1(n_83), .A2(n_122), .B1(n_894), .B2(n_897), .C1(n_903), .C2(n_910), .Y(n_893) );
OAI22xp5_ASAP7_75t_SL g800 ( .A1(n_84), .A2(n_102), .B1(n_801), .B2(n_802), .Y(n_800) );
OAI21xp33_ASAP7_75t_L g815 ( .A1(n_84), .A2(n_705), .B(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g1066 ( .A(n_85), .Y(n_1066) );
INVx1_ASAP7_75t_L g331 ( .A(n_86), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_88), .A2(n_110), .B1(n_380), .B2(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g1541 ( .A1(n_89), .A2(n_203), .B1(n_958), .B2(n_1057), .Y(n_1541) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_90), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_91), .Y(n_742) );
INVx1_ASAP7_75t_L g520 ( .A(n_92), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_92), .A2(n_225), .B1(n_553), .B2(n_555), .C(n_558), .Y(n_552) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_93), .Y(n_290) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_93), .B(n_288), .Y(n_1203) );
AOI22xp33_ASAP7_75t_SL g1161 ( .A1(n_94), .A2(n_281), .B1(n_549), .B2(n_1162), .Y(n_1161) );
AOI21xp33_ASAP7_75t_L g1186 ( .A1(n_94), .A2(n_953), .B(n_1187), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_96), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_97), .Y(n_1020) );
OAI211xp5_ASAP7_75t_SL g1119 ( .A1(n_98), .A2(n_1120), .B(n_1121), .C(n_1127), .Y(n_1119) );
AOI221xp5_ASAP7_75t_SL g666 ( .A1(n_99), .A2(n_274), .B1(n_422), .B2(n_667), .C(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g743 ( .A(n_100), .Y(n_743) );
OAI211xp5_ASAP7_75t_L g794 ( .A1(n_101), .A2(n_795), .B(n_796), .C(n_797), .Y(n_794) );
INVxp33_ASAP7_75t_SL g817 ( .A(n_101), .Y(n_817) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_102), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_103), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_104), .A2(n_265), .B1(n_936), .B2(n_937), .Y(n_1173) );
INVx1_ASAP7_75t_L g1181 ( .A(n_104), .Y(n_1181) );
INVx1_ASAP7_75t_L g1206 ( .A(n_105), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_105), .B(n_1205), .Y(n_1211) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_106), .A2(n_238), .B1(n_583), .B2(n_586), .Y(n_582) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_106), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_107), .A2(n_189), .B1(n_1202), .B2(n_1207), .Y(n_1228) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_108), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g1531 ( .A1(n_109), .A2(n_130), .B1(n_424), .B2(n_431), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_109), .A2(n_169), .B1(n_982), .B2(n_1544), .Y(n_1543) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_110), .A2(n_179), .B1(n_950), .B2(n_951), .C(n_953), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_111), .A2(n_171), .B1(n_936), .B2(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g962 ( .A(n_111), .Y(n_962) );
INVx1_ASAP7_75t_L g1069 ( .A(n_112), .Y(n_1069) );
INVx2_ASAP7_75t_L g326 ( .A(n_113), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_113), .B(n_324), .Y(n_341) );
INVx1_ASAP7_75t_L g386 ( .A(n_113), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_114), .A2(n_152), .B1(n_376), .B2(n_562), .Y(n_624) );
INVx1_ASAP7_75t_L g636 ( .A(n_114), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g1518 ( .A1(n_115), .A2(n_275), .B1(n_1519), .B2(n_1522), .Y(n_1518) );
INVx1_ASAP7_75t_L g533 ( .A(n_116), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_117), .A2(n_146), .B1(n_487), .B2(n_493), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_117), .A2(n_213), .B1(n_561), .B2(n_563), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_118), .A2(n_136), .B1(n_671), .B2(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g702 ( .A(n_118), .Y(n_702) );
INVx1_ASAP7_75t_L g751 ( .A(n_119), .Y(n_751) );
NAND2xp33_ASAP7_75t_SL g775 ( .A(n_119), .B(n_422), .Y(n_775) );
INVx1_ASAP7_75t_L g1086 ( .A(n_120), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_121), .B(n_333), .Y(n_1104) );
INVx1_ASAP7_75t_L g851 ( .A(n_122), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_123), .A2(n_227), .B1(n_431), .B2(n_438), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_124), .A2(n_249), .B1(n_355), .B2(n_614), .C(n_615), .Y(n_613) );
XNOR2xp5_ASAP7_75t_L g595 ( .A(n_125), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g1094 ( .A(n_126), .Y(n_1094) );
XOR2x2_ASAP7_75t_L g918 ( .A(n_127), .B(n_919), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_128), .A2(n_269), .B1(n_883), .B2(n_885), .C(n_887), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_129), .A2(n_245), .B1(n_865), .B2(n_930), .Y(n_1427) );
AOI22xp33_ASAP7_75t_SL g1549 ( .A1(n_130), .A2(n_234), .B1(n_696), .B2(n_985), .Y(n_1549) );
AOI22xp33_ASAP7_75t_SL g984 ( .A1(n_131), .A2(n_148), .B1(n_367), .B2(n_985), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_131), .A2(n_185), .B1(n_887), .B2(n_990), .C(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g898 ( .A(n_133), .Y(n_898) );
INVxp67_ASAP7_75t_SL g1158 ( .A(n_134), .Y(n_1158) );
OAI211xp5_ASAP7_75t_L g1175 ( .A1(n_134), .A2(n_955), .B(n_1176), .C(n_1180), .Y(n_1175) );
AOI22xp33_ASAP7_75t_SL g1164 ( .A1(n_135), .A2(n_260), .B1(n_549), .B2(n_1162), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_135), .A2(n_281), .B1(n_432), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g714 ( .A(n_136), .Y(n_714) );
INVx1_ASAP7_75t_L g1255 ( .A(n_137), .Y(n_1255) );
INVx1_ASAP7_75t_L g971 ( .A(n_138), .Y(n_971) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_139), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_140), .A2(n_270), .B1(n_583), .B2(n_586), .Y(n_603) );
INVxp33_ASAP7_75t_SL g645 ( .A(n_140), .Y(n_645) );
NAND5xp2_ASAP7_75t_L g651 ( .A(n_141), .B(n_652), .C(n_686), .D(n_703), .E(n_711), .Y(n_651) );
INVx1_ASAP7_75t_L g720 ( .A(n_141), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_142), .A2(n_551), .B(n_562), .Y(n_752) );
INVx1_ASAP7_75t_L g777 ( .A(n_143), .Y(n_777) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_146), .A2(n_261), .B1(n_547), .B2(n_549), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_147), .A2(n_174), .B1(n_460), .B2(n_779), .Y(n_1432) );
OAI211xp5_ASAP7_75t_SL g1434 ( .A1(n_147), .A2(n_1120), .B(n_1435), .C(n_1440), .Y(n_1434) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_148), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_149), .A2(n_186), .B1(n_1210), .B2(n_1257), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1459 ( .A1(n_149), .A2(n_1460), .B1(n_1463), .B2(n_1552), .Y(n_1459) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_149), .A2(n_1466), .B1(n_1550), .B2(n_1551), .Y(n_1465) );
INVxp67_ASAP7_75t_SL g1551 ( .A(n_149), .Y(n_1551) );
INVx1_ASAP7_75t_L g1155 ( .A(n_150), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1183 ( .A1(n_150), .A2(n_153), .B1(n_911), .B2(n_944), .C(n_1184), .Y(n_1183) );
BUFx3_ASAP7_75t_L g318 ( .A(n_151), .Y(n_318) );
INVx1_ASAP7_75t_L g630 ( .A(n_152), .Y(n_630) );
INVx1_ASAP7_75t_L g1156 ( .A(n_153), .Y(n_1156) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_155), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_156), .A2(n_243), .B1(n_388), .B2(n_869), .Y(n_1165) );
AOI221xp5_ASAP7_75t_L g1177 ( .A1(n_156), .A2(n_188), .B1(n_425), .B2(n_426), .C(n_1037), .Y(n_1177) );
INVx1_ASAP7_75t_L g923 ( .A(n_157), .Y(n_923) );
INVx1_ASAP7_75t_L g610 ( .A(n_158), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_158), .A2(n_206), .B1(n_425), .B2(n_628), .C(n_629), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g1259 ( .A1(n_160), .A2(n_204), .B1(n_1202), .B2(n_1207), .Y(n_1259) );
INVx1_ASAP7_75t_L g1074 ( .A(n_161), .Y(n_1074) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_162), .A2(n_460), .B(n_873), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g1222 ( .A1(n_163), .A2(n_222), .B1(n_1210), .B2(n_1218), .Y(n_1222) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_164), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g926 ( .A1(n_165), .A2(n_241), .B1(n_367), .B2(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g598 ( .A(n_166), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_167), .A2(n_212), .B1(n_659), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_167), .A2(n_205), .B1(n_563), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g1034 ( .A(n_168), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g1536 ( .A1(n_169), .A2(n_234), .B1(n_1537), .B2(n_1538), .Y(n_1536) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_170), .Y(n_390) );
INVx1_ASAP7_75t_L g961 ( .A(n_171), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_172), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_173), .A2(n_213), .B1(n_493), .B2(n_516), .C(n_518), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_173), .A2(n_219), .B1(n_365), .B2(n_388), .C(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g977 ( .A1(n_175), .A2(n_185), .B1(n_365), .B2(n_870), .Y(n_977) );
INVx1_ASAP7_75t_L g1000 ( .A(n_175), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_176), .A2(n_255), .B1(n_432), .B2(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1479 ( .A(n_177), .Y(n_1479) );
OAI211xp5_ASAP7_75t_L g1506 ( .A1(n_177), .A2(n_1507), .B(n_1508), .C(n_1510), .Y(n_1506) );
OAI21xp5_ASAP7_75t_SL g1042 ( .A1(n_178), .A2(n_1043), .B(n_1044), .Y(n_1042) );
INVx1_ASAP7_75t_L g618 ( .A(n_181), .Y(n_618) );
INVx1_ASAP7_75t_L g875 ( .A(n_182), .Y(n_875) );
INVx1_ASAP7_75t_L g730 ( .A(n_184), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_184), .B(n_583), .Y(n_732) );
INVx1_ASAP7_75t_L g856 ( .A(n_187), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g1450 ( .A1(n_191), .A2(n_245), .B1(n_883), .B2(n_885), .C(n_1065), .Y(n_1450) );
AOI22xp5_ASAP7_75t_L g1415 ( .A1(n_192), .A2(n_1416), .B1(n_1453), .B2(n_1454), .Y(n_1415) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_192), .Y(n_1453) );
AOI21xp33_ASAP7_75t_L g812 ( .A1(n_193), .A2(n_425), .B(n_663), .Y(n_812) );
INVx1_ASAP7_75t_L g823 ( .A(n_193), .Y(n_823) );
INVx1_ASAP7_75t_L g710 ( .A(n_194), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_195), .Y(n_350) );
OAI211xp5_ASAP7_75t_L g1050 ( .A1(n_196), .A2(n_894), .B(n_1051), .C(n_1058), .Y(n_1050) );
INVx1_ASAP7_75t_L g1101 ( .A(n_196), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_197), .A2(n_259), .B1(n_1037), .B2(n_1063), .C(n_1065), .Y(n_1062) );
INVx1_ASAP7_75t_L g1077 ( .A(n_197), .Y(n_1077) );
INVx1_ASAP7_75t_L g1071 ( .A(n_198), .Y(n_1071) );
OAI332xp33_ASAP7_75t_SL g1075 ( .A1(n_198), .A2(n_698), .A3(n_837), .B1(n_1076), .B2(n_1082), .B3(n_1083), .C1(n_1089), .C2(n_1093), .Y(n_1075) );
INVx1_ASAP7_75t_L g403 ( .A(n_199), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_200), .Y(n_940) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_201), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_202), .A2(n_214), .B1(n_367), .B2(n_985), .Y(n_1140) );
AOI22xp33_ASAP7_75t_SL g1545 ( .A1(n_203), .A2(n_215), .B1(n_863), .B2(n_985), .Y(n_1545) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_205), .A2(n_248), .B1(n_422), .B2(n_661), .C(n_663), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_206), .A2(n_557), .B(n_558), .Y(n_623) );
INVx1_ASAP7_75t_L g395 ( .A(n_207), .Y(n_395) );
XOR2x2_ASAP7_75t_L g787 ( .A(n_208), .B(n_788), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_209), .A2(n_263), .B1(n_417), .B2(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g825 ( .A(n_209), .Y(n_825) );
INVxp67_ASAP7_75t_SL g1116 ( .A(n_210), .Y(n_1116) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_210), .A2(n_255), .B1(n_371), .B2(n_980), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g1431 ( .A(n_211), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_212), .A2(n_248), .B1(n_563), .B2(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_R g768 ( .A(n_216), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_217), .B(n_1151), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_217), .A2(n_1169), .B1(n_1170), .B2(n_1189), .Y(n_1168) );
INVx1_ASAP7_75t_L g1191 ( .A(n_217), .Y(n_1191) );
OA22x2_ASAP7_75t_L g1109 ( .A1(n_218), .A2(n_1110), .B1(n_1144), .B2(n_1145), .Y(n_1109) );
CKINVDCx16_ASAP7_75t_R g1144 ( .A(n_218), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_219), .A2(n_225), .B1(n_497), .B2(n_500), .C(n_504), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_220), .A2(n_236), .B1(n_460), .B2(n_779), .Y(n_941) );
INVx1_ASAP7_75t_L g725 ( .A(n_222), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_223), .A2(n_242), .B1(n_429), .B2(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1092 ( .A(n_223), .Y(n_1092) );
INVx1_ASAP7_75t_L g1421 ( .A(n_224), .Y(n_1421) );
OAI221xp5_ASAP7_75t_SL g1445 ( .A1(n_224), .A2(n_276), .B1(n_910), .B2(n_998), .C(n_1446), .Y(n_1445) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_226), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_226), .A2(n_230), .B1(n_575), .B2(n_577), .C(n_579), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_228), .A2(n_269), .B1(n_553), .B2(n_860), .Y(n_859) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_228), .Y(n_904) );
OAI211xp5_ASAP7_75t_SL g604 ( .A1(n_229), .A2(n_572), .B(n_579), .C(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g641 ( .A(n_229), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_230), .A2(n_240), .B1(n_507), .B2(n_512), .C(n_513), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_231), .Y(n_799) );
INVx1_ASAP7_75t_L g1068 ( .A(n_232), .Y(n_1068) );
BUFx3_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
INVx1_ASAP7_75t_L g408 ( .A(n_235), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g954 ( .A1(n_236), .A2(n_955), .B(n_956), .C(n_960), .Y(n_954) );
XOR2x2_ASAP7_75t_L g964 ( .A(n_237), .B(n_965), .Y(n_964) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_238), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_239), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_240), .A2(n_244), .B1(n_565), .B2(n_568), .Y(n_564) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_241), .Y(n_947) );
INVx1_ASAP7_75t_L g1079 ( .A(n_242), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_244), .Y(n_539) );
INVx1_ASAP7_75t_L g330 ( .A(n_246), .Y(n_330) );
INVx1_ASAP7_75t_L g344 ( .A(n_246), .Y(n_344) );
INVx2_ASAP7_75t_L g363 ( .A(n_246), .Y(n_363) );
XNOR2x1_ASAP7_75t_L g1013 ( .A(n_247), .B(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g631 ( .A(n_249), .Y(n_631) );
INVx1_ASAP7_75t_L g740 ( .A(n_250), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_250), .A2(n_280), .B1(n_659), .B2(n_665), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_251), .B(n_425), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g1240 ( .A1(n_252), .A2(n_271), .B1(n_1202), .B2(n_1207), .Y(n_1240) );
INVx1_ASAP7_75t_L g475 ( .A(n_254), .Y(n_475) );
INVx1_ASAP7_75t_L g1131 ( .A(n_256), .Y(n_1131) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_258), .A2(n_460), .B(n_469), .Y(n_459) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_259), .Y(n_1090) );
INVx1_ASAP7_75t_L g1185 ( .A(n_260), .Y(n_1185) );
INVx1_ASAP7_75t_L g519 ( .A(n_261), .Y(n_519) );
INVx1_ASAP7_75t_L g1253 ( .A(n_262), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g831 ( .A(n_263), .Y(n_831) );
INVx1_ASAP7_75t_L g1182 ( .A(n_265), .Y(n_1182) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_266), .Y(n_612) );
INVx1_ASAP7_75t_L g1441 ( .A(n_267), .Y(n_1441) );
INVx1_ASAP7_75t_L g914 ( .A(n_268), .Y(n_914) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_270), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_273), .Y(n_798) );
INVx1_ASAP7_75t_L g1477 ( .A(n_275), .Y(n_1477) );
INVx1_ASAP7_75t_L g1422 ( .A(n_276), .Y(n_1422) );
INVx1_ASAP7_75t_L g809 ( .A(n_277), .Y(n_809) );
INVx1_ASAP7_75t_L g1472 ( .A(n_279), .Y(n_1472) );
INVx1_ASAP7_75t_L g749 ( .A(n_280), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_306), .B(n_1192), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1462 ( .A(n_285), .B(n_294), .Y(n_1462) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1458 ( .A(n_287), .B(n_290), .Y(n_1458) );
INVx1_ASAP7_75t_L g1553 ( .A(n_287), .Y(n_1553) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_290), .B(n_1553), .Y(n_1555) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g1495 ( .A(n_294), .B(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g427 ( .A(n_295), .B(n_305), .Y(n_427) );
AND2x4_ASAP7_75t_L g449 ( .A(n_295), .B(n_304), .Y(n_449) );
AND2x4_ASAP7_75t_SL g1461 ( .A(n_296), .B(n_1462), .Y(n_1461) );
INVxp67_ASAP7_75t_SL g1490 ( .A(n_296), .Y(n_1490) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g495 ( .A(n_299), .Y(n_495) );
BUFx4f_ASAP7_75t_L g672 ( .A(n_299), .Y(n_672) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
AND2x2_ASAP7_75t_L g413 ( .A(n_301), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g419 ( .A(n_301), .Y(n_419) );
AND2x2_ASAP7_75t_L g423 ( .A(n_301), .B(n_302), .Y(n_423) );
INVx1_ASAP7_75t_L g464 ( .A(n_301), .Y(n_464) );
NAND2x1_ASAP7_75t_L g503 ( .A(n_301), .B(n_302), .Y(n_503) );
INVx1_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
INVx2_ASAP7_75t_L g414 ( .A(n_302), .Y(n_414) );
AND2x2_ASAP7_75t_L g418 ( .A(n_302), .B(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g454 ( .A(n_302), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_302), .B(n_419), .Y(n_492) );
OR2x2_ASAP7_75t_L g499 ( .A(n_302), .B(n_348), .Y(n_499) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g1488 ( .A(n_304), .Y(n_1488) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g1471 ( .A(n_305), .Y(n_1471) );
AND2x4_ASAP7_75t_L g1482 ( .A(n_305), .B(n_463), .Y(n_1482) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_1007), .B2(n_1008), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
XNOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_477), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_310) );
INVx1_ASAP7_75t_L g476 ( .A(n_311), .Y(n_476) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_400), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_331), .B1(n_332), .B2(n_350), .C(n_351), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_313), .A2(n_332), .B1(n_1016), .B2(n_1017), .C(n_1018), .Y(n_1015) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx5_ASAP7_75t_L g843 ( .A(n_314), .Y(n_843) );
OR2x6_ASAP7_75t_L g314 ( .A(n_315), .B(n_327), .Y(n_314) );
INVx2_ASAP7_75t_L g573 ( .A(n_315), .Y(n_573) );
OR2x2_ASAP7_75t_L g779 ( .A(n_315), .B(n_327), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_316), .B(n_322), .Y(n_315) );
INVx8_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
BUFx3_ASAP7_75t_L g562 ( .A(n_316), .Y(n_562) );
AND2x2_ASAP7_75t_L g566 ( .A(n_316), .B(n_567), .Y(n_566) );
BUFx3_ASAP7_75t_L g827 ( .A(n_316), .Y(n_827) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_316), .Y(n_833) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x4_ASAP7_75t_L g372 ( .A(n_317), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_318), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g355 ( .A(n_318), .B(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_318), .Y(n_377) );
OR2x2_ASAP7_75t_L g736 ( .A(n_318), .B(n_320), .Y(n_736) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g373 ( .A(n_321), .Y(n_373) );
AND2x4_ASAP7_75t_L g357 ( .A(n_322), .B(n_343), .Y(n_357) );
AND2x6_ASAP7_75t_L g576 ( .A(n_322), .B(n_393), .Y(n_576) );
AND2x2_ASAP7_75t_L g578 ( .A(n_322), .B(n_399), .Y(n_578) );
INVx1_ASAP7_75t_L g581 ( .A(n_322), .Y(n_581) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NAND3x1_ASAP7_75t_L g384 ( .A(n_323), .B(n_385), .C(n_386), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_323), .B(n_386), .Y(n_551) );
INVx1_ASAP7_75t_L g1501 ( .A(n_323), .Y(n_1501) );
OR2x6_ASAP7_75t_L g1504 ( .A(n_323), .B(n_1505), .Y(n_1504) );
AND2x4_ASAP7_75t_L g1509 ( .A(n_323), .B(n_355), .Y(n_1509) );
OR2x4_ASAP7_75t_L g1521 ( .A(n_323), .B(n_736), .Y(n_1521) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
NAND2xp33_ASAP7_75t_SL g559 ( .A(n_324), .B(n_326), .Y(n_559) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND3x4_ASAP7_75t_L g360 ( .A(n_326), .B(n_361), .C(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g744 ( .A(n_326), .B(n_361), .Y(n_744) );
HB1xp67_ASAP7_75t_L g1526 ( .A(n_326), .Y(n_1526) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g461 ( .A(n_328), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g512 ( .A(n_328), .B(n_462), .Y(n_512) );
INVx1_ASAP7_75t_L g543 ( .A(n_328), .Y(n_543) );
INVx1_ASAP7_75t_L g1496 ( .A(n_328), .Y(n_1496) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g340 ( .A(n_329), .Y(n_340) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_331), .A2(n_416), .B1(n_420), .B2(n_428), .C(n_433), .Y(n_415) );
AOI211x1_ASAP7_75t_L g846 ( .A1(n_332), .A2(n_847), .B(n_848), .C(n_872), .Y(n_846) );
AOI21xp33_ASAP7_75t_SL g939 ( .A1(n_332), .A2(n_940), .B(n_941), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g966 ( .A1(n_332), .A2(n_967), .B(n_968), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_332), .A2(n_1131), .B(n_1132), .Y(n_1130) );
NAND2xp33_ASAP7_75t_L g1166 ( .A(n_332), .B(n_1167), .Y(n_1166) );
AOI21xp5_ASAP7_75t_L g1430 ( .A1(n_332), .A2(n_1431), .B(n_1432), .Y(n_1430) );
INVx8_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_342), .Y(n_333) );
INVx1_ASAP7_75t_L g715 ( .A(n_334), .Y(n_715) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
BUFx3_ASAP7_75t_L g611 ( .A(n_335), .Y(n_611) );
INVx1_ASAP7_75t_L g1081 ( .A(n_335), .Y(n_1081) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_336), .Y(n_739) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g1505 ( .A(n_337), .Y(n_1505) );
INVx2_ASAP7_75t_L g356 ( .A(n_338), .Y(n_356) );
INVx1_ASAP7_75t_L g468 ( .A(n_338), .Y(n_468) );
OR2x2_ASAP7_75t_L g465 ( .A(n_339), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g472 ( .A(n_339), .Y(n_472) );
INVx1_ASAP7_75t_L g708 ( .A(n_339), .Y(n_708) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_340), .B(n_427), .Y(n_505) );
INVx1_ASAP7_75t_L g639 ( .A(n_340), .Y(n_639) );
OR2x2_ASAP7_75t_L g821 ( .A(n_340), .B(n_559), .Y(n_821) );
HB1xp67_ASAP7_75t_L g1528 ( .A(n_340), .Y(n_1528) );
INVx1_ASAP7_75t_L g567 ( .A(n_341), .Y(n_567) );
INVx1_ASAP7_75t_L g585 ( .A(n_341), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_342), .B(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g525 ( .A(n_343), .Y(n_525) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_344), .B(n_407), .Y(n_530) );
INVx1_ASAP7_75t_L g526 ( .A(n_345), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AND2x6_ASAP7_75t_L g433 ( .A(n_346), .B(n_422), .Y(n_433) );
AND2x2_ASAP7_75t_L g452 ( .A(n_346), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_346), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_346), .B(n_363), .Y(n_509) );
INVx1_ASAP7_75t_L g681 ( .A(n_346), .Y(n_681) );
AND2x2_ASAP7_75t_L g406 ( .A(n_347), .B(n_407), .Y(n_406) );
INVx3_ASAP7_75t_L g430 ( .A(n_347), .Y(n_430) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_347), .Y(n_658) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_348), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g351 ( .A(n_352), .B(n_358), .C(n_389), .Y(n_351) );
AND5x1_ASAP7_75t_L g788 ( .A(n_352), .B(n_789), .C(n_818), .D(n_834), .E(n_841), .Y(n_788) );
INVx2_ASAP7_75t_SL g938 ( .A(n_352), .Y(n_938) );
NAND4xp75_ASAP7_75t_L g965 ( .A(n_352), .B(n_966), .C(n_969), .D(n_986), .Y(n_965) );
NAND3xp33_ASAP7_75t_SL g1018 ( .A(n_352), .B(n_1019), .C(n_1022), .Y(n_1018) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_353), .A2(n_676), .B1(n_700), .B2(n_701), .C(n_702), .Y(n_699) );
INVx3_ASAP7_75t_L g857 ( .A(n_353), .Y(n_857) );
NOR3xp33_ASAP7_75t_L g1133 ( .A(n_353), .B(n_1134), .C(n_1143), .Y(n_1133) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
BUFx2_ASAP7_75t_L g1425 ( .A(n_354), .Y(n_1425) );
BUFx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g367 ( .A(n_355), .Y(n_367) );
BUFx3_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
INVx2_ASAP7_75t_L g554 ( .A(n_355), .Y(n_554) );
AND2x2_ASAP7_75t_L g569 ( .A(n_355), .B(n_567), .Y(n_569) );
BUFx2_ASAP7_75t_L g689 ( .A(n_355), .Y(n_689) );
INVx1_ASAP7_75t_L g378 ( .A(n_356), .Y(n_378) );
NAND2x1_ASAP7_75t_L g392 ( .A(n_357), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g396 ( .A(n_357), .B(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_SL g700 ( .A(n_357), .B(n_393), .Y(n_700) );
AND2x4_ASAP7_75t_SL g701 ( .A(n_357), .B(n_397), .Y(n_701) );
AND2x2_ASAP7_75t_L g852 ( .A(n_357), .B(n_393), .Y(n_852) );
AOI33xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_364), .A3(n_368), .B1(n_379), .B2(n_381), .B3(n_387), .Y(n_358) );
AOI33xp33_ASAP7_75t_L g858 ( .A1(n_359), .A2(n_859), .A3(n_862), .B1(n_864), .B2(n_866), .B3(n_868), .Y(n_858) );
AOI33xp33_ASAP7_75t_L g976 ( .A1(n_359), .A2(n_933), .A3(n_977), .B1(n_978), .B2(n_981), .B3(n_984), .Y(n_976) );
AOI33xp33_ASAP7_75t_L g1423 ( .A1(n_359), .A2(n_381), .A3(n_1424), .B1(n_1426), .B2(n_1427), .B3(n_1428), .Y(n_1423) );
NAND3xp33_ASAP7_75t_L g1542 ( .A(n_359), .B(n_1543), .C(n_1545), .Y(n_1542) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI33xp33_ASAP7_75t_L g687 ( .A1(n_360), .A2(n_688), .A3(n_690), .B1(n_693), .B2(n_695), .B3(n_697), .Y(n_687) );
AOI33xp33_ASAP7_75t_L g925 ( .A1(n_360), .A2(n_926), .A3(n_929), .B1(n_932), .B2(n_933), .B3(n_934), .Y(n_925) );
INVx1_ASAP7_75t_L g1028 ( .A(n_360), .Y(n_1028) );
AOI33xp33_ASAP7_75t_L g1137 ( .A1(n_360), .A2(n_1138), .A3(n_1139), .B1(n_1140), .B2(n_1141), .B3(n_1142), .Y(n_1137) );
AOI33xp33_ASAP7_75t_L g1159 ( .A1(n_360), .A2(n_933), .A3(n_1160), .B1(n_1161), .B2(n_1164), .B3(n_1165), .Y(n_1159) );
INVx3_ASAP7_75t_L g1513 ( .A(n_361), .Y(n_1513) );
INVx1_ASAP7_75t_L g589 ( .A(n_362), .Y(n_589) );
OAI31xp33_ASAP7_75t_SL g602 ( .A1(n_362), .A2(n_603), .A3(n_604), .B(n_608), .Y(n_602) );
OAI31xp33_ASAP7_75t_L g731 ( .A1(n_362), .A2(n_732), .A3(n_733), .B(n_753), .Y(n_731) );
INVx2_ASAP7_75t_SL g963 ( .A(n_362), .Y(n_963) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g458 ( .A(n_363), .Y(n_458) );
INVx8_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g471 ( .A(n_366), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_366), .Y(n_614) );
INVx3_ASAP7_75t_L g869 ( .A(n_366), .Y(n_869) );
INVx2_ASAP7_75t_L g1024 ( .A(n_366), .Y(n_1024) );
INVx1_ASAP7_75t_L g871 ( .A(n_367), .Y(n_871) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g473 ( .A(n_371), .B(n_472), .Y(n_473) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_371), .Y(n_979) );
INVx3_ASAP7_75t_L g1078 ( .A(n_371), .Y(n_1078) );
BUFx8_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g548 ( .A(n_372), .Y(n_548) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_372), .Y(n_557) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_372), .Y(n_692) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g863 ( .A(n_375), .Y(n_863) );
INVx5_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g380 ( .A(n_376), .Y(n_380) );
BUFx2_ASAP7_75t_L g549 ( .A(n_376), .Y(n_549) );
BUFx12f_ASAP7_75t_L g563 ( .A(n_376), .Y(n_563) );
AND2x4_ASAP7_75t_L g587 ( .A(n_376), .B(n_585), .Y(n_587) );
BUFx3_ASAP7_75t_L g980 ( .A(n_376), .Y(n_980) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx2_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g467 ( .A(n_377), .B(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g1514 ( .A(n_377), .Y(n_1514) );
INVx1_ASAP7_75t_L g399 ( .A(n_378), .Y(n_399) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g828 ( .A(n_383), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g1546 ( .A(n_383), .B(n_1547), .C(n_1549), .Y(n_1546) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g867 ( .A(n_384), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_395), .B2(n_396), .Y(n_389) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_390), .A2(n_395), .B1(n_435), .B2(n_437), .C1(n_439), .C2(n_450), .Y(n_434) );
AOI221x1_ASAP7_75t_L g818 ( .A1(n_391), .A2(n_396), .B1(n_792), .B2(n_798), .C(n_819), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_391), .A2(n_396), .B1(n_923), .B2(n_924), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_391), .A2(n_396), .B1(n_971), .B2(n_972), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_391), .A2(n_396), .B1(n_1066), .B2(n_1101), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_391), .A2(n_396), .B1(n_1155), .B2(n_1156), .Y(n_1154) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AO22x1_ASAP7_75t_L g850 ( .A1(n_396), .A2(n_851), .B1(n_852), .B2(n_853), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_396), .A2(n_852), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_455), .B(n_459), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_415), .C(n_434), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_409), .B2(n_410), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_403), .A2(n_409), .B1(n_470), .B2(n_473), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_404), .A2(n_1441), .B1(n_1442), .B2(n_1443), .Y(n_1440) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_405), .A2(n_411), .B1(n_974), .B2(n_975), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g1032 ( .A1(n_405), .A2(n_411), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_405), .B(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_405), .A2(n_411), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g542 ( .A(n_406), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g880 ( .A(n_406), .Y(n_880) );
AND2x4_ASAP7_75t_L g411 ( .A(n_407), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g416 ( .A(n_407), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_407), .B(n_422), .Y(n_436) );
AND2x2_ASAP7_75t_L g593 ( .A(n_407), .B(n_412), .Y(n_593) );
AND2x2_ASAP7_75t_L g655 ( .A(n_407), .B(n_531), .Y(n_655) );
BUFx2_ASAP7_75t_L g682 ( .A(n_407), .Y(n_682) );
HB1xp67_ASAP7_75t_L g1493 ( .A(n_408), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_410), .A2(n_879), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_410), .A2(n_879), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_411), .A2(n_874), .B1(n_875), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_411), .A2(n_655), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
INVx1_ASAP7_75t_L g1444 ( .A(n_411), .Y(n_1444) );
INVx2_ASAP7_75t_L g447 ( .A(n_412), .Y(n_447) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_412), .Y(n_886) );
INVx1_ASAP7_75t_L g1064 ( .A(n_412), .Y(n_1064) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g425 ( .A(n_413), .Y(n_425) );
INVx2_ASAP7_75t_L g662 ( .A(n_413), .Y(n_662) );
AND2x4_ASAP7_75t_L g1492 ( .A(n_413), .B(n_1493), .Y(n_1492) );
NAND2xp5_ASAP7_75t_R g892 ( .A(n_416), .B(n_856), .Y(n_892) );
INVx2_ASAP7_75t_SL g955 ( .A(n_416), .Y(n_955) );
INVx3_ASAP7_75t_L g1120 ( .A(n_416), .Y(n_1120) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_417), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g432 ( .A(n_418), .Y(n_432) );
INVx2_ASAP7_75t_L g532 ( .A(n_418), .Y(n_532) );
BUFx3_ASAP7_75t_L g659 ( .A(n_418), .Y(n_659) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g628 ( .A(n_422), .Y(n_628) );
BUFx3_ASAP7_75t_L g950 ( .A(n_422), .Y(n_950) );
INVx1_ASAP7_75t_L g991 ( .A(n_422), .Y(n_991) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_422), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_422), .B(n_1488), .Y(n_1487) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
BUFx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g1054 ( .A(n_425), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_425), .Y(n_1123) );
INVx4_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g637 ( .A(n_427), .B(n_638), .Y(n_637) );
INVx4_ASAP7_75t_L g668 ( .A(n_427), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g803 ( .A(n_427), .B(n_804), .C(n_805), .D(n_807), .Y(n_803) );
INVx1_ASAP7_75t_SL g887 ( .A(n_427), .Y(n_887) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g438 ( .A(n_430), .Y(n_438) );
INVx2_ASAP7_75t_L g665 ( .A(n_430), .Y(n_665) );
INVx1_ASAP7_75t_L g806 ( .A(n_430), .Y(n_806) );
INVx2_ASAP7_75t_L g889 ( .A(n_430), .Y(n_889) );
INVx1_ASAP7_75t_L g958 ( .A(n_430), .Y(n_958) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g891 ( .A(n_432), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_433), .A2(n_882), .B(n_888), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_433), .A2(n_957), .B(n_959), .Y(n_956) );
AOI21xp5_ASAP7_75t_SL g988 ( .A1(n_433), .A2(n_989), .B(n_994), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1035 ( .A1(n_433), .A2(n_655), .B1(n_1016), .B2(n_1036), .C(n_1038), .Y(n_1035) );
INVx1_ASAP7_75t_L g1058 ( .A(n_433), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_433), .A2(n_1122), .B(n_1124), .Y(n_1121) );
AOI21xp5_ASAP7_75t_L g1176 ( .A1(n_433), .A2(n_1177), .B(n_1178), .Y(n_1176) );
AOI21xp5_ASAP7_75t_L g1435 ( .A1(n_433), .A2(n_1436), .B(n_1439), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_435), .B(n_792), .Y(n_791) );
AOI222xp33_ASAP7_75t_L g1039 ( .A1(n_435), .A2(n_452), .B1(n_1020), .B2(n_1021), .C1(n_1040), .C2(n_1041), .Y(n_1039) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g896 ( .A(n_436), .Y(n_896) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g884 ( .A(n_443), .Y(n_884) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g952 ( .A(n_447), .Y(n_952) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g663 ( .A(n_449), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_449), .A2(n_501), .B1(n_898), .B2(n_899), .C(n_902), .Y(n_897) );
INVx2_ASAP7_75t_L g953 ( .A(n_449), .Y(n_953) );
INVx2_ASAP7_75t_L g1065 ( .A(n_449), .Y(n_1065) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_452), .A2(n_1061), .B1(n_1062), .B2(n_1066), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_452), .B(n_1114), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_453), .A2(n_676), .B1(n_677), .B2(n_679), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_453), .A2(n_677), .B1(n_798), .B2(n_799), .Y(n_797) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
INVx1_ASAP7_75t_L g913 ( .A(n_454), .Y(n_913) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_454), .B(n_1471), .Y(n_1485) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_455), .A2(n_877), .B(n_893), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_455), .A2(n_1031), .B(n_1042), .Y(n_1030) );
OAI21xp5_ASAP7_75t_L g1049 ( .A1(n_455), .A2(n_1050), .B(n_1059), .Y(n_1049) );
OAI21xp5_ASAP7_75t_SL g1111 ( .A1(n_455), .A2(n_1112), .B(n_1119), .Y(n_1111) );
OAI21xp5_ASAP7_75t_L g1174 ( .A1(n_455), .A2(n_1175), .B(n_1183), .Y(n_1174) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_457), .B(n_587), .Y(n_784) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g521 ( .A(n_458), .B(n_522), .Y(n_521) );
OR2x6_ASAP7_75t_L g698 ( .A(n_458), .B(n_551), .Y(n_698) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_458), .B(n_551), .Y(n_1025) );
INVx2_ASAP7_75t_L g1073 ( .A(n_460), .Y(n_1073) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
INVx2_ASAP7_75t_SL g643 ( .A(n_461), .Y(n_643) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_461), .B(n_465), .Y(n_1043) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g712 ( .A(n_465), .Y(n_712) );
INVx3_ASAP7_75t_L g622 ( .A(n_466), .Y(n_622) );
INVx4_ASAP7_75t_L g1088 ( .A(n_466), .Y(n_1088) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g580 ( .A(n_467), .Y(n_580) );
BUFx2_ASAP7_75t_L g1517 ( .A(n_468), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_470), .A2(n_473), .B1(n_874), .B2(n_875), .Y(n_873) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x4_ASAP7_75t_L g713 ( .A(n_471), .B(n_472), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_471), .A2(n_696), .B1(n_729), .B2(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g937 ( .A(n_473), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_473), .A2(n_713), .B1(n_974), .B2(n_975), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_473), .B(n_1068), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
AO22x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_917), .B1(n_1005), .B2(n_1006), .Y(n_477) );
XOR2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_647), .Y(n_478) );
XNOR2x1_ASAP7_75t_L g1006 ( .A(n_479), .B(n_647), .Y(n_1006) );
BUFx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
XNOR2x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_595), .Y(n_481) );
XNOR2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_594), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_544), .Y(n_483) );
NAND3xp33_ASAP7_75t_SL g484 ( .A(n_485), .B(n_523), .C(n_538), .Y(n_484) );
AOI211xp5_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_496), .B(n_506), .C(n_515), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g999 ( .A1(n_488), .A2(n_494), .B1(n_1000), .B2(n_1001), .C(n_1002), .Y(n_999) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g632 ( .A(n_490), .Y(n_632) );
INVx4_ASAP7_75t_L g802 ( .A(n_490), .Y(n_802) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_490), .Y(n_909) );
INVx1_ASAP7_75t_L g1448 ( .A(n_490), .Y(n_1448) );
INVx8_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g517 ( .A(n_491), .Y(n_517) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_491), .B(n_1471), .Y(n_1476) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_495), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
OAI22x1_ASAP7_75t_SL g635 ( .A1(n_495), .A2(n_612), .B1(n_632), .B2(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_498), .A2(n_501), .B1(n_519), .B2(n_520), .C(n_521), .Y(n_518) );
BUFx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g773 ( .A(n_499), .Y(n_773) );
BUFx2_ASAP7_75t_L g801 ( .A(n_499), .Y(n_801) );
BUFx2_ASAP7_75t_L g901 ( .A(n_499), .Y(n_901) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
BUFx4f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x6_ASAP7_75t_L g513 ( .A(n_502), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g674 ( .A(n_502), .Y(n_674) );
BUFx4f_ASAP7_75t_L g684 ( .A(n_502), .Y(n_684) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g536 ( .A(n_503), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_504), .A2(n_513), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g642 ( .A(n_507), .Y(n_642) );
INVx2_ASAP7_75t_SL g767 ( .A(n_507), .Y(n_767) );
NAND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g514 ( .A(n_508), .Y(n_514) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_SL g765 ( .A(n_512), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_513), .Y(n_646) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_521), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_521), .B(n_762), .Y(n_761) );
INVx4_ASAP7_75t_L g1534 ( .A(n_521), .Y(n_1534) );
AOI222xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_527), .B1(n_528), .B2(n_533), .C1(n_534), .C2(n_537), .Y(n_523) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_524), .A2(n_645), .B(n_646), .Y(n_644) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g640 ( .A1(n_528), .A2(n_606), .B1(n_618), .B2(n_641), .C1(n_642), .C2(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g780 ( .A(n_528), .Y(n_780) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g535 ( .A(n_530), .B(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g769 ( .A(n_530), .B(n_536), .Y(n_769) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g995 ( .A(n_532), .Y(n_995) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_533), .A2(n_571), .B(n_574), .C(n_582), .Y(n_570) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_534), .A2(n_607), .B1(n_627), .B2(n_633), .C1(n_634), .C2(n_637), .Y(n_626) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g811 ( .A(n_536), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_541), .B(n_837), .Y(n_836) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_542), .A2(n_592), .B1(n_729), .B2(n_730), .Y(n_728) );
AND2x4_ASAP7_75t_L g592 ( .A(n_543), .B(n_593), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_570), .B(n_588), .C(n_590), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_550), .B1(n_552), .B2(n_560), .C(n_564), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x6_ASAP7_75t_SL g583 ( .A(n_548), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g707 ( .A(n_548), .Y(n_707) );
BUFx2_ASAP7_75t_L g931 ( .A(n_548), .Y(n_931) );
BUFx2_ASAP7_75t_L g983 ( .A(n_548), .Y(n_983) );
INVx3_ASAP7_75t_L g616 ( .A(n_551), .Y(n_616) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g696 ( .A(n_554), .Y(n_696) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_556), .A2(n_610), .B1(n_611), .B2(n_612), .C(n_613), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_556), .A2(n_580), .B1(n_742), .B2(n_743), .C(n_744), .Y(n_741) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g746 ( .A(n_557), .Y(n_746) );
INVx5_ASAP7_75t_L g830 ( .A(n_557), .Y(n_830) );
INVx2_ASAP7_75t_SL g1163 ( .A(n_557), .Y(n_1163) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g865 ( .A(n_563), .Y(n_865) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_566), .A2(n_569), .B1(n_598), .B2(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx4_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_576), .A2(n_578), .B1(n_606), .B2(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_579), .A2(n_734), .B1(n_741), .B2(n_745), .C(n_750), .Y(n_733) );
OR2x6_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g1097 ( .A(n_580), .Y(n_1097) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_585), .Y(n_757) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_588), .Y(n_814) );
INVx1_ASAP7_75t_L g1452 ( .A(n_588), .Y(n_1452) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI21x1_ASAP7_75t_L g652 ( .A1(n_589), .A2(n_653), .B(n_685), .Y(n_652) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_589), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_592), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g709 ( .A(n_592), .Y(n_709) );
AOI211x1_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_599), .C(n_625), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_617), .C(n_619), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_611), .A2(n_809), .B1(n_830), .B2(n_831), .C(n_832), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_611), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1089) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B(n_623), .C(n_624), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g750 ( .A1(n_621), .A2(n_751), .B(n_752), .Y(n_750) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g1507 ( .A(n_622), .Y(n_1507) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_640), .C(n_644), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g1535 ( .A(n_637), .B(n_1536), .C(n_1541), .Y(n_1535) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AO22x2_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_844), .B1(n_915), .B2(n_916), .Y(n_647) );
INVx1_ASAP7_75t_L g915 ( .A(n_648), .Y(n_915) );
XNOR2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_787), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_724), .B1(n_785), .B2(n_786), .Y(n_649) );
INVx1_ASAP7_75t_L g786 ( .A(n_650), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_717), .C(n_721), .Y(n_650) );
INVx1_ASAP7_75t_L g718 ( .A(n_652), .Y(n_718) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B1(n_664), .B2(n_666), .Y(n_656) );
INVx3_ASAP7_75t_L g1126 ( .A(n_658), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g1179 ( .A(n_658), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_658), .B(n_1471), .Y(n_1470) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g667 ( .A(n_662), .Y(n_667) );
INVx2_ASAP7_75t_L g993 ( .A(n_667), .Y(n_993) );
HB1xp67_ASAP7_75t_L g1537 ( .A(n_667), .Y(n_1537) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_680), .B1(n_682), .B2(n_683), .Y(n_669) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx4_ASAP7_75t_L g795 ( .A(n_672), .Y(n_795) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_672), .Y(n_906) );
OAI211xp5_ASAP7_75t_L g1184 ( .A1(n_673), .A2(n_1185), .B(n_1186), .C(n_1188), .Y(n_1184) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g796 ( .A(n_674), .Y(n_796) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI222xp33_ASAP7_75t_L g711 ( .A1(n_679), .A2(n_712), .B1(n_713), .B2(n_714), .C1(n_715), .C2(n_716), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_680), .A2(n_682), .B1(n_794), .B2(n_800), .Y(n_793) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2x1_ASAP7_75t_L g912 ( .A(n_681), .B(n_913), .Y(n_912) );
OAI211xp5_ASAP7_75t_L g1115 ( .A1(n_684), .A2(n_1116), .B(n_1117), .C(n_1118), .Y(n_1115) );
INVx1_ASAP7_75t_L g719 ( .A(n_686), .Y(n_719) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_699), .Y(n_686) );
HB1xp67_ASAP7_75t_L g1544 ( .A(n_689), .Y(n_1544) );
INVx2_ASAP7_75t_L g1091 ( .A(n_691), .Y(n_1091) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_692), .Y(n_694) );
AND2x4_ASAP7_75t_L g1500 ( .A(n_692), .B(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g1141 ( .A(n_698), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g1019 ( .A1(n_700), .A2(n_701), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_700), .A2(n_701), .B1(n_1114), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g723 ( .A(n_703), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .Y(n_703) );
NAND2x1_ASAP7_75t_L g704 ( .A(n_705), .B(n_709), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_706), .A2(n_713), .B1(n_1033), .B2(n_1034), .Y(n_1044) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVxp67_ASAP7_75t_L g840 ( .A(n_708), .Y(n_840) );
INVx1_ASAP7_75t_L g722 ( .A(n_711), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_712), .A2(n_715), .B1(n_799), .B2(n_817), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_720), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g785 ( .A(n_724), .Y(n_785) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_758), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_731), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B1(n_738), .B2(n_740), .Y(n_734) );
BUFx4f_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g839 ( .A(n_736), .Y(n_839) );
BUFx3_ASAP7_75t_L g1084 ( .A(n_736), .Y(n_1084) );
BUFx3_ASAP7_75t_L g1095 ( .A(n_736), .Y(n_1095) );
OR2x4_ASAP7_75t_L g1523 ( .A(n_736), .B(n_1501), .Y(n_1523) );
INVx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g748 ( .A(n_739), .Y(n_748) );
INVx3_ASAP7_75t_L g824 ( .A(n_739), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g771 ( .A1(n_742), .A2(n_772), .B(n_774), .C(n_775), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_746), .A2(n_823), .B1(n_824), .B2(n_825), .C(n_826), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_755), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_776), .C(n_781), .Y(n_758) );
NOR3xp33_ASAP7_75t_SL g759 ( .A(n_760), .B(n_768), .C(n_770), .Y(n_759) );
OAI21xp5_ASAP7_75t_SL g760 ( .A1(n_761), .A2(n_763), .B(n_764), .Y(n_760) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_814), .B(n_815), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .C(n_803), .D(n_808), .Y(n_790) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B(n_812), .C(n_813), .Y(n_808) );
INVx5_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI22xp5_ASAP7_75t_SL g819 ( .A1(n_820), .A2(n_822), .B1(n_828), .B2(n_829), .Y(n_819) );
BUFx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx8_ASAP7_75t_L g1082 ( .A(n_821), .Y(n_1082) );
INVx2_ASAP7_75t_SL g861 ( .A(n_827), .Y(n_861) );
INVx1_ASAP7_75t_L g928 ( .A(n_827), .Y(n_928) );
BUFx3_ASAP7_75t_L g985 ( .A(n_827), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
OR2x6_ASAP7_75t_L g837 ( .A(n_838), .B(n_840), .Y(n_837) );
OR2x2_ASAP7_75t_L g936 ( .A(n_838), .B(n_840), .Y(n_936) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_843), .B(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_843), .B(n_1069), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_843), .B(n_1158), .Y(n_1157) );
INVx2_ASAP7_75t_L g916 ( .A(n_844), .Y(n_916) );
XOR2x2_ASAP7_75t_L g844 ( .A(n_845), .B(n_914), .Y(n_844) );
NAND2xp5_ASAP7_75t_SL g845 ( .A(n_846), .B(n_876), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_858), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_854), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g854 ( .A(n_855), .B(n_857), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g1099 ( .A(n_857), .B(n_1100), .C(n_1102), .D(n_1103), .Y(n_1099) );
NAND4xp25_ASAP7_75t_SL g1153 ( .A(n_857), .B(n_1154), .C(n_1157), .D(n_1159), .Y(n_1153) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
BUFx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx2_ASAP7_75t_L g933 ( .A(n_867), .Y(n_933) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND3xp33_ASAP7_75t_SL g877 ( .A(n_878), .B(n_881), .C(n_892), .Y(n_877) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g1540 ( .A(n_884), .Y(n_1540) );
BUFx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g944 ( .A(n_895), .Y(n_944) );
INVx2_ASAP7_75t_L g998 ( .A(n_895), .Y(n_998) );
INVx4_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx4_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_905), .B1(n_907), .B2(n_908), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g946 ( .A1(n_905), .A2(n_908), .B1(n_947), .B2(n_948), .C(n_949), .Y(n_946) );
OAI221xp5_ASAP7_75t_L g1446 ( .A1(n_905), .A2(n_1447), .B1(n_1448), .B2(n_1449), .C(n_1450), .Y(n_1446) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx5_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx2_ASAP7_75t_L g945 ( .A(n_912), .Y(n_945) );
INVx1_ASAP7_75t_L g1005 ( .A(n_917), .Y(n_1005) );
XNOR2x1_ASAP7_75t_L g917 ( .A(n_918), .B(n_964), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_939), .C(n_942), .Y(n_919) );
NOR3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_935), .C(n_938), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .Y(n_921) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
NOR3xp33_ASAP7_75t_L g1418 ( .A(n_938), .B(n_1419), .C(n_1429), .Y(n_1418) );
OAI21xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_954), .B(n_963), .Y(n_942) );
AOI222xp33_ASAP7_75t_L g1478 ( .A1(n_950), .A2(n_1479), .B1(n_1480), .B2(n_1483), .C1(n_1484), .C2(n_1485), .Y(n_1478) );
BUFx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
AND3x1_ASAP7_75t_L g969 ( .A(n_970), .B(n_973), .C(n_976), .Y(n_969) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
OAI21xp5_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_997), .B(n_1004), .Y(n_986) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g1003 ( .A(n_991), .Y(n_1003) );
INVx1_ASAP7_75t_L g1055 ( .A(n_991), .Y(n_1055) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
XNOR2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1106), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1045), .B1(n_1046), .B2(n_1105), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1013), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1030), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1026), .B1(n_1027), .B2(n_1029), .Y(n_1022) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1035), .C(n_1039), .Y(n_1031) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1037), .Y(n_1438) );
INVxp67_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
NOR3xp33_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1099), .C(n_1104), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1072), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1056), .Y(n_1051) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1054), .Y(n_1187) );
NAND3xp33_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1067), .C(n_1070), .Y(n_1059) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_1064), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B(n_1075), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1171 ( .A1(n_1073), .A2(n_1172), .B(n_1173), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1076) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1078), .Y(n_1548) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1083) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B1(n_1096), .B2(n_1098), .Y(n_1093) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
XOR2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1146), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1110), .Y(n_1145) );
NAND3xp33_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1130), .C(n_1133), .Y(n_1110) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1137), .Y(n_1134) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
NAND2x1p5_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1168), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1166), .Y(n_1151) );
INVxp67_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
NOR2xp33_ASAP7_75t_SL g1189 ( .A(n_1153), .B(n_1190), .Y(n_1189) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1166), .B(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1174), .Y(n_1170) );
OAI221xp5_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1411), .B1(n_1415), .B2(n_1455), .C(n_1459), .Y(n_1192) );
AND3x1_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1340), .C(n_1376), .Y(n_1193) );
NOR3xp33_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1271), .C(n_1329), .Y(n_1194) );
OAI221xp5_ASAP7_75t_L g1195 ( .A1(n_1196), .A2(n_1198), .B1(n_1248), .B2(n_1261), .C(n_1264), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1223), .B1(n_1229), .B2(n_1238), .C(n_1242), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1214), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1199), .B(n_1289), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_1199), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1199), .B(n_1343), .Y(n_1342) );
OAI211xp5_ASAP7_75t_SL g1377 ( .A1(n_1199), .A2(n_1378), .B(n_1381), .C(n_1393), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1199), .B(n_1275), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1408 ( .A(n_1199), .B(n_1409), .Y(n_1408) );
INVx4_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx4_ASAP7_75t_L g1231 ( .A(n_1200), .Y(n_1231) );
NAND2xp5_ASAP7_75t_SL g1246 ( .A(n_1200), .B(n_1247), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1200), .B(n_1247), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1200), .B(n_1332), .Y(n_1331) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_1200), .B(n_1263), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1200), .B(n_1299), .Y(n_1386) );
AND2x4_ASAP7_75t_SL g1200 ( .A(n_1201), .B(n_1209), .Y(n_1200) );
AND2x4_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
AND2x6_ASAP7_75t_L g1207 ( .A(n_1203), .B(n_1208), .Y(n_1207) );
AND2x6_ASAP7_75t_L g1210 ( .A(n_1203), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1203), .B(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1203), .B(n_1213), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1203), .B(n_1204), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1203), .B(n_1213), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1206), .Y(n_1204) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1207), .Y(n_1254) );
OAI21xp5_ASAP7_75t_L g1552 ( .A1(n_1213), .A2(n_1553), .B(n_1554), .Y(n_1552) );
INVxp67_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1215), .B(n_1231), .Y(n_1374) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1220), .Y(n_1215) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1216), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1216), .B(n_1239), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1216), .B(n_1247), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1216), .B(n_1238), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1216), .B(n_1239), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1385 ( .A(n_1216), .B(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1216), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1219), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1220), .B(n_1244), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1220), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1220), .B(n_1297), .Y(n_1321) );
AOI222xp33_ASAP7_75t_L g1407 ( .A1(n_1220), .A2(n_1343), .B1(n_1349), .B2(n_1357), .C1(n_1408), .C2(n_1410), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1222), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1221), .B(n_1222), .Y(n_1247) );
OAI321xp33_ASAP7_75t_L g1329 ( .A1(n_1223), .A2(n_1330), .A3(n_1333), .B1(n_1334), .B2(n_1335), .C(n_1336), .Y(n_1329) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1224), .B(n_1258), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_1224), .B(n_1231), .Y(n_1363) );
NOR2xp33_ASAP7_75t_L g1366 ( .A(n_1224), .B(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1225), .B(n_1234), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_1225), .B(n_1235), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1225), .B(n_1266), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1225), .B(n_1276), .Y(n_1283) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1225), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1225), .B(n_1258), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1225), .B(n_1258), .Y(n_1388) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1226), .B(n_1276), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1228), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1232), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1230), .B(n_1262), .Y(n_1285) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_1230), .B(n_1290), .C(n_1293), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1230), .B(n_1234), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1230), .B(n_1233), .Y(n_1410) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1231), .B(n_1234), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1231), .B(n_1251), .Y(n_1323) );
NAND2x1_ASAP7_75t_L g1400 ( .A(n_1231), .B(n_1401), .Y(n_1400) );
NOR2xp33_ASAP7_75t_L g1242 ( .A(n_1232), .B(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1233), .B(n_1332), .Y(n_1335) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1234), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1234), .B(n_1266), .Y(n_1345) );
OAI31xp33_ASAP7_75t_L g1391 ( .A1(n_1234), .A2(n_1239), .A3(n_1284), .B(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1235), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1289 ( .A(n_1238), .B(n_1290), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1238), .B(n_1247), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1238), .B(n_1247), .Y(n_1372) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1239), .B(n_1245), .Y(n_1244) );
NAND2x1p5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1246), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1244), .B(n_1296), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1344 ( .A(n_1244), .B(n_1290), .Y(n_1344) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1244), .Y(n_1379) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1246), .Y(n_1308) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1247), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1247), .B(n_1396), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1247), .B(n_1303), .Y(n_1401) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1247), .B(n_1396), .Y(n_1409) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
NOR2xp33_ASAP7_75t_SL g1249 ( .A(n_1250), .B(n_1258), .Y(n_1249) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1250), .Y(n_1311) );
A2O1A1Ixp33_ASAP7_75t_L g1317 ( .A1(n_1250), .A2(n_1299), .B(n_1318), .C(n_1320), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1250), .B(n_1265), .Y(n_1398) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1253), .B1(n_1254), .B2(n_1255), .C(n_1256), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1414 ( .A(n_1257), .Y(n_1414) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1258), .Y(n_1262) );
INVx3_ASAP7_75t_L g1266 ( .A(n_1258), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1261), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1263), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1392 ( .A(n_1262), .B(n_1269), .C(n_1297), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1267), .Y(n_1264) );
NAND3xp33_ASAP7_75t_L g1389 ( .A(n_1265), .B(n_1297), .C(n_1390), .Y(n_1389) );
CKINVDCx14_ASAP7_75t_R g1265 ( .A(n_1266), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1266), .B(n_1275), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1266), .B(n_1328), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1266), .B(n_1349), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1270), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1298), .C(n_1313), .Y(n_1271) );
AOI21xp5_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1281), .B(n_1282), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1277), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1274), .B(n_1306), .Y(n_1305) );
O2A1O1Ixp33_ASAP7_75t_L g1370 ( .A1(n_1274), .A2(n_1371), .B(n_1373), .C(n_1375), .Y(n_1370) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1275), .B(n_1281), .Y(n_1291) );
OAI22xp5_ASAP7_75t_SL g1322 ( .A1(n_1275), .A2(n_1310), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
OAI221xp5_ASAP7_75t_L g1399 ( .A1(n_1275), .A2(n_1400), .B1(n_1402), .B2(n_1403), .C(n_1407), .Y(n_1399) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AOI222xp33_ASAP7_75t_L g1393 ( .A1(n_1277), .A2(n_1293), .B1(n_1321), .B2(n_1348), .C1(n_1394), .C2(n_1395), .Y(n_1393) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1280), .Y(n_1278) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1279), .Y(n_1316) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1280), .Y(n_1307) );
OAI211xp5_ASAP7_75t_SL g1346 ( .A1(n_1280), .A2(n_1347), .B(n_1350), .C(n_1352), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1280), .B(n_1290), .Y(n_1354) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1281), .Y(n_1375) );
OAI322xp33_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1284), .A3(n_1286), .B1(n_1287), .B2(n_1291), .C1(n_1292), .C2(n_1294), .Y(n_1282) );
CKINVDCx5p33_ASAP7_75t_R g1349 ( .A(n_1283), .Y(n_1349) );
CKINVDCx14_ASAP7_75t_R g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1286), .Y(n_1368) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1290), .B(n_1307), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1290), .B(n_1297), .Y(n_1332) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1297), .B(n_1316), .Y(n_1356) );
A2O1A1Ixp33_ASAP7_75t_R g1298 ( .A1(n_1299), .A2(n_1300), .B(n_1304), .C(n_1309), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1299), .B(n_1351), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1299), .B(n_1320), .Y(n_1364) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1299), .Y(n_1402) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
AOI21xp33_ASAP7_75t_SL g1341 ( .A1(n_1301), .A2(n_1342), .B(n_1345), .Y(n_1341) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1303), .B(n_1316), .Y(n_1315) );
AOI211xp5_ASAP7_75t_L g1381 ( .A1(n_1303), .A2(n_1382), .B(n_1383), .C(n_1391), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1303), .B(n_1308), .Y(n_1406) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1312), .Y(n_1310) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1311), .Y(n_1334) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1312), .Y(n_1394) );
AOI222xp33_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1317), .B1(n_1321), .B2(n_1322), .C1(n_1325), .C2(n_1326), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
OAI21xp5_ASAP7_75t_L g1336 ( .A1(n_1321), .A2(n_1337), .B(n_1339), .Y(n_1336) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1321), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1324), .B(n_1325), .Y(n_1351) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1325), .Y(n_1360) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_1328), .Y(n_1357) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1376 ( .A1(n_1333), .A2(n_1377), .B1(n_1397), .B2(n_1399), .Y(n_1376) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OAI31xp33_ASAP7_75t_L g1340 ( .A1(n_1334), .A2(n_1341), .A3(n_1346), .B(n_1358), .Y(n_1340) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
OAI221xp5_ASAP7_75t_L g1358 ( .A1(n_1344), .A2(n_1359), .B1(n_1362), .B2(n_1364), .C(n_1365), .Y(n_1358) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
OAI21xp33_ASAP7_75t_L g1352 ( .A1(n_1353), .A2(n_1355), .B(n_1357), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_1354), .B(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1361), .Y(n_1359) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1364), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1370), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1369), .Y(n_1367) );
CKINVDCx14_ASAP7_75t_R g1371 ( .A(n_1372), .Y(n_1371) );
INVxp67_ASAP7_75t_SL g1373 ( .A(n_1374), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1380), .Y(n_1378) );
OAI21xp33_ASAP7_75t_L g1383 ( .A1(n_1384), .A2(n_1387), .B(n_1389), .Y(n_1383) );
INVxp33_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
INVxp67_ASAP7_75t_SL g1403 ( .A(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
CKINVDCx20_ASAP7_75t_R g1411 ( .A(n_1412), .Y(n_1411) );
CKINVDCx20_ASAP7_75t_R g1412 ( .A(n_1413), .Y(n_1412) );
INVx4_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1416), .Y(n_1454) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
NAND3xp33_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1430), .C(n_1433), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1423), .Y(n_1419) );
OAI21xp5_ASAP7_75t_L g1433 ( .A1(n_1434), .A2(n_1445), .B(n_1451), .Y(n_1433) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
CKINVDCx5p33_ASAP7_75t_R g1455 ( .A(n_1456), .Y(n_1455) );
BUFx3_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
BUFx3_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
BUFx4f_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1466), .Y(n_1550) );
NAND3xp33_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1497), .C(n_1529), .Y(n_1466) );
OAI21xp5_ASAP7_75t_L g1467 ( .A1(n_1468), .A2(n_1489), .B(n_1494), .Y(n_1467) );
NAND3xp33_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1478), .C(n_1486), .Y(n_1468) );
AOI22xp5_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1472), .B1(n_1473), .B2(n_1477), .Y(n_1469) );
INVx2_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx2_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx2_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_1483), .A2(n_1484), .B1(n_1511), .B2(n_1515), .Y(n_1510) );
INVx3_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx3_ASAP7_75t_SL g1491 ( .A(n_1492), .Y(n_1491) );
BUFx2_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
OAI31xp33_ASAP7_75t_L g1497 ( .A1(n_1498), .A2(n_1506), .A3(n_1518), .B(n_1524), .Y(n_1497) );
INVxp67_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx2_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
CKINVDCx8_ASAP7_75t_R g1508 ( .A(n_1509), .Y(n_1508) );
BUFx3_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1514), .Y(n_1512) );
AND2x4_ASAP7_75t_L g1516 ( .A(n_1513), .B(n_1517), .Y(n_1516) );
BUFx6f_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx2_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx2_ASAP7_75t_SL g1520 ( .A(n_1521), .Y(n_1520) );
BUFx3_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
AND2x4_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1527), .Y(n_1524) );
INVx1_ASAP7_75t_SL g1525 ( .A(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
AND4x1_ASAP7_75t_L g1529 ( .A(n_1530), .B(n_1535), .C(n_1542), .D(n_1546), .Y(n_1529) );
NAND3xp33_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1532), .C(n_1533), .Y(n_1530) );
INVx2_ASAP7_75t_SL g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
endmodule