module fake_jpeg_9177_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_182;
wire n_19;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_25),
.B1(n_31),
.B2(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_67),
.B1(n_25),
.B2(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx11_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_50),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_32),
.CI(n_39),
.CON(n_88),
.SN(n_88)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_68),
.C(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_29),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g114 ( 
.A(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_71),
.B(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_17),
.B1(n_33),
.B2(n_26),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_59),
.B1(n_58),
.B2(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_33),
.B1(n_26),
.B2(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_61),
.B1(n_60),
.B2(n_56),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_89),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_39),
.B(n_28),
.C(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_19),
.Y(n_103)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_98),
.B1(n_69),
.B2(n_70),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_115),
.Y(n_121)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_119),
.B1(n_75),
.B2(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_104),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_83),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AND2x6_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_32),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_84),
.B(n_32),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_59),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_41),
.B(n_58),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_115),
.B(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_74),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_49),
.B1(n_54),
.B2(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_113),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_143),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_76),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_139),
.C(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_134),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_104),
.B1(n_112),
.B2(n_105),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_142),
.B(n_144),
.Y(n_158)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_109),
.B1(n_107),
.B2(n_98),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_84),
.C(n_89),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_92),
.B1(n_64),
.B2(n_20),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_119),
.B1(n_96),
.B2(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_83),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_147),
.A2(n_148),
.B1(n_138),
.B2(n_49),
.Y(n_192)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_141),
.B1(n_129),
.B2(n_94),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_117),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_121),
.B(n_105),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_161),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_135),
.B(n_143),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_99),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_170),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_117),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_101),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_182),
.C(n_184),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_129),
.B1(n_141),
.B2(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_173),
.B1(n_185),
.B2(n_150),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_141),
.B1(n_137),
.B2(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_122),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_169),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_138),
.B1(n_124),
.B2(n_121),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_194),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_161),
.B(n_158),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_80),
.B(n_109),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_146),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_154),
.B1(n_145),
.B2(n_152),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_87),
.B1(n_132),
.B2(n_73),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_206),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_165),
.C(n_151),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_209),
.C(n_191),
.Y(n_218)
);

NOR2x1_ASAP7_75t_R g205 ( 
.A(n_178),
.B(n_155),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_184),
.C(n_176),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_155),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_194),
.B1(n_193),
.B2(n_154),
.Y(n_224)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_154),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_212),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_170),
.C(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_172),
.B1(n_188),
.B2(n_187),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_179),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_221),
.C(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_185),
.C(n_176),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_234),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_224),
.A2(n_228),
.B1(n_231),
.B2(n_62),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_179),
.C(n_145),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_214),
.B1(n_203),
.B2(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_73),
.C(n_132),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_41),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_156),
.B1(n_87),
.B2(n_62),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_212),
.B1(n_210),
.B2(n_213),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_233),
.A2(n_201),
.B1(n_204),
.B2(n_216),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_156),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_24),
.B1(n_1),
.B2(n_3),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_215),
.B1(n_201),
.B2(n_85),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_233),
.B1(n_230),
.B2(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_62),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_246),
.C(n_250),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_23),
.B1(n_24),
.B2(n_2),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_11),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_41),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_52),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_10),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_23),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_226),
.C(n_246),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_248),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_229),
.B1(n_222),
.B2(n_234),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_236),
.B(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_10),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_85),
.B1(n_24),
.B2(n_23),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_24),
.B1(n_1),
.B2(n_3),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_10),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_267),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_268),
.B(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_269),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_9),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_8),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_15),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_252),
.C(n_259),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_277),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_257),
.C(n_4),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_251),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_258),
.B(n_260),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_6),
.B(n_7),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_256),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_283),
.C(n_285),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_270),
.B(n_252),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_12),
.C(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_6),
.B1(n_7),
.B2(n_13),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_288),
.B(n_291),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_286),
.B(n_6),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_290),
.A3(n_7),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_0),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_293),
.C(n_0),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_0),
.B(n_22),
.Y(n_296)
);


endmodule