module fake_netlist_1_5862_n_707 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_707);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_707;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_62), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_1), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_5), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_60), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_5), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_30), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_42), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_27), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_56), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_83), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_57), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_18), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_49), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_63), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_3), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_34), .Y(n_109) );
NOR2xp67_ASAP7_75t_L g110 ( .A(n_29), .B(n_21), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_80), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_3), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_50), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_24), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_31), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_59), .Y(n_120) );
NOR2xp67_ASAP7_75t_L g121 ( .A(n_43), .B(n_87), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_9), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_68), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_51), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_47), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_125), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_116), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_108), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_116), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_95), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_125), .Y(n_134) );
INVx5_ASAP7_75t_L g135 ( .A(n_116), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_92), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_94), .A2(n_0), .B1(n_2), .B2(n_4), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_94), .B(n_4), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_125), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_102), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_145), .B(n_107), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_126), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_132), .B(n_91), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_126), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_145), .B(n_93), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_138), .B(n_101), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_141), .B(n_113), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_141), .B(n_97), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_129), .B(n_106), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_144), .B(n_122), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
INVx2_ASAP7_75t_SL g162 ( .A(n_129), .Y(n_162) );
OAI22xp33_ASAP7_75t_L g163 ( .A1(n_131), .A2(n_124), .B1(n_96), .B2(n_106), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_133), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_133), .B(n_119), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_133), .B(n_98), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
INVx1_ASAP7_75t_SL g169 ( .A(n_134), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_142), .B(n_100), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_142), .B(n_103), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_139), .B(n_102), .Y(n_172) );
NAND2xp33_ASAP7_75t_SL g173 ( .A(n_140), .B(n_109), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_139), .B(n_119), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
INVxp67_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_139), .B(n_104), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_146), .A2(n_120), .B1(n_99), .B2(n_105), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_143), .B(n_112), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_169), .B(n_120), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_158), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_148), .B(n_123), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_159), .B(n_6), .Y(n_189) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_157), .B(n_143), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
AOI221xp5_ASAP7_75t_L g192 ( .A1(n_163), .A2(n_146), .B1(n_104), .B2(n_111), .C(n_114), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_181), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_156), .B(n_143), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_157), .A2(n_143), .B1(n_146), .B2(n_111), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_153), .B(n_114), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_181), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_155), .B(n_115), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_179), .B(n_115), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_135), .B(n_110), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_158), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_179), .B(n_167), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_165), .B(n_146), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_160), .B(n_135), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_160), .B(n_135), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_157), .A2(n_158), .B1(n_166), .B2(n_173), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_157), .B(n_135), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_158), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_151), .B(n_110), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
INVxp33_ASAP7_75t_L g214 ( .A(n_174), .Y(n_214) );
BUFx12f_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_157), .B(n_121), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_152), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_170), .B(n_121), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g220 ( .A1(n_158), .A2(n_136), .B1(n_130), .B2(n_128), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_171), .B(n_17), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_194), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_194), .Y(n_223) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_215), .B(n_166), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_218), .A2(n_174), .B(n_172), .C(n_162), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_184), .B(n_162), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_203), .A2(n_180), .B(n_177), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_215), .A2(n_166), .B1(n_168), .B2(n_149), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_189), .B(n_166), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_184), .B(n_149), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_218), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_215), .A2(n_166), .B1(n_168), .B2(n_149), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_191), .B(n_168), .Y(n_233) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_201), .A2(n_177), .B(n_175), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_195), .A2(n_166), .B(n_176), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_192), .A2(n_175), .B1(n_178), .B2(n_164), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_204), .A2(n_178), .B(n_164), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_182), .B(n_175), .Y(n_238) );
OR2x6_ASAP7_75t_SL g239 ( .A(n_189), .B(n_6), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_209), .A2(n_161), .B1(n_136), .B2(n_130), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_214), .B(n_7), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_184), .B(n_161), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_197), .A2(n_217), .B(n_190), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_212), .B(n_8), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_187), .B(n_9), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_200), .A2(n_136), .B(n_130), .C(n_128), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_202), .B(n_10), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_183), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_219), .A2(n_136), .B(n_130), .Y(n_250) );
OA22x2_ASAP7_75t_L g251 ( .A1(n_199), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_210), .A2(n_136), .B(n_130), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_225), .A2(n_221), .B(n_186), .C(n_211), .Y(n_253) );
CKINVDCx6p67_ASAP7_75t_R g254 ( .A(n_239), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_227), .A2(n_196), .B(n_207), .C(n_208), .Y(n_255) );
BUFx4f_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_222), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_233), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_234), .A2(n_198), .B(n_216), .Y(n_259) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_227), .A2(n_250), .A3(n_247), .B(n_252), .Y(n_260) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_250), .A2(n_198), .B(n_216), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_223), .B(n_202), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_241), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_229), .B(n_202), .Y(n_264) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_246), .B(n_220), .C(n_184), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_243), .A2(n_213), .B(n_206), .Y(n_267) );
OAI22x1_ASAP7_75t_L g268 ( .A1(n_245), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_206), .B(n_198), .C(n_193), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_231), .B(n_248), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_252), .A2(n_206), .B(n_183), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_257), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_257), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_266), .B(n_249), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_263), .B(n_238), .Y(n_275) );
INVx6_ASAP7_75t_L g276 ( .A(n_264), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_270), .B(n_248), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_258), .B(n_228), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_256), .B(n_251), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_256), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_254), .B(n_232), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_268), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_269), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_259), .A2(n_237), .B(n_240), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_262), .B(n_251), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_259), .A2(n_237), .B(n_235), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_264), .B(n_226), .Y(n_288) );
NOR2x1_ASAP7_75t_SL g289 ( .A(n_261), .B(n_184), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_264), .B(n_262), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_255), .B(n_224), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_271), .A2(n_226), .B(n_242), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_255), .B(n_236), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_273), .B(n_261), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_281), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_291), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_283), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_272), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_273), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_273), .B(n_268), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_291), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_274), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_293), .A2(n_271), .B(n_267), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_279), .B(n_254), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_275), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_292), .A2(n_253), .B(n_265), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_290), .B(n_260), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_285), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g328 ( .A(n_282), .B(n_127), .C(n_128), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_297), .Y(n_333) );
OR2x2_ASAP7_75t_SL g334 ( .A(n_318), .B(n_292), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_326), .B(n_290), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_326), .B(n_290), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_299), .A2(n_278), .B(n_277), .C(n_281), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_311), .B(n_290), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_311), .B(n_294), .Y(n_341) );
OR2x2_ASAP7_75t_SL g342 ( .A(n_318), .B(n_278), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_315), .B(n_294), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_284), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_303), .B(n_284), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_313), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_301), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_302), .B(n_295), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_312), .A2(n_288), .B1(n_281), .B2(n_276), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_302), .B(n_288), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
NOR2xp67_ASAP7_75t_L g359 ( .A(n_323), .B(n_280), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_308), .B(n_288), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_295), .Y(n_362) );
BUFx4f_ASAP7_75t_SL g363 ( .A(n_319), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_313), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_306), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_320), .B(n_260), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_320), .B(n_321), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_306), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_307), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_320), .B(n_260), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_319), .B(n_276), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_321), .B(n_260), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_296), .B(n_276), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_296), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_321), .B(n_293), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_313), .B(n_276), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_307), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_327), .B(n_276), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_307), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_309), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_313), .B(n_13), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_327), .B(n_14), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_309), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_314), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_317), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_309), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_310), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_310), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_317), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_359), .B(n_324), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_358), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_355), .B(n_357), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_355), .B(n_324), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_357), .B(n_310), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_388), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_348), .B(n_316), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_362), .B(n_330), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_341), .B(n_330), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_341), .B(n_330), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_348), .B(n_15), .Y(n_406) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_359), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_365), .B(n_314), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_362), .B(n_325), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_364), .B(n_325), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_364), .B(n_325), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_367), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_335), .B(n_128), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_360), .B(n_15), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_351), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_335), .B(n_128), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_353), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_338), .B(n_328), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_336), .B(n_127), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_353), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_354), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_367), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_354), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_331), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_331), .Y(n_427) );
NAND2x1p5_ASAP7_75t_SL g428 ( .A(n_350), .B(n_230), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_336), .B(n_127), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_337), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_344), .B(n_127), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_365), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_361), .B(n_20), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_345), .B(n_337), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_343), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_340), .B(n_253), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_375), .B(n_22), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_361), .B(n_23), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
OR2x6_ASAP7_75t_SL g440 ( .A(n_342), .B(n_25), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_373), .B(n_26), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_373), .B(n_28), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_340), .B(n_32), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_363), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_347), .B(n_33), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_371), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_366), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_371), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_345), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_383), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_385), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_347), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_381), .B(n_35), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_381), .B(n_36), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_370), .B(n_37), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_369), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_392), .B(n_38), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_388), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_392), .B(n_39), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_352), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_375), .B(n_40), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_375), .B(n_41), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_375), .B(n_44), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_389), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_374), .B(n_45), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_369), .Y(n_467) );
OR2x6_ASAP7_75t_SL g468 ( .A(n_342), .B(n_46), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_389), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_372), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_350), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_380), .B(n_48), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_380), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_382), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_390), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_386), .B(n_52), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_390), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_474), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_413), .B(n_391), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_394), .B(n_370), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_453), .B(n_391), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_432), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_397), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_398), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_395), .B(n_386), .Y(n_485) );
OAI22xp33_ASAP7_75t_SL g486 ( .A1(n_440), .A2(n_379), .B1(n_384), .B2(n_376), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_396), .B(n_339), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_401), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_414), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_452), .B(n_368), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_400), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_414), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_415), .A2(n_356), .B1(n_368), .B2(n_378), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_444), .B(n_334), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_461), .B(n_378), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_402), .B(n_333), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_396), .B(n_333), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_417), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_434), .B(n_332), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_399), .B(n_332), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_399), .B(n_387), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_419), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_422), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_415), .B(n_387), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_400), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_423), .B(n_387), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_418), .B(n_387), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_425), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_426), .B(n_427), .Y(n_510) );
OR2x6_ASAP7_75t_L g511 ( .A(n_407), .B(n_387), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_430), .B(n_334), .Y(n_512) );
A2O1A1O1Ixp25_ASAP7_75t_L g513 ( .A1(n_420), .A2(n_53), .B(n_54), .C(n_55), .D(n_58), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_471), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_435), .B(n_61), .Y(n_515) );
OR2x6_ASAP7_75t_L g516 ( .A(n_400), .B(n_205), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_439), .B(n_64), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_434), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_424), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_457), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_424), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_421), .B(n_65), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_421), .B(n_66), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_449), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_429), .B(n_67), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_404), .B(n_69), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_405), .B(n_71), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_409), .B(n_73), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_431), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_409), .B(n_74), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_406), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_410), .B(n_75), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_409), .B(n_77), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_410), .B(n_411), .Y(n_537) );
OAI21xp33_ASAP7_75t_SL g538 ( .A1(n_451), .A2(n_78), .B(n_79), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_451), .B(n_81), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_446), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_446), .B(n_82), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_448), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_451), .B(n_84), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_411), .B(n_85), .Y(n_544) );
BUFx2_ASAP7_75t_SL g545 ( .A(n_459), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_412), .B(n_88), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_459), .B(n_89), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_450), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_459), .B(n_90), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_450), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_412), .B(n_185), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_471), .B(n_185), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_465), .B(n_188), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_465), .B(n_475), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_441), .B(n_188), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_440), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_469), .B(n_188), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_475), .B(n_193), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_441), .B(n_205), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_458), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_477), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_403), .B(n_205), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g563 ( .A(n_556), .B(n_463), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_482), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_518), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_478), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_534), .B(n_403), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_483), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_485), .B(n_408), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_537), .B(n_477), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_506), .B(n_408), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_502), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_480), .B(n_456), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_493), .A2(n_468), .B1(n_456), .B2(n_437), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_488), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_537), .B(n_436), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_487), .B(n_393), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_503), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_490), .B(n_442), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_479), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_504), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_497), .B(n_442), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_509), .Y(n_585) );
XNOR2xp5_ASAP7_75t_L g586 ( .A(n_500), .B(n_454), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_495), .B(n_496), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_520), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_499), .B(n_464), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_521), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_525), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_538), .A2(n_420), .B(n_472), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_526), .Y(n_594) );
NOR2x1p5_ASAP7_75t_L g595 ( .A(n_512), .B(n_468), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_527), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_481), .B(n_464), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_554), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_501), .B(n_462), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_514), .B(n_463), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_481), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_489), .Y(n_602) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_492), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_505), .B(n_463), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
NAND2x1_ASAP7_75t_L g607 ( .A(n_511), .B(n_437), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_494), .A2(n_466), .B1(n_437), .B2(n_416), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_548), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_538), .A2(n_476), .B(n_472), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_491), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_550), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_540), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_486), .A2(n_466), .B1(n_428), .B2(n_445), .C(n_443), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_561), .B(n_476), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_508), .B(n_455), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_545), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_532), .B(n_455), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_552), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_551), .B(n_454), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_507), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_551), .B(n_428), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_486), .B(n_460), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_491), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_557), .Y(n_626) );
OAI21xp33_ASAP7_75t_SL g627 ( .A1(n_618), .A2(n_511), .B(n_560), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_603), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_565), .B(n_560), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_587), .B(n_535), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_624), .B(n_513), .C(n_535), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_588), .B(n_546), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_611), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_618), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_572), .B(n_546), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_568), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_625), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_564), .A2(n_544), .B1(n_515), .B2(n_517), .C(n_528), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_573), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g641 ( .A(n_615), .B(n_524), .C(n_523), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_624), .A2(n_563), .B(n_593), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_575), .A2(n_555), .B1(n_531), .B2(n_530), .C(n_529), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_593), .A2(n_531), .B1(n_549), .B2(n_547), .C1(n_543), .C2(n_539), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_576), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_578), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_625), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_583), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_563), .A2(n_536), .B1(n_533), .B2(n_552), .Y(n_650) );
INVx4_ASAP7_75t_L g651 ( .A(n_600), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_585), .Y(n_652) );
INVxp33_ASAP7_75t_L g653 ( .A(n_586), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_582), .B(n_562), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_607), .A2(n_516), .B(n_558), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_620), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_569), .B(n_516), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_566), .Y(n_658) );
AOI32xp33_ASAP7_75t_L g659 ( .A1(n_600), .A2(n_513), .A3(n_559), .B1(n_433), .B2(n_438), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_610), .B(n_541), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_622), .B(n_558), .Y(n_661) );
NOR4xp25_ASAP7_75t_L g662 ( .A(n_635), .B(n_592), .C(n_589), .D(n_594), .Y(n_662) );
AOI211x1_ASAP7_75t_SL g663 ( .A1(n_631), .A2(n_610), .B(n_623), .C(n_577), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_642), .A2(n_608), .B(n_619), .C(n_581), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_643), .B(n_621), .C(n_581), .D(n_626), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_628), .B(n_591), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_634), .B(n_596), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_637), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_635), .A2(n_567), .A3(n_570), .B1(n_574), .B2(n_597), .C1(n_590), .C2(n_584), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g670 ( .A(n_659), .B(n_595), .C(n_579), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_640), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_653), .A2(n_598), .B1(n_606), .B2(n_612), .C(n_609), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_632), .A2(n_614), .B1(n_571), .B2(n_616), .C(n_599), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_645), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_660), .A2(n_617), .A3(n_605), .B1(n_616), .B2(n_602), .C1(n_613), .C2(n_604), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_646), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_644), .A2(n_205), .B1(n_553), .B2(n_641), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_647), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_649), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_633), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_656), .A2(n_654), .B1(n_651), .B2(n_636), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_655), .A2(n_656), .B(n_658), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_639), .A2(n_638), .B(n_652), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_650), .B(n_638), .C(n_661), .D(n_629), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_630), .A2(n_653), .B1(n_642), .B2(n_632), .C(n_635), .Y(n_685) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_648), .A2(n_642), .B1(n_653), .B2(n_635), .C1(n_627), .C2(n_643), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_657), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_670), .B(n_683), .Y(n_688) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_682), .B(n_684), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_664), .B(n_669), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_666), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_681), .B(n_687), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_662), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_688), .B(n_663), .C(n_686), .D(n_685), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_689), .B(n_677), .C(n_672), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_692), .B(n_674), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_695), .B(n_690), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_696), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_697), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_698), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_693), .B1(n_691), .B2(n_694), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_700), .B(n_671), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_701), .A2(n_699), .B1(n_680), .B2(n_676), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_702), .B(n_667), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_704), .A2(n_679), .B(n_678), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_705), .B(n_665), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_675), .B(n_673), .C(n_668), .Y(n_707) );
endmodule