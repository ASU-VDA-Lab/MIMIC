module fake_ibex_1276_n_6652 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1079, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_1080, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_1081, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_1083, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_1082, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1078, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_1073, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_6652);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1079;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_1080;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_1081;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_1083;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_1082;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1078;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_1073;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_6652;

wire n_4557;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_6616;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_6602;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_3979;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5969;
wire n_5920;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_6185;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6483;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_5397;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_2982;
wire n_2634;
wire n_3124;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3988;
wire n_3406;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6461;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_4437;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_5319;
wire n_2260;
wire n_4724;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_6448;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5488;
wire n_3107;
wire n_5465;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6361;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_1832;
wire n_3718;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_4878;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_2463;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4924;
wire n_2238;
wire n_6398;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_6480;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_6498;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6590;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_3261;
wire n_5324;
wire n_6547;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_6643;
wire n_6569;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6548;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_5436;
wire n_4887;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_5152;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_1523;
wire n_1086;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5595;
wire n_5334;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_2555;
wire n_1587;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6573;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6189;
wire n_6167;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3896;
wire n_3533;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_4650;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4542;
wire n_4122;
wire n_5021;
wire n_2819;
wire n_5523;
wire n_5456;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_6632;
wire n_1589;
wire n_2717;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_5214;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1566;
wire n_1464;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_3331;
wire n_2999;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_3449;
wire n_2923;
wire n_2990;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5992;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5349;
wire n_5054;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_965),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_983),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_845),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_881),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1002),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_10),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_755),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_598),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_982),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_83),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_703),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_420),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_574),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_293),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_510),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1070),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_134),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_998),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_976),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_615),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_599),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1009),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1008),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_628),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_762),
.Y(n_1108)
);

BUFx10_ASAP7_75t_L g1109 ( 
.A(n_643),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_972),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_581),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_596),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_756),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_614),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_727),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_808),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_961),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_643),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_343),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_711),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_193),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_471),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_558),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_654),
.Y(n_1124)
);

BUFx10_ASAP7_75t_L g1125 ( 
.A(n_380),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_422),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_253),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_830),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_542),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_959),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_77),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_146),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_257),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_10),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_29),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_984),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_897),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_214),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_296),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_579),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_447),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_445),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_488),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_833),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_967),
.Y(n_1145)
);

CKINVDCx16_ASAP7_75t_R g1146 ( 
.A(n_708),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1078),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_475),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_258),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1067),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_72),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_308),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_911),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_821),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_955),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_104),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1011),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_227),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_569),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_872),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1046),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_853),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_975),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_40),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_962),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_61),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_993),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_960),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_703),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_607),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_483),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_649),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_861),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_332),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_366),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_274),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_389),
.Y(n_1177)
);

CKINVDCx16_ASAP7_75t_R g1178 ( 
.A(n_349),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_22),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_18),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1047),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_629),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_624),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1075),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_682),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_395),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_319),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_992),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_400),
.Y(n_1189)
);

CKINVDCx14_ASAP7_75t_R g1190 ( 
.A(n_619),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_939),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_620),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_476),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_790),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_740),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_98),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1082),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_275),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_895),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_132),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_93),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1032),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_316),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1055),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_505),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_952),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_805),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_38),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_691),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_620),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_536),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_461),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_967),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1041),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_636),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_975),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_863),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1036),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_37),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_869),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_221),
.Y(n_1221)
);

BUFx10_ASAP7_75t_L g1222 ( 
.A(n_184),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_618),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_709),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_115),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_417),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_985),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_210),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_419),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_456),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_49),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_456),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_980),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_974),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_483),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_877),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_388),
.Y(n_1237)
);

BUFx2_ASAP7_75t_SL g1238 ( 
.A(n_20),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_202),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_934),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_410),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_146),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_318),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_678),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_851),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1017),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_940),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_651),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_423),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1075),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_26),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_420),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_239),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1021),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_190),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_393),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1082),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_585),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_425),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_981),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_526),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_511),
.Y(n_1262)
);

BUFx8_ASAP7_75t_SL g1263 ( 
.A(n_105),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_896),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_921),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_827),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_565),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_573),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_75),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_200),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_568),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_264),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_570),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_484),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_390),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_515),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_989),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_402),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_435),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_992),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_969),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_975),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_986),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_704),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_482),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_503),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_771),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_692),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1073),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_466),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_880),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_921),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_852),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_194),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_898),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_842),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1004),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_631),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_165),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_966),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_628),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_5),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_798),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_605),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_963),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_210),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_794),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_326),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_260),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_845),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_721),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_638),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_944),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1076),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_921),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_760),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_718),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_672),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_17),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_22),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_602),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_401),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1010),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_714),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_857),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_701),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1052),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_623),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_899),
.Y(n_1329)
);

BUFx8_ASAP7_75t_SL g1330 ( 
.A(n_766),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_935),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_799),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_841),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_289),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_970),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_218),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1063),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_438),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_39),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_425),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1024),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_278),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_806),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_457),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_219),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_139),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_125),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_37),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_606),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_195),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_519),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_689),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_364),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_987),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_462),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_907),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1048),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_238),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_389),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_18),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_147),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_207),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_932),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1077),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_257),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_578),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_163),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_35),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_701),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_137),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1035),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_172),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_844),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_127),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_922),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_283),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_339),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_33),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_26),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_800),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_314),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_343),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1048),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_124),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_971),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_646),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_623),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_768),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_951),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_513),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_410),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_367),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_11),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_270),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_54),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_682),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_349),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_483),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_134),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_530),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_41),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_684),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_358),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_305),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_415),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1014),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1063),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_945),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_348),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1007),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_284),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1062),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_476),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_321),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_354),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_187),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_53),
.Y(n_1417)
);

CKINVDCx16_ASAP7_75t_R g1418 ( 
.A(n_1072),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_863),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_658),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_300),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_634),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_49),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_194),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_730),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_208),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_319),
.Y(n_1427)
);

CKINVDCx16_ASAP7_75t_R g1428 ( 
.A(n_889),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_92),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_147),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_741),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_631),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_148),
.Y(n_1433)
);

CKINVDCx16_ASAP7_75t_R g1434 ( 
.A(n_970),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1000),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_640),
.Y(n_1436)
);

BUFx5_ASAP7_75t_L g1437 ( 
.A(n_1006),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_991),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_125),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_924),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_711),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_450),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_25),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_387),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_542),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_878),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_885),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_325),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_976),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_145),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_836),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_206),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_259),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_430),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_324),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_292),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_104),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_411),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_680),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_372),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_654),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_248),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_409),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_557),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_848),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_905),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_188),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_419),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_588),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_330),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_252),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_475),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_564),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_268),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_86),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_624),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_943),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_900),
.Y(n_1478)
);

BUFx2_ASAP7_75t_SL g1479 ( 
.A(n_416),
.Y(n_1479)
);

BUFx10_ASAP7_75t_L g1480 ( 
.A(n_1053),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_228),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_997),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_685),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1061),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_978),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_14),
.Y(n_1486)
);

CKINVDCx16_ASAP7_75t_R g1487 ( 
.A(n_887),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_734),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_226),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1012),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_698),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_33),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_285),
.Y(n_1493)
);

CKINVDCx16_ASAP7_75t_R g1494 ( 
.A(n_671),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_847),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_502),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1005),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_728),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_130),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_15),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_754),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1034),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_551),
.Y(n_1503)
);

CKINVDCx16_ASAP7_75t_R g1504 ( 
.A(n_211),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_935),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_342),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1029),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_384),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_495),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_345),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_849),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_805),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_389),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_457),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_258),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_776),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_973),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_754),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_337),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_310),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_676),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_69),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_994),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_179),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_775),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_254),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_492),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_440),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_648),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_845),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_855),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_347),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_841),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_49),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_770),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_452),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_252),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_777),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_100),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_289),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_51),
.Y(n_1542)
);

BUFx10_ASAP7_75t_L g1543 ( 
.A(n_440),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_233),
.Y(n_1544)
);

BUFx10_ASAP7_75t_L g1545 ( 
.A(n_83),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_728),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_648),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_984),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_512),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_117),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_698),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_463),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_470),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_663),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_396),
.Y(n_1555)
);

BUFx10_ASAP7_75t_L g1556 ( 
.A(n_1076),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_645),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_867),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_412),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_30),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1001),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_964),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1008),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_265),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_977),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_433),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_355),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_827),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_64),
.Y(n_1569)
);

BUFx10_ASAP7_75t_L g1570 ( 
.A(n_938),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_117),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_94),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_827),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_22),
.Y(n_1574)
);

INVxp67_ASAP7_75t_R g1575 ( 
.A(n_1080),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_836),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_11),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_805),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_100),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_137),
.Y(n_1580)
);

BUFx5_ASAP7_75t_L g1581 ( 
.A(n_501),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_446),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_776),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_134),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_406),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_606),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1065),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_451),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_417),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_547),
.Y(n_1590)
);

CKINVDCx16_ASAP7_75t_R g1591 ( 
.A(n_309),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_990),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_997),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_449),
.Y(n_1594)
);

BUFx8_ASAP7_75t_SL g1595 ( 
.A(n_1052),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_191),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_76),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_350),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_949),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_74),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_102),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_622),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_995),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_647),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_493),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_831),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_726),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_324),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_468),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_782),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1047),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_214),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_51),
.Y(n_1613)
);

CKINVDCx16_ASAP7_75t_R g1614 ( 
.A(n_881),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_530),
.Y(n_1615)
);

BUFx5_ASAP7_75t_L g1616 ( 
.A(n_703),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_542),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_865),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_338),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_883),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_868),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_813),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_379),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_588),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_987),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_622),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_661),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_613),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_340),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_722),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_183),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1027),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_691),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_475),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_412),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_997),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_12),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_395),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1003),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_257),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_634),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_318),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_510),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_540),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1013),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_527),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_378),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_935),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_492),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1015),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_604),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_260),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_400),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_684),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_194),
.Y(n_1655)
);

BUFx10_ASAP7_75t_L g1656 ( 
.A(n_430),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_988),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_806),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_994),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_303),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_78),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_714),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_99),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1079),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_968),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_530),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_262),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_270),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_55),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_368),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_521),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_117),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_410),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1064),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_613),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1025),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_390),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_682),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_294),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_841),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_980),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_946),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_742),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_999),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_109),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_31),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_341),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_527),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_738),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_289),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_447),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_631),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_294),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_158),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_200),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_996),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_90),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_979),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_851),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1004),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_438),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_754),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_916),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1050),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_580),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_188),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1062),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_559),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_799),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_889),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_455),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_285),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_423),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_85),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_208),
.Y(n_1715)
);

BUFx10_ASAP7_75t_L g1716 ( 
.A(n_878),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_700),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_847),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_68),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_920),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1073),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_161),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_733),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_266),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_521),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_826),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_740),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_248),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_663),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1728),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1728),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_1263),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1728),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1190),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1190),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1437),
.Y(n_1736)
);

CKINVDCx16_ASAP7_75t_R g1737 ( 
.A(n_1095),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1243),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1263),
.Y(n_1739)
);

INVxp67_ASAP7_75t_SL g1740 ( 
.A(n_1243),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1330),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1108),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1243),
.Y(n_1743)
);

CKINVDCx16_ASAP7_75t_R g1744 ( 
.A(n_1118),
.Y(n_1744)
);

CKINVDCx16_ASAP7_75t_R g1745 ( 
.A(n_1133),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1378),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1330),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1378),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1378),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1595),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1402),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1282),
.Y(n_1752)
);

CKINVDCx16_ASAP7_75t_R g1753 ( 
.A(n_1146),
.Y(n_1753)
);

INVxp33_ASAP7_75t_L g1754 ( 
.A(n_1094),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1595),
.Y(n_1755)
);

CKINVDCx20_ASAP7_75t_R g1756 ( 
.A(n_1087),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1402),
.Y(n_1757)
);

CKINVDCx16_ASAP7_75t_R g1758 ( 
.A(n_1178),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1402),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1307),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1398),
.Y(n_1761)
);

INVxp33_ASAP7_75t_L g1762 ( 
.A(n_1113),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1525),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1437),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1261),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1617),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1637),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1698),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1705),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1437),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1276),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1168),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1168),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_1087),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1368),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1428),
.Y(n_1776)
);

CKINVDCx16_ASAP7_75t_R g1777 ( 
.A(n_1434),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1109),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1368),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1487),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1391),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1391),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1104),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1421),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1421),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1494),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1457),
.Y(n_1787)
);

CKINVDCx16_ASAP7_75t_R g1788 ( 
.A(n_1504),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1457),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1523),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1523),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1684),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1684),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1101),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1103),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1105),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1650),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1110),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1707),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1104),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1480),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1591),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1162),
.Y(n_1803)
);

CKINVDCx16_ASAP7_75t_R g1804 ( 
.A(n_1614),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1162),
.Y(n_1805)
);

BUFx2_ASAP7_75t_SL g1806 ( 
.A(n_1109),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1121),
.Y(n_1807)
);

CKINVDCx20_ASAP7_75t_R g1808 ( 
.A(n_1120),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1437),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1129),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1131),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1437),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1437),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1136),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1137),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1480),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1143),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1120),
.Y(n_1818)
);

CKINVDCx20_ASAP7_75t_R g1819 ( 
.A(n_1175),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1145),
.Y(n_1820)
);

CKINVDCx20_ASAP7_75t_R g1821 ( 
.A(n_1175),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1720),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1148),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1196),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1084),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1169),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1151),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1085),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1086),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1171),
.Y(n_1830)
);

INVxp67_ASAP7_75t_SL g1831 ( 
.A(n_1196),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1153),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1155),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1160),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1320),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1166),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1320),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1514),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1172),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1089),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1180),
.Y(n_1841)
);

CKINVDCx16_ASAP7_75t_R g1842 ( 
.A(n_1109),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1182),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1090),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1183),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1185),
.Y(n_1846)
);

INVxp33_ASAP7_75t_SL g1847 ( 
.A(n_1575),
.Y(n_1847)
);

CKINVDCx14_ASAP7_75t_R g1848 ( 
.A(n_1125),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1188),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1192),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1437),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_1187),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1193),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1201),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1209),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1091),
.Y(n_1856)
);

INVxp67_ASAP7_75t_SL g1857 ( 
.A(n_1326),
.Y(n_1857)
);

INVxp33_ASAP7_75t_SL g1858 ( 
.A(n_1092),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1581),
.Y(n_1859)
);

CKINVDCx20_ASAP7_75t_R g1860 ( 
.A(n_1187),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1540),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1210),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1326),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_1384),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1212),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1581),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1219),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1220),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1799),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1736),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1764),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1734),
.B(n_1707),
.Y(n_1872)
);

OA21x2_ASAP7_75t_L g1873 ( 
.A1(n_1770),
.A2(n_1119),
.B(n_1111),
.Y(n_1873)
);

INVx4_ASAP7_75t_L g1874 ( 
.A(n_1842),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1730),
.A2(n_1119),
.B(n_1111),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1809),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1735),
.B(n_1093),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1812),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1813),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1778),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1848),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1786),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1851),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1740),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1742),
.A2(n_1232),
.B1(n_1288),
.B2(n_1227),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1778),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1859),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1866),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1740),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1749),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1742),
.B(n_1384),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1731),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1733),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1772),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1752),
.B(n_1474),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1754),
.Y(n_1896)
);

AND2x6_ASAP7_75t_L g1897 ( 
.A(n_1771),
.B(n_1474),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1824),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1773),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1775),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1738),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1746),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1748),
.Y(n_1903)
);

BUFx8_ASAP7_75t_L g1904 ( 
.A(n_1797),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1751),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1749),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1779),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1835),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1762),
.B(n_1125),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1765),
.B(n_1125),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1752),
.B(n_1511),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1835),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1825),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1765),
.A2(n_1232),
.B1(n_1288),
.B2(n_1227),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1757),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1759),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1781),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1782),
.Y(n_1918)
);

BUFx8_ASAP7_75t_L g1919 ( 
.A(n_1760),
.Y(n_1919)
);

OA21x2_ASAP7_75t_L g1920 ( 
.A1(n_1794),
.A2(n_1127),
.B(n_1124),
.Y(n_1920)
);

INVx4_ASAP7_75t_L g1921 ( 
.A(n_1828),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1822),
.B(n_1163),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1801),
.B(n_1511),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1803),
.B(n_1805),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1784),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1785),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1756),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1847),
.A2(n_1441),
.B1(n_1470),
.B2(n_1310),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1803),
.B(n_1096),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1837),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1816),
.B(n_1694),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1787),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1761),
.B(n_1694),
.Y(n_1933)
);

BUFx8_ASAP7_75t_L g1934 ( 
.A(n_1763),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1837),
.Y(n_1935)
);

NAND2xp33_ASAP7_75t_L g1936 ( 
.A(n_1795),
.B(n_1581),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1826),
.B(n_1163),
.Y(n_1937)
);

OA21x2_ASAP7_75t_L g1938 ( 
.A1(n_1796),
.A2(n_1127),
.B(n_1124),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1766),
.B(n_1181),
.Y(n_1939)
);

CKINVDCx6p67_ASAP7_75t_R g1940 ( 
.A(n_1737),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1857),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1805),
.B(n_1097),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1789),
.Y(n_1943)
);

BUFx8_ASAP7_75t_L g1944 ( 
.A(n_1767),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1830),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1790),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1791),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1829),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1792),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1743),
.B(n_1098),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1793),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1858),
.B(n_1246),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1857),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1798),
.Y(n_1954)
);

INVx5_ASAP7_75t_L g1955 ( 
.A(n_1806),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1863),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1838),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1863),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1807),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1840),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1831),
.B(n_1102),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1810),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1768),
.B(n_1418),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1811),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1864),
.Y(n_1965)
);

NAND2xp33_ASAP7_75t_L g1966 ( 
.A(n_1814),
.B(n_1581),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1815),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1861),
.A2(n_1441),
.B1(n_1470),
.B2(n_1310),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1769),
.B(n_1181),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1844),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1856),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1864),
.B(n_1106),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1817),
.B(n_1820),
.Y(n_1973)
);

CKINVDCx16_ASAP7_75t_R g1974 ( 
.A(n_1744),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1823),
.B(n_1107),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1827),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1832),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1833),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1745),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1834),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1753),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1776),
.Y(n_1982)
);

OA21x2_ASAP7_75t_L g1983 ( 
.A1(n_1836),
.A2(n_1200),
.B(n_1191),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1839),
.B(n_1112),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1841),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1843),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1845),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1846),
.B(n_1849),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_SL g1989 ( 
.A(n_1758),
.B(n_1163),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1850),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1739),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1853),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1854),
.B(n_1114),
.Y(n_1993)
);

INVx4_ASAP7_75t_L g1994 ( 
.A(n_1777),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1788),
.A2(n_1116),
.B1(n_1117),
.B2(n_1115),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1855),
.Y(n_1996)
);

NOR2x1_ASAP7_75t_L g1997 ( 
.A(n_1862),
.B(n_1221),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1865),
.B(n_1867),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1868),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1780),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1802),
.B(n_1099),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1804),
.B(n_1222),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1741),
.B(n_1147),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1747),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1750),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1755),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1732),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1774),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1783),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1860),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1800),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1808),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1818),
.B(n_1122),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1852),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1819),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1821),
.B(n_1150),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1799),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1799),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1734),
.B(n_1123),
.Y(n_2019)
);

OAI21x1_ASAP7_75t_L g2020 ( 
.A1(n_1730),
.A2(n_1200),
.B(n_1191),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1740),
.Y(n_2021)
);

XNOR2xp5_ASAP7_75t_L g2022 ( 
.A(n_1756),
.B(n_1475),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1740),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1740),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1799),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1740),
.Y(n_2026)
);

CKINVDCx6p67_ASAP7_75t_R g2027 ( 
.A(n_1842),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1799),
.Y(n_2028)
);

INVx4_ASAP7_75t_L g2029 ( 
.A(n_1842),
.Y(n_2029)
);

BUFx12f_ASAP7_75t_L g2030 ( 
.A(n_1739),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1734),
.B(n_1161),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1799),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1786),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1799),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1740),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1740),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1740),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1740),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1799),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1799),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1799),
.Y(n_2041)
);

CKINVDCx8_ASAP7_75t_R g2042 ( 
.A(n_1842),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1740),
.Y(n_2043)
);

AND2x6_ASAP7_75t_L g2044 ( 
.A(n_1778),
.B(n_1088),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1799),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1740),
.Y(n_2046)
);

BUFx12f_ASAP7_75t_L g2047 ( 
.A(n_1739),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1740),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1842),
.B(n_1581),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1799),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1799),
.Y(n_2051)
);

AND2x6_ASAP7_75t_L g2052 ( 
.A(n_1778),
.B(n_1088),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1740),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1734),
.B(n_1126),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1778),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1799),
.Y(n_2056)
);

OAI21x1_ASAP7_75t_L g2057 ( 
.A1(n_1730),
.A2(n_1273),
.B(n_1251),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1848),
.Y(n_2058)
);

OA21x2_ASAP7_75t_L g2059 ( 
.A1(n_1736),
.A2(n_1273),
.B(n_1251),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1734),
.B(n_1128),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1799),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1734),
.B(n_1130),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1740),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1799),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1824),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1734),
.B(n_1218),
.Y(n_2066)
);

AND2x6_ASAP7_75t_L g2067 ( 
.A(n_1778),
.B(n_1088),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1742),
.A2(n_1477),
.B1(n_1478),
.B2(n_1475),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_1778),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1799),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1754),
.B(n_1222),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1754),
.B(n_1222),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_1734),
.B(n_1257),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1734),
.B(n_1327),
.Y(n_2074)
);

INVx5_ASAP7_75t_L g2075 ( 
.A(n_1778),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1740),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1848),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1778),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1799),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1799),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_1734),
.B(n_1502),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_1778),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_SL g2083 ( 
.A1(n_1756),
.A2(n_1478),
.B1(n_1529),
.B2(n_1477),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1742),
.A2(n_1539),
.B1(n_1559),
.B2(n_1529),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1740),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1740),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1740),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1799),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1740),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1742),
.A2(n_1559),
.B1(n_1576),
.B2(n_1539),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1848),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1754),
.B(n_1374),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1734),
.B(n_1132),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1734),
.B(n_1134),
.Y(n_2094)
);

INVx2_ASAP7_75t_SL g2095 ( 
.A(n_1896),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_2032),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1875),
.Y(n_2097)
);

INVxp33_ASAP7_75t_L g2098 ( 
.A(n_1909),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1917),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2020),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2057),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1920),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1925),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1909),
.B(n_1374),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1920),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1938),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1938),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1983),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1983),
.Y(n_2109)
);

AOI21x1_ASAP7_75t_L g2110 ( 
.A1(n_1873),
.A2(n_1230),
.B(n_1226),
.Y(n_2110)
);

INVxp67_ASAP7_75t_L g2111 ( 
.A(n_1882),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1918),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1918),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_2071),
.Y(n_2114)
);

INVxp33_ASAP7_75t_L g2115 ( 
.A(n_2071),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1873),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1947),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1947),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1915),
.Y(n_2119)
);

INVx4_ASAP7_75t_L g2120 ( 
.A(n_1955),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2059),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1915),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_2072),
.B(n_1374),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2059),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1962),
.Y(n_2125)
);

NAND2xp33_ASAP7_75t_L g2126 ( 
.A(n_1897),
.B(n_1581),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_2044),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1962),
.Y(n_2128)
);

CKINVDCx6p67_ASAP7_75t_R g2129 ( 
.A(n_2027),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1964),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_SL g2131 ( 
.A(n_1989),
.B(n_1576),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1964),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1986),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1986),
.Y(n_2134)
);

INVxp67_ASAP7_75t_SL g2135 ( 
.A(n_1945),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1926),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1932),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_2072),
.B(n_1377),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1943),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1880),
.B(n_1135),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_2092),
.B(n_1377),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2092),
.B(n_1377),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1949),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1951),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1957),
.B(n_1448),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1910),
.B(n_1448),
.Y(n_2146)
);

AOI21x1_ASAP7_75t_L g2147 ( 
.A1(n_1916),
.A2(n_1236),
.B(n_1235),
.Y(n_2147)
);

NAND2xp33_ASAP7_75t_L g2148 ( 
.A(n_1897),
.B(n_1581),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1910),
.B(n_1448),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1924),
.B(n_1616),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1869),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_2044),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1894),
.Y(n_2153)
);

BUFx6f_ASAP7_75t_L g2154 ( 
.A(n_2044),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2017),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_1922),
.B(n_1937),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2018),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1899),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1922),
.A2(n_1139),
.B1(n_1140),
.B2(n_1138),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2025),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2028),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1900),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2039),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1937),
.B(n_1450),
.Y(n_2164)
);

NAND3xp33_ASAP7_75t_L g2165 ( 
.A(n_1952),
.B(n_1142),
.C(n_1141),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1955),
.B(n_1450),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1907),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1940),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2040),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1955),
.B(n_1450),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2041),
.Y(n_2171)
);

INVx8_ASAP7_75t_L g2172 ( 
.A(n_1897),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_2055),
.B(n_1144),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_2052),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1946),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2056),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_2069),
.B(n_1149),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1959),
.B(n_1616),
.Y(n_2178)
);

AO21x2_ASAP7_75t_L g2179 ( 
.A1(n_1936),
.A2(n_1245),
.B(n_1239),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2061),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1976),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2064),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2079),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2088),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_2065),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1892),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_2075),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1893),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1901),
.Y(n_2189)
);

NAND3xp33_ASAP7_75t_L g2190 ( 
.A(n_1995),
.B(n_1154),
.C(n_1152),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1902),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1891),
.B(n_1483),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1930),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1903),
.Y(n_2194)
);

BUFx6f_ASAP7_75t_L g2195 ( 
.A(n_2052),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_2077),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1905),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1930),
.Y(n_2198)
);

NOR2x1p5_ASAP7_75t_L g2199 ( 
.A(n_1874),
.B(n_1156),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1916),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1954),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1884),
.Y(n_2202)
);

CKINVDCx20_ASAP7_75t_R g2203 ( 
.A(n_1927),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1889),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1890),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1967),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1895),
.B(n_1483),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1980),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1906),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_2032),
.Y(n_2210)
);

INVx2_ASAP7_75t_SL g2211 ( 
.A(n_2091),
.Y(n_2211)
);

INVxp67_ASAP7_75t_SL g2212 ( 
.A(n_2033),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1985),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_SL g2214 ( 
.A(n_2029),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2021),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_2052),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1987),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_SL g2218 ( 
.A(n_1994),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1929),
.B(n_1616),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2023),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2024),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1911),
.B(n_1483),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2026),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1942),
.B(n_1616),
.Y(n_2224)
);

AND2x6_ASAP7_75t_L g2225 ( 
.A(n_2002),
.B(n_1284),
.Y(n_2225)
);

CKINVDCx6p67_ASAP7_75t_R g2226 ( 
.A(n_2030),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1972),
.B(n_1616),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_2067),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2035),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2036),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_2075),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2037),
.Y(n_2232)
);

AOI21x1_ASAP7_75t_L g2233 ( 
.A1(n_1870),
.A2(n_1258),
.B(n_1247),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2038),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1992),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1996),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_2075),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1961),
.B(n_1616),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1871),
.Y(n_2239)
);

AOI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_1963),
.A2(n_1158),
.B1(n_1159),
.B2(n_1157),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1871),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_2078),
.B(n_1164),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_2034),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2043),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2031),
.B(n_1543),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2046),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1888),
.Y(n_2247)
);

NOR2x1p5_ASAP7_75t_L g2248 ( 
.A(n_1881),
.B(n_1165),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2066),
.B(n_2073),
.Y(n_2249)
);

AND3x2_ASAP7_75t_L g2250 ( 
.A(n_1981),
.B(n_1585),
.C(n_1577),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2002),
.B(n_1543),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1888),
.Y(n_2252)
);

BUFx6f_ASAP7_75t_L g2253 ( 
.A(n_2067),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1950),
.B(n_2048),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2053),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_2082),
.B(n_1886),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2063),
.Y(n_2257)
);

AND3x2_ASAP7_75t_L g2258 ( 
.A(n_1981),
.B(n_1585),
.C(n_1577),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2076),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2085),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1948),
.B(n_1543),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2074),
.B(n_1545),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2086),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_1923),
.B(n_1344),
.Y(n_2264)
);

INVx2_ASAP7_75t_SL g2265 ( 
.A(n_1898),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2087),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2089),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2081),
.B(n_1545),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1908),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_1877),
.B(n_1167),
.Y(n_2270)
);

INVx2_ASAP7_75t_SL g2271 ( 
.A(n_1898),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1912),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_1975),
.B(n_1545),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1935),
.Y(n_2274)
);

OR2x2_ASAP7_75t_L g2275 ( 
.A(n_1974),
.B(n_1215),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_2058),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1941),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1953),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1956),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1958),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1965),
.B(n_1616),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1984),
.B(n_1170),
.Y(n_2282)
);

INVx8_ASAP7_75t_L g2283 ( 
.A(n_1931),
.Y(n_2283)
);

BUFx8_ASAP7_75t_SL g2284 ( 
.A(n_2047),
.Y(n_2284)
);

INVx2_ASAP7_75t_SL g2285 ( 
.A(n_1970),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1988),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1977),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1978),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1990),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1948),
.B(n_1570),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_1921),
.B(n_1570),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_1993),
.B(n_1570),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1999),
.Y(n_2293)
);

AND3x2_ASAP7_75t_L g2294 ( 
.A(n_1979),
.B(n_1631),
.C(n_1618),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1933),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2034),
.Y(n_2296)
);

INVx3_ASAP7_75t_L g2297 ( 
.A(n_2045),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2045),
.Y(n_2298)
);

AO21x2_ASAP7_75t_L g2299 ( 
.A1(n_1966),
.A2(n_1275),
.B(n_1265),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2050),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2050),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1997),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_2051),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1939),
.Y(n_2304)
);

INVxp67_ASAP7_75t_SL g2305 ( 
.A(n_1971),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1969),
.Y(n_2306)
);

INVx3_ASAP7_75t_L g2307 ( 
.A(n_2051),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2070),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_2019),
.B(n_1173),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2070),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2080),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2080),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1973),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1998),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1876),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2054),
.B(n_1656),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2060),
.B(n_1656),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1878),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1879),
.Y(n_2319)
);

INVx2_ASAP7_75t_SL g2320 ( 
.A(n_1872),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2062),
.B(n_1174),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1883),
.Y(n_2322)
);

AOI21x1_ASAP7_75t_L g2323 ( 
.A1(n_1887),
.A2(n_1293),
.B(n_1280),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2067),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2093),
.B(n_1176),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2049),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2094),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_2000),
.B(n_1656),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2001),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2003),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1913),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1960),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2016),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_1982),
.B(n_1177),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2042),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_1914),
.B(n_1716),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_1885),
.B(n_1716),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2004),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2005),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1991),
.B(n_1716),
.Y(n_2340)
);

CKINVDCx6p67_ASAP7_75t_R g2341 ( 
.A(n_2007),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2006),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_2013),
.B(n_1284),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2068),
.B(n_1480),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2084),
.B(n_1179),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2090),
.B(n_1556),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1904),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2008),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1968),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_L g2350 ( 
.A(n_1928),
.B(n_1189),
.C(n_1186),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1919),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_1934),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2015),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2022),
.B(n_1556),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1944),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2009),
.Y(n_2356)
);

AND2x6_ASAP7_75t_L g2357 ( 
.A(n_2007),
.B(n_1295),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2014),
.B(n_1195),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2083),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2022),
.B(n_1556),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2011),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2012),
.B(n_1198),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2011),
.Y(n_2363)
);

CKINVDCx20_ASAP7_75t_R g2364 ( 
.A(n_2010),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_1952),
.B(n_1203),
.C(n_1199),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1917),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1924),
.B(n_1205),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1924),
.B(n_1206),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1875),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1875),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1875),
.Y(n_2371)
);

AOI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_1910),
.A2(n_1208),
.B1(n_1211),
.B2(n_1207),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1917),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1917),
.Y(n_2374)
);

NAND2xp33_ASAP7_75t_L g2375 ( 
.A(n_1897),
.B(n_1088),
.Y(n_2375)
);

INVxp33_ASAP7_75t_L g2376 ( 
.A(n_1896),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1875),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1875),
.Y(n_2378)
);

INVx1_ASAP7_75t_SL g2379 ( 
.A(n_1896),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_1909),
.B(n_1295),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1875),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_1909),
.B(n_1335),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1917),
.Y(n_2383)
);

NAND2xp33_ASAP7_75t_SL g2384 ( 
.A(n_2077),
.B(n_1213),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1917),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1875),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1875),
.Y(n_2387)
);

INVx4_ASAP7_75t_L g2388 ( 
.A(n_1955),
.Y(n_2388)
);

AO21x2_ASAP7_75t_L g2389 ( 
.A1(n_1875),
.A2(n_1302),
.B(n_1300),
.Y(n_2389)
);

BUFx3_ASAP7_75t_L g2390 ( 
.A(n_2032),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_1875),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_1920),
.Y(n_2392)
);

INVx2_ASAP7_75t_SL g2393 ( 
.A(n_1896),
.Y(n_2393)
);

INVx2_ASAP7_75t_SL g2394 ( 
.A(n_1896),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_1875),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_1896),
.B(n_1216),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_1880),
.B(n_1217),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1875),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1875),
.Y(n_2399)
);

CKINVDCx6p67_ASAP7_75t_R g2400 ( 
.A(n_2027),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1920),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2200),
.Y(n_2402)
);

OAI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2116),
.A2(n_1306),
.B(n_1304),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2286),
.Y(n_2404)
);

INVx2_ASAP7_75t_SL g2405 ( 
.A(n_2379),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2129),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2220),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2111),
.B(n_1618),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2220),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2102),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2327),
.B(n_1223),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2102),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2221),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2221),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2223),
.Y(n_2415)
);

XOR2x2_ASAP7_75t_L g2416 ( 
.A(n_2250),
.B(n_1631),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2102),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2223),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2229),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2229),
.Y(n_2420)
);

OAI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2116),
.A2(n_1315),
.B(n_1312),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2327),
.B(n_1225),
.Y(n_2422)
);

OAI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2121),
.A2(n_1324),
.B(n_1319),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2104),
.B(n_1228),
.Y(n_2424)
);

XOR2xp5_ASAP7_75t_L g2425 ( 
.A(n_2203),
.B(n_1661),
.Y(n_2425)
);

XNOR2x2_ASAP7_75t_L g2426 ( 
.A(n_2131),
.B(n_1342),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2095),
.B(n_1661),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2230),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2230),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2232),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2232),
.Y(n_2431)
);

XOR2xp5_ASAP7_75t_L g2432 ( 
.A(n_2168),
.B(n_1710),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2400),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2393),
.B(n_1710),
.Y(n_2434)
);

INVx2_ASAP7_75t_SL g2435 ( 
.A(n_2394),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_2226),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_SL g2437 ( 
.A(n_2335),
.B(n_1711),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2098),
.B(n_1711),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2234),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2234),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2396),
.B(n_1197),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2244),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2109),
.Y(n_2443)
);

XNOR2x2_ASAP7_75t_L g2444 ( 
.A(n_2350),
.B(n_1409),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2244),
.Y(n_2445)
);

XNOR2x2_ASAP7_75t_L g2446 ( 
.A(n_2354),
.B(n_1422),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2246),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2246),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2259),
.Y(n_2449)
);

OR2x2_ASAP7_75t_L g2450 ( 
.A(n_2275),
.B(n_2376),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2259),
.Y(n_2451)
);

XNOR2x2_ASAP7_75t_L g2452 ( 
.A(n_2360),
.B(n_1424),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2109),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2266),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2266),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2109),
.Y(n_2456)
);

CKINVDCx20_ASAP7_75t_R g2457 ( 
.A(n_2364),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2269),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2392),
.Y(n_2459)
);

CKINVDCx20_ASAP7_75t_R g2460 ( 
.A(n_2284),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_SL g2461 ( 
.A(n_2355),
.B(n_1197),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2269),
.Y(n_2462)
);

INVxp33_ASAP7_75t_L g2463 ( 
.A(n_2261),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2135),
.B(n_1357),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2212),
.B(n_1357),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2193),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2198),
.Y(n_2467)
);

INVxp33_ASAP7_75t_L g2468 ( 
.A(n_2290),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2251),
.B(n_1484),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2202),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2204),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2205),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2209),
.Y(n_2473)
);

INVx4_ASAP7_75t_L g2474 ( 
.A(n_2172),
.Y(n_2474)
);

OR2x6_ASAP7_75t_L g2475 ( 
.A(n_2347),
.B(n_1238),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2215),
.Y(n_2476)
);

OAI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2121),
.A2(n_1331),
.B(n_1329),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2257),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2115),
.B(n_1229),
.Y(n_2479)
);

INVx1_ASAP7_75t_SL g2480 ( 
.A(n_2196),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2274),
.Y(n_2481)
);

XNOR2xp5_ASAP7_75t_L g2482 ( 
.A(n_2258),
.B(n_1484),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2279),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2255),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_2156),
.B(n_1231),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2336),
.B(n_1676),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2142),
.B(n_1676),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2260),
.Y(n_2488)
);

OAI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2369),
.A2(n_2391),
.B(n_2370),
.Y(n_2489)
);

NAND2x1p5_ASAP7_75t_L g2490 ( 
.A(n_2285),
.B(n_1499),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2254),
.B(n_1233),
.Y(n_2491)
);

AND2x2_ASAP7_75t_SL g2492 ( 
.A(n_2352),
.B(n_1721),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_SL g2493 ( 
.A(n_2351),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2097),
.A2(n_1352),
.B(n_1335),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2263),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2267),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2114),
.B(n_1234),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2249),
.B(n_1237),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2272),
.Y(n_2499)
);

CKINVDCx5p33_ASAP7_75t_R g2500 ( 
.A(n_2214),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2127),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_L g2502 ( 
.A(n_2145),
.B(n_1240),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2277),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2164),
.B(n_2123),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2338),
.B(n_1651),
.Y(n_2505)
);

INVxp33_ASAP7_75t_L g2506 ( 
.A(n_2291),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2278),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2280),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2127),
.B(n_1241),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_2214),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2293),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2287),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2288),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2289),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2099),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2103),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2138),
.B(n_1242),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2136),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2313),
.B(n_1244),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2137),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2392),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2392),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2366),
.Y(n_2523)
);

INVxp67_ASAP7_75t_SL g2524 ( 
.A(n_2401),
.Y(n_2524)
);

AND2x6_ASAP7_75t_L g2525 ( 
.A(n_2105),
.B(n_1352),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2373),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2374),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2383),
.Y(n_2528)
);

INVxp33_ASAP7_75t_L g2529 ( 
.A(n_2362),
.Y(n_2529)
);

INVxp67_ASAP7_75t_L g2530 ( 
.A(n_2211),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2141),
.B(n_2342),
.Y(n_2531)
);

OR2x6_ASAP7_75t_L g2532 ( 
.A(n_2352),
.B(n_1479),
.Y(n_2532)
);

XNOR2x2_ASAP7_75t_L g2533 ( 
.A(n_2337),
.B(n_1558),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2385),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2139),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2342),
.B(n_1248),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2143),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2144),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_SL g2539 ( 
.A(n_2276),
.B(n_2218),
.Y(n_2539)
);

CKINVDCx20_ASAP7_75t_R g2540 ( 
.A(n_2341),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2305),
.B(n_1721),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2201),
.Y(n_2542)
);

AND2x6_ASAP7_75t_L g2543 ( 
.A(n_2106),
.B(n_2107),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2206),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2208),
.Y(n_2545)
);

CKINVDCx20_ASAP7_75t_R g2546 ( 
.A(n_2384),
.Y(n_2546)
);

XOR2xp5_ASAP7_75t_L g2547 ( 
.A(n_2159),
.B(n_1249),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2218),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2401),
.Y(n_2549)
);

INVxp33_ASAP7_75t_L g2550 ( 
.A(n_2344),
.Y(n_2550)
);

XOR2xp5_ASAP7_75t_L g2551 ( 
.A(n_2359),
.B(n_1252),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2372),
.B(n_1253),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2213),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2217),
.Y(n_2554)
);

CKINVDCx16_ASAP7_75t_R g2555 ( 
.A(n_2225),
.Y(n_2555)
);

XOR2xp5_ASAP7_75t_L g2556 ( 
.A(n_2359),
.B(n_1255),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2235),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2236),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2346),
.B(n_1256),
.Y(n_2559)
);

OR2x2_ASAP7_75t_SL g2560 ( 
.A(n_2349),
.B(n_1674),
.Y(n_2560)
);

XNOR2x2_ASAP7_75t_L g2561 ( 
.A(n_2240),
.B(n_1561),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2245),
.B(n_1259),
.Y(n_2562)
);

INVx2_ASAP7_75t_SL g2563 ( 
.A(n_2283),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2262),
.B(n_1260),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2186),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2188),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2189),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2191),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2338),
.B(n_1334),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2194),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2331),
.B(n_1339),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2197),
.Y(n_2572)
);

XOR2x2_ASAP7_75t_L g2573 ( 
.A(n_2294),
.B(n_0),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2281),
.Y(n_2574)
);

INVxp67_ASAP7_75t_SL g2575 ( 
.A(n_2401),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2380),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2185),
.B(n_1262),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2382),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2270),
.B(n_1264),
.Y(n_2579)
);

XOR2xp5_ASAP7_75t_L g2580 ( 
.A(n_2190),
.B(n_2165),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2181),
.Y(n_2581)
);

NOR2xp67_ASAP7_75t_L g2582 ( 
.A(n_2365),
.B(n_0),
.Y(n_2582)
);

CKINVDCx14_ASAP7_75t_R g2583 ( 
.A(n_2357),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2309),
.B(n_1266),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2178),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2153),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2325),
.B(n_1267),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2264),
.B(n_1268),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2268),
.B(n_1269),
.Y(n_2589)
);

INVx2_ASAP7_75t_SL g2590 ( 
.A(n_2283),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2162),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2225),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2264),
.B(n_1270),
.Y(n_2593)
);

INVxp33_ASAP7_75t_SL g2594 ( 
.A(n_2334),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2167),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_SL g2596 ( 
.A(n_2172),
.B(n_1271),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2175),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2322),
.Y(n_2598)
);

XNOR2x2_ASAP7_75t_L g2599 ( 
.A(n_2333),
.B(n_1566),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2345),
.B(n_1272),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2322),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2120),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2146),
.B(n_1274),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2108),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2158),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2149),
.B(n_1277),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2158),
.Y(n_2607)
);

NOR2xp67_ASAP7_75t_L g2608 ( 
.A(n_2329),
.B(n_0),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2304),
.Y(n_2609)
);

INVx2_ASAP7_75t_SL g2610 ( 
.A(n_2120),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2306),
.Y(n_2611)
);

AOI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2100),
.A2(n_1381),
.B(n_1365),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2332),
.B(n_1346),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2321),
.B(n_1278),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2329),
.B(n_1279),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2348),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2320),
.B(n_1281),
.Y(n_2617)
);

XOR2xp5_ASAP7_75t_L g2618 ( 
.A(n_2333),
.B(n_1283),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2339),
.B(n_1350),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2353),
.Y(n_2620)
);

CKINVDCx20_ASAP7_75t_R g2621 ( 
.A(n_2388),
.Y(n_2621)
);

OAI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2369),
.A2(n_1354),
.B(n_1351),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2151),
.Y(n_2623)
);

INVx1_ASAP7_75t_SL g2624 ( 
.A(n_2357),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2155),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2157),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2160),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2389),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2096),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2161),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2163),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2169),
.Y(n_2632)
);

INVx1_ASAP7_75t_SL g2633 ( 
.A(n_2357),
.Y(n_2633)
);

INVx2_ASAP7_75t_SL g2634 ( 
.A(n_2388),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2225),
.Y(n_2635)
);

XNOR2xp5_ASAP7_75t_L g2636 ( 
.A(n_2199),
.B(n_1285),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2171),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2176),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2180),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_SL g2640 ( 
.A(n_2225),
.B(n_1286),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2182),
.Y(n_2641)
);

INVxp33_ASAP7_75t_L g2642 ( 
.A(n_2330),
.Y(n_2642)
);

XNOR2x2_ASAP7_75t_L g2643 ( 
.A(n_2140),
.B(n_1612),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2183),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_SL g2645 ( 
.A(n_2127),
.B(n_1287),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2184),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2295),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2227),
.Y(n_2648)
);

BUFx8_ASAP7_75t_L g2649 ( 
.A(n_2357),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2238),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2101),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2328),
.B(n_1355),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2150),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2371),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2302),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2219),
.Y(n_2656)
);

CKINVDCx20_ASAP7_75t_R g2657 ( 
.A(n_2210),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2192),
.B(n_2207),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2367),
.B(n_1290),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2368),
.B(n_1291),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2224),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2233),
.Y(n_2662)
);

XNOR2x2_ASAP7_75t_L g2663 ( 
.A(n_2173),
.B(n_1647),
.Y(n_2663)
);

OR2x2_ASAP7_75t_L g2664 ( 
.A(n_2356),
.B(n_1702),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_2248),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2323),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2314),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2147),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2282),
.B(n_1292),
.Y(n_2669)
);

NOR2xp67_ASAP7_75t_L g2670 ( 
.A(n_2358),
.B(n_1),
.Y(n_2670)
);

AND2x6_ASAP7_75t_L g2671 ( 
.A(n_2152),
.B(n_1365),
.Y(n_2671)
);

INVxp33_ASAP7_75t_SL g2672 ( 
.A(n_2177),
.Y(n_2672)
);

INVxp33_ASAP7_75t_L g2673 ( 
.A(n_2361),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2315),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2318),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2242),
.B(n_1294),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2397),
.B(n_1296),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2319),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2187),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2187),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2231),
.Y(n_2681)
);

NAND2xp33_ASAP7_75t_SL g2682 ( 
.A(n_2152),
.B(n_2154),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2231),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2237),
.Y(n_2684)
);

NOR2xp67_ASAP7_75t_L g2685 ( 
.A(n_2340),
.B(n_1),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2237),
.Y(n_2686)
);

XOR2x2_ASAP7_75t_L g2687 ( 
.A(n_2222),
.B(n_2316),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2370),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2391),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2326),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2265),
.B(n_1297),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2256),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2166),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2170),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_L g2695 ( 
.A(n_2317),
.B(n_1298),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2124),
.Y(n_2696)
);

XNOR2xp5_ASAP7_75t_L g2697 ( 
.A(n_2343),
.B(n_2273),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2292),
.B(n_1299),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2271),
.B(n_1301),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2110),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2308),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2310),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2296),
.Y(n_2703)
);

CKINVDCx20_ASAP7_75t_R g2704 ( 
.A(n_2390),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2298),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2300),
.Y(n_2706)
);

XOR2xp5_ASAP7_75t_L g2707 ( 
.A(n_2363),
.B(n_1303),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2243),
.B(n_1305),
.Y(n_2708)
);

AND2x2_ASAP7_75t_SL g2709 ( 
.A(n_2126),
.B(n_1381),
.Y(n_2709)
);

OR2x2_ASAP7_75t_L g2710 ( 
.A(n_2243),
.B(n_1718),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2377),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2311),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2152),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_L g2714 ( 
.A(n_2297),
.B(n_1308),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2297),
.B(n_1309),
.Y(n_2715)
);

NAND2xp33_ASAP7_75t_SL g2716 ( 
.A(n_2154),
.B(n_1311),
.Y(n_2716)
);

XOR2xp5_ASAP7_75t_L g2717 ( 
.A(n_2154),
.B(n_1313),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2312),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2378),
.Y(n_2719)
);

BUFx6f_ASAP7_75t_L g2720 ( 
.A(n_2174),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2301),
.Y(n_2721)
);

BUFx2_ASAP7_75t_R g2722 ( 
.A(n_2179),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2301),
.B(n_1316),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2303),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2303),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_2307),
.B(n_1317),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2307),
.B(n_1318),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2174),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2299),
.B(n_1321),
.Y(n_2729)
);

INVxp33_ASAP7_75t_L g2730 ( 
.A(n_2112),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2381),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_L g2732 ( 
.A(n_2148),
.B(n_1322),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2113),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2117),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2386),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2118),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2125),
.B(n_1323),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2387),
.Y(n_2738)
);

INVxp67_ASAP7_75t_L g2739 ( 
.A(n_2375),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2395),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2398),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2174),
.Y(n_2742)
);

XOR2xp5_ASAP7_75t_L g2743 ( 
.A(n_2195),
.B(n_1325),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_L g2744 ( 
.A(n_2128),
.B(n_1328),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_2130),
.Y(n_2745)
);

XNOR2xp5_ASAP7_75t_L g2746 ( 
.A(n_2132),
.B(n_1332),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2195),
.B(n_1333),
.Y(n_2747)
);

NOR2xp67_ASAP7_75t_L g2748 ( 
.A(n_2133),
.B(n_1),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2399),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2134),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2119),
.B(n_1336),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2122),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2195),
.B(n_1338),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2324),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2216),
.B(n_1340),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2216),
.B(n_1343),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2324),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_SL g2758 ( 
.A(n_2216),
.B(n_1345),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2228),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2228),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2228),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2253),
.Y(n_2762)
);

INVx4_ASAP7_75t_SL g2763 ( 
.A(n_2253),
.Y(n_2763)
);

XOR2xp5_ASAP7_75t_L g2764 ( 
.A(n_2253),
.B(n_1347),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2239),
.Y(n_2765)
);

INVxp33_ASAP7_75t_L g2766 ( 
.A(n_2241),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2247),
.B(n_1348),
.Y(n_2767)
);

OAI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2252),
.A2(n_1369),
.B(n_1361),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2286),
.B(n_1379),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2286),
.Y(n_2770)
);

CKINVDCx20_ASAP7_75t_R g2771 ( 
.A(n_2129),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2098),
.B(n_1349),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2097),
.A2(n_1455),
.B(n_1393),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_SL g2774 ( 
.A(n_2131),
.B(n_1353),
.Y(n_2774)
);

CKINVDCx20_ASAP7_75t_R g2775 ( 
.A(n_2129),
.Y(n_2775)
);

OR2x2_ASAP7_75t_L g2776 ( 
.A(n_2379),
.B(n_1356),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2286),
.Y(n_2777)
);

OR2x6_ASAP7_75t_L g2778 ( 
.A(n_2347),
.B(n_1393),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2286),
.Y(n_2779)
);

CKINVDCx5p33_ASAP7_75t_R g2780 ( 
.A(n_2129),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2200),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2286),
.B(n_1358),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2098),
.B(n_1359),
.Y(n_2783)
);

INVxp67_ASAP7_75t_SL g2784 ( 
.A(n_2095),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2286),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2286),
.Y(n_2786)
);

XOR2x2_ASAP7_75t_L g2787 ( 
.A(n_2250),
.B(n_2),
.Y(n_2787)
);

AND2x2_ASAP7_75t_L g2788 ( 
.A(n_2379),
.B(n_1360),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2286),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2286),
.B(n_1362),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2404),
.B(n_2770),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2777),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2779),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2785),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2786),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2789),
.B(n_1363),
.Y(n_2796)
);

INVxp67_ASAP7_75t_SL g2797 ( 
.A(n_2405),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2738),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2769),
.B(n_1366),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2511),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2769),
.B(n_1367),
.Y(n_2801)
);

BUFx8_ASAP7_75t_L g2802 ( 
.A(n_2493),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2667),
.B(n_1370),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2550),
.B(n_1372),
.Y(n_2804)
);

BUFx2_ASAP7_75t_L g2805 ( 
.A(n_2457),
.Y(n_2805)
);

NOR3xp33_ASAP7_75t_SL g2806 ( 
.A(n_2665),
.B(n_1375),
.C(n_1373),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2470),
.Y(n_2807)
);

A2O1A1Ixp33_ASAP7_75t_L g2808 ( 
.A1(n_2653),
.A2(n_1488),
.B(n_1489),
.C(n_1455),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2471),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2491),
.B(n_1376),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2740),
.Y(n_2811)
);

INVx5_ASAP7_75t_L g2812 ( 
.A(n_2671),
.Y(n_2812)
);

NAND2x1p5_ASAP7_75t_L g2813 ( 
.A(n_2474),
.B(n_1100),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2407),
.B(n_1382),
.Y(n_2814)
);

INVx2_ASAP7_75t_SL g2815 ( 
.A(n_2540),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_SL g2816 ( 
.A(n_2480),
.B(n_1385),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2472),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2409),
.B(n_1386),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2594),
.B(n_1388),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2473),
.Y(n_2820)
);

AND2x6_ASAP7_75t_L g2821 ( 
.A(n_2624),
.B(n_1100),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_SL g2822 ( 
.A(n_2774),
.B(n_1392),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2413),
.B(n_1394),
.Y(n_2823)
);

INVxp67_ASAP7_75t_L g2824 ( 
.A(n_2437),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2414),
.B(n_1395),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2476),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2478),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2741),
.Y(n_2828)
);

OAI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2461),
.A2(n_1399),
.B1(n_1400),
.B2(n_1397),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2481),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2483),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2463),
.B(n_1401),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2489),
.A2(n_1389),
.B(n_1387),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2403),
.A2(n_1489),
.B1(n_1517),
.B2(n_1488),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2415),
.B(n_1405),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2640),
.B(n_1406),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2418),
.B(n_1408),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_SL g2838 ( 
.A(n_2555),
.B(n_1410),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2450),
.B(n_1411),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_SL g2840 ( 
.A(n_2435),
.B(n_1413),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2512),
.Y(n_2841)
);

INVx4_ASAP7_75t_L g2842 ( 
.A(n_2474),
.Y(n_2842)
);

INVx4_ASAP7_75t_L g2843 ( 
.A(n_2436),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2468),
.B(n_1417),
.Y(n_2844)
);

INVx2_ASAP7_75t_SL g2845 ( 
.A(n_2490),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2600),
.B(n_1420),
.Y(n_2846)
);

INVx5_ASAP7_75t_L g2847 ( 
.A(n_2671),
.Y(n_2847)
);

AOI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2700),
.A2(n_1549),
.B(n_1517),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2505),
.B(n_1423),
.Y(n_2849)
);

INVxp67_ASAP7_75t_L g2850 ( 
.A(n_2788),
.Y(n_2850)
);

AND2x6_ASAP7_75t_SL g2851 ( 
.A(n_2532),
.B(n_1390),
.Y(n_2851)
);

NOR3xp33_ASAP7_75t_L g2852 ( 
.A(n_2559),
.B(n_1250),
.C(n_1214),
.Y(n_2852)
);

O2A1O1Ixp33_ASAP7_75t_L g2853 ( 
.A1(n_2411),
.A2(n_1403),
.B(n_1404),
.C(n_1396),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2749),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2419),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2506),
.B(n_1425),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2408),
.B(n_1430),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2505),
.B(n_1431),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2659),
.B(n_1433),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2487),
.A2(n_1438),
.B1(n_1439),
.B2(n_1435),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2513),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2660),
.B(n_1440),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2541),
.B(n_1444),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2569),
.B(n_1445),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2569),
.B(n_1446),
.Y(n_2865)
);

INVx8_ASAP7_75t_L g2866 ( 
.A(n_2532),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2464),
.B(n_1449),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2614),
.B(n_1451),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2465),
.B(n_1454),
.Y(n_2869)
);

AOI22xp33_ASAP7_75t_L g2870 ( 
.A1(n_2486),
.A2(n_1462),
.B1(n_1463),
.B2(n_1459),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2469),
.B(n_1464),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_SL g2872 ( 
.A(n_2530),
.B(n_1465),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2422),
.B(n_1466),
.Y(n_2873)
);

INVx4_ASAP7_75t_L g2874 ( 
.A(n_2406),
.Y(n_2874)
);

OR2x6_ASAP7_75t_L g2875 ( 
.A(n_2475),
.B(n_1549),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2596),
.B(n_2645),
.Y(n_2876)
);

OAI221xp5_ASAP7_75t_L g2877 ( 
.A1(n_2438),
.A2(n_1469),
.B1(n_1471),
.B2(n_1468),
.C(n_1467),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2427),
.A2(n_1473),
.B1(n_1481),
.B2(n_1472),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2514),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_SL g2880 ( 
.A(n_2758),
.B(n_1485),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_2672),
.B(n_1486),
.Y(n_2881)
);

INVx2_ASAP7_75t_SL g2882 ( 
.A(n_2657),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2529),
.B(n_1490),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2420),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2579),
.B(n_1492),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2584),
.B(n_1495),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2587),
.B(n_1496),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_2425),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_2776),
.B(n_1497),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2784),
.B(n_1501),
.Y(n_2890)
);

AOI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2434),
.A2(n_1506),
.B1(n_1508),
.B2(n_1503),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2441),
.B(n_1509),
.Y(n_2892)
);

INVx2_ASAP7_75t_SL g2893 ( 
.A(n_2704),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2428),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2484),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2488),
.Y(n_2896)
);

AOI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2547),
.A2(n_1512),
.B1(n_1513),
.B2(n_1510),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2782),
.B(n_1516),
.Y(n_2898)
);

CKINVDCx5p33_ASAP7_75t_R g2899 ( 
.A(n_2771),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2429),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2688),
.A2(n_1415),
.B(n_1414),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2495),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2790),
.B(n_1518),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2664),
.B(n_1519),
.Y(n_2904)
);

INVx2_ASAP7_75t_SL g2905 ( 
.A(n_2475),
.Y(n_2905)
);

INVx2_ASAP7_75t_SL g2906 ( 
.A(n_2621),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_SL g2907 ( 
.A(n_2592),
.B(n_1521),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_2759),
.Y(n_2908)
);

BUFx3_ASAP7_75t_L g2909 ( 
.A(n_2775),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2466),
.B(n_2467),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2552),
.B(n_1522),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2430),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_SL g2913 ( 
.A(n_2635),
.B(n_1524),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2618),
.B(n_1526),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2431),
.B(n_1530),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2439),
.B(n_1531),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2496),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_L g2918 ( 
.A(n_2502),
.B(n_1533),
.Y(n_2918)
);

CKINVDCx5p33_ASAP7_75t_R g2919 ( 
.A(n_2460),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2689),
.A2(n_2654),
.B(n_2651),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2440),
.Y(n_2921)
);

AOI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2479),
.A2(n_1536),
.B1(n_1537),
.B2(n_1535),
.Y(n_2922)
);

O2A1O1Ixp5_ASAP7_75t_L g2923 ( 
.A1(n_2494),
.A2(n_1592),
.B(n_1672),
.C(n_1580),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2442),
.B(n_1538),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2577),
.B(n_1544),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2445),
.B(n_2447),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2499),
.Y(n_2927)
);

INVx2_ASAP7_75t_SL g2928 ( 
.A(n_2778),
.Y(n_2928)
);

BUFx5_ASAP7_75t_L g2929 ( 
.A(n_2543),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2424),
.B(n_1546),
.Y(n_2930)
);

NAND3xp33_ASAP7_75t_SL g2931 ( 
.A(n_2546),
.B(n_1552),
.C(n_1550),
.Y(n_2931)
);

INVx2_ASAP7_75t_SL g2932 ( 
.A(n_2778),
.Y(n_2932)
);

AOI22xp33_ASAP7_75t_L g2933 ( 
.A1(n_2533),
.A2(n_1554),
.B1(n_1557),
.B2(n_1553),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2448),
.B(n_1560),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2449),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2772),
.A2(n_1563),
.B1(n_1564),
.B2(n_1562),
.Y(n_2936)
);

INVx3_ASAP7_75t_L g2937 ( 
.A(n_2501),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2503),
.Y(n_2938)
);

INVx4_ASAP7_75t_L g2939 ( 
.A(n_2433),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2451),
.B(n_1565),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2492),
.B(n_1567),
.Y(n_2941)
);

INVx5_ASAP7_75t_L g2942 ( 
.A(n_2671),
.Y(n_2942)
);

NOR2x2_ASAP7_75t_L g2943 ( 
.A(n_2432),
.B(n_1580),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2454),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2446),
.A2(n_1571),
.B1(n_1572),
.B2(n_1569),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2560),
.B(n_1578),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2452),
.A2(n_2561),
.B1(n_2593),
.B2(n_2588),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_SL g2948 ( 
.A(n_2649),
.B(n_1579),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2507),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2497),
.B(n_1584),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2455),
.B(n_1589),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2458),
.B(n_2462),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2711),
.A2(n_1426),
.B(n_1419),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2649),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2619),
.B(n_1596),
.Y(n_2955)
);

INVx2_ASAP7_75t_SL g2956 ( 
.A(n_2500),
.Y(n_2956)
);

OAI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2668),
.A2(n_1429),
.B(n_1427),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2709),
.B(n_1601),
.Y(n_2958)
);

INVx2_ASAP7_75t_SL g2959 ( 
.A(n_2510),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2508),
.Y(n_2960)
);

O2A1O1Ixp33_ASAP7_75t_L g2961 ( 
.A1(n_2519),
.A2(n_1436),
.B(n_1442),
.C(n_1432),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2642),
.B(n_1602),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_SL g2963 ( 
.A(n_2783),
.B(n_1603),
.Y(n_2963)
);

NAND2x1p5_ASAP7_75t_L g2964 ( 
.A(n_2501),
.B(n_1100),
.Y(n_2964)
);

O2A1O1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2669),
.A2(n_1447),
.B(n_1452),
.C(n_1443),
.Y(n_2965)
);

AOI221xp5_ASAP7_75t_L g2966 ( 
.A1(n_2536),
.A2(n_1606),
.B1(n_1613),
.B2(n_1605),
.C(n_1604),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2619),
.B(n_1615),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2498),
.B(n_1619),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2571),
.B(n_1621),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2571),
.B(n_1622),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2515),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2613),
.B(n_1624),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2746),
.B(n_1625),
.Y(n_2973)
);

OR2x6_ASAP7_75t_L g2974 ( 
.A(n_2563),
.B(n_2590),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2696),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2516),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2562),
.B(n_1626),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2676),
.B(n_1627),
.Y(n_2978)
);

AND2x6_ASAP7_75t_L g2979 ( 
.A(n_2633),
.B(n_1100),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2622),
.B(n_2574),
.Y(n_2980)
);

AOI22xp33_ASAP7_75t_L g2981 ( 
.A1(n_2485),
.A2(n_1634),
.B1(n_1639),
.B2(n_1629),
.Y(n_2981)
);

INVx2_ASAP7_75t_SL g2982 ( 
.A(n_2548),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2518),
.Y(n_2983)
);

INVxp67_ASAP7_75t_SL g2984 ( 
.A(n_2717),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2539),
.B(n_1640),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2613),
.B(n_1643),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2564),
.B(n_1648),
.Y(n_2987)
);

INVx6_ASAP7_75t_L g2988 ( 
.A(n_2629),
.Y(n_2988)
);

AND2x6_ASAP7_75t_SL g2989 ( 
.A(n_2416),
.B(n_2482),
.Y(n_2989)
);

BUFx5_ASAP7_75t_L g2990 ( 
.A(n_2543),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2531),
.B(n_1649),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2691),
.B(n_1652),
.Y(n_2992)
);

OR2x2_ASAP7_75t_L g2993 ( 
.A(n_2743),
.B(n_1654),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2729),
.B(n_1655),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2589),
.B(n_1657),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2520),
.B(n_1660),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2604),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2719),
.Y(n_2998)
);

A2O1A1Ixp33_ASAP7_75t_L g2999 ( 
.A1(n_2648),
.A2(n_1672),
.B(n_1683),
.C(n_1592),
.Y(n_2999)
);

INVx2_ASAP7_75t_SL g3000 ( 
.A(n_2764),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2617),
.A2(n_1666),
.B1(n_1668),
.B2(n_1662),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_L g3002 ( 
.A1(n_2599),
.A2(n_1670),
.B1(n_1675),
.B2(n_1669),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2523),
.B(n_1677),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2526),
.B(n_1678),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2527),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2747),
.B(n_1680),
.Y(n_3006)
);

NAND3xp33_ASAP7_75t_L g3007 ( 
.A(n_2582),
.B(n_1224),
.C(n_1194),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2731),
.A2(n_1456),
.B(n_1453),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2697),
.B(n_1681),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2643),
.A2(n_1685),
.B1(n_1686),
.B2(n_1682),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2528),
.B(n_1687),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2534),
.B(n_1688),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_SL g3013 ( 
.A(n_2753),
.B(n_2755),
.Y(n_3013)
);

AND2x6_ASAP7_75t_SL g3014 ( 
.A(n_2780),
.B(n_1458),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2735),
.Y(n_3015)
);

INVx8_ASAP7_75t_L g3016 ( 
.A(n_2671),
.Y(n_3016)
);

INVxp67_ASAP7_75t_L g3017 ( 
.A(n_2710),
.Y(n_3017)
);

O2A1O1Ixp5_ASAP7_75t_L g3018 ( 
.A1(n_2612),
.A2(n_1683),
.B(n_1476),
.C(n_1482),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2609),
.B(n_1689),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2421),
.A2(n_1194),
.B1(n_1380),
.B2(n_1224),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_SL g3021 ( 
.A(n_2423),
.B(n_1690),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2699),
.B(n_1691),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2611),
.B(n_1693),
.Y(n_3023)
);

OR2x2_ASAP7_75t_L g3024 ( 
.A(n_2707),
.B(n_1695),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2692),
.B(n_2616),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2620),
.B(n_1696),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2652),
.B(n_1697),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2658),
.B(n_1700),
.Y(n_3028)
);

AND2x6_ASAP7_75t_SL g3029 ( 
.A(n_2787),
.B(n_1460),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2652),
.B(n_1703),
.Y(n_3030)
);

BUFx3_ASAP7_75t_L g3031 ( 
.A(n_2426),
.Y(n_3031)
);

AOI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2615),
.A2(n_1708),
.B1(n_1709),
.B2(n_1706),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2647),
.B(n_1712),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2504),
.B(n_1713),
.Y(n_3034)
);

INVx2_ASAP7_75t_SL g3035 ( 
.A(n_2708),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2517),
.B(n_1715),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2477),
.B(n_1717),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2576),
.B(n_1719),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2578),
.B(n_1722),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2677),
.B(n_1723),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2598),
.Y(n_3041)
);

BUFx3_ASAP7_75t_L g3042 ( 
.A(n_2602),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2580),
.B(n_2723),
.Y(n_3043)
);

A2O1A1Ixp33_ASAP7_75t_L g3044 ( 
.A1(n_2650),
.A2(n_1493),
.B(n_1498),
.C(n_1491),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2767),
.B(n_1725),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2601),
.B(n_1726),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2581),
.B(n_1729),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2535),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2537),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_2583),
.A2(n_1194),
.B1(n_1380),
.B2(n_1224),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2656),
.B(n_1704),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2586),
.B(n_1500),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2538),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_SL g3054 ( 
.A(n_2661),
.B(n_1184),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2768),
.B(n_1202),
.Y(n_3055)
);

AND2x6_ASAP7_75t_SL g3056 ( 
.A(n_2573),
.B(n_1505),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2670),
.B(n_2501),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2542),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2591),
.B(n_1515),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2663),
.A2(n_1204),
.B1(n_1289),
.B2(n_1254),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2595),
.B(n_1520),
.Y(n_3061)
);

INVxp67_ASAP7_75t_L g3062 ( 
.A(n_2714),
.Y(n_3062)
);

HB1xp67_ASAP7_75t_L g3063 ( 
.A(n_2608),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2597),
.B(n_1527),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2402),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_L g3066 ( 
.A1(n_2603),
.A2(n_1337),
.B1(n_1341),
.B2(n_1314),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2606),
.B(n_2695),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2655),
.B(n_1528),
.Y(n_3068)
);

BUFx6f_ASAP7_75t_L g3069 ( 
.A(n_2713),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2693),
.B(n_1532),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2781),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2694),
.B(n_1534),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2662),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2698),
.B(n_1364),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2544),
.Y(n_3075)
);

INVx2_ASAP7_75t_SL g3076 ( 
.A(n_2687),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2666),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2545),
.Y(n_3078)
);

INVxp67_ASAP7_75t_L g3079 ( 
.A(n_2715),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2713),
.B(n_1371),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2553),
.Y(n_3081)
);

AOI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2636),
.A2(n_1407),
.B1(n_1412),
.B2(n_1383),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2554),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2557),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2685),
.B(n_1541),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_2444),
.A2(n_1587),
.B1(n_1611),
.B2(n_1507),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2558),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2713),
.B(n_1632),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2605),
.B(n_1664),
.Y(n_3089)
);

INVxp67_ASAP7_75t_L g3090 ( 
.A(n_2726),
.Y(n_3090)
);

NOR2x1_ASAP7_75t_L g3091 ( 
.A(n_2509),
.B(n_1542),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_L g3092 ( 
.A(n_2607),
.B(n_1547),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2732),
.A2(n_1551),
.B1(n_1555),
.B2(n_1548),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2673),
.B(n_1568),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2565),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2551),
.B(n_1573),
.Y(n_3096)
);

AND2x4_ASAP7_75t_SL g3097 ( 
.A(n_2720),
.B(n_1194),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2556),
.B(n_2727),
.Y(n_3098)
);

OAI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2722),
.A2(n_1380),
.B1(n_1416),
.B2(n_1224),
.Y(n_3099)
);

BUFx3_ASAP7_75t_L g3100 ( 
.A(n_2610),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2628),
.A2(n_1582),
.B(n_1574),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2525),
.B(n_1583),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2566),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2525),
.B(n_1586),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_SL g3105 ( 
.A(n_2720),
.B(n_1588),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2567),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_2720),
.B(n_1590),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2568),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2570),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2572),
.Y(n_3110)
);

NAND3xp33_ASAP7_75t_L g3111 ( 
.A(n_2773),
.B(n_1416),
.C(n_1380),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2674),
.Y(n_3112)
);

NOR2xp33_ASAP7_75t_L g3113 ( 
.A(n_2679),
.B(n_1593),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2675),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2525),
.B(n_1594),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2525),
.B(n_1597),
.Y(n_3116)
);

AND2x6_ASAP7_75t_SL g3117 ( 
.A(n_2737),
.B(n_1598),
.Y(n_3117)
);

O2A1O1Ixp5_ASAP7_75t_L g3118 ( 
.A1(n_2524),
.A2(n_1600),
.B(n_1607),
.C(n_1599),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2678),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2623),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2690),
.B(n_1608),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_2716),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_2585),
.A2(n_1610),
.B(n_1609),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2680),
.B(n_1620),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2625),
.B(n_1623),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2744),
.B(n_1628),
.Y(n_3126)
);

INVx8_ASAP7_75t_L g3127 ( 
.A(n_2728),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_2410),
.A2(n_1633),
.B(n_1630),
.Y(n_3128)
);

NAND2x1p5_ASAP7_75t_L g3129 ( 
.A(n_2728),
.B(n_1416),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_SL g3130 ( 
.A(n_2728),
.B(n_1636),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_L g3131 ( 
.A1(n_2626),
.A2(n_1641),
.B1(n_1642),
.B2(n_1638),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2634),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2751),
.B(n_1644),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2627),
.B(n_1645),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2630),
.B(n_1646),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2756),
.B(n_1653),
.Y(n_3136)
);

BUFx12f_ASAP7_75t_SL g3137 ( 
.A(n_2763),
.Y(n_3137)
);

INVx2_ASAP7_75t_SL g3138 ( 
.A(n_2681),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2631),
.B(n_1658),
.Y(n_3139)
);

OAI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2575),
.A2(n_1663),
.B(n_1659),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2632),
.Y(n_3141)
);

AND2x6_ASAP7_75t_L g3142 ( 
.A(n_2760),
.B(n_1416),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2637),
.B(n_1665),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_2683),
.B(n_2),
.Y(n_3144)
);

INVx2_ASAP7_75t_SL g3145 ( 
.A(n_2684),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2638),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2639),
.Y(n_3147)
);

OR2x6_ASAP7_75t_L g3148 ( 
.A(n_2686),
.B(n_1667),
.Y(n_3148)
);

AOI22xp33_ASAP7_75t_L g3149 ( 
.A1(n_2641),
.A2(n_1673),
.B1(n_1679),
.B2(n_1671),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2763),
.B(n_1692),
.Y(n_3150)
);

OAI22xp5_ASAP7_75t_SL g3151 ( 
.A1(n_2644),
.A2(n_1701),
.B1(n_1714),
.B2(n_1699),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2646),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2543),
.B(n_1724),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2543),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2701),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2702),
.Y(n_3156)
);

OR2x6_ASAP7_75t_L g3157 ( 
.A(n_2748),
.B(n_1727),
.Y(n_3157)
);

BUFx6f_ASAP7_75t_L g3158 ( 
.A(n_2412),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2754),
.B(n_1461),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2757),
.B(n_1461),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2417),
.B(n_1461),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_2730),
.B(n_2),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2733),
.Y(n_3163)
);

AO22x1_ASAP7_75t_L g3164 ( 
.A1(n_2766),
.A2(n_1635),
.B1(n_1461),
.B2(n_5),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2721),
.B(n_3),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2734),
.Y(n_3166)
);

AOI22xp33_ASAP7_75t_L g3167 ( 
.A1(n_2703),
.A2(n_1635),
.B1(n_5),
.B2(n_3),
.Y(n_3167)
);

NAND2xp33_ASAP7_75t_L g3168 ( 
.A(n_2761),
.B(n_1635),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2724),
.B(n_3),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2705),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2736),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2706),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2443),
.B(n_1635),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2712),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_3174)
);

AND2x4_ASAP7_75t_L g3175 ( 
.A(n_2725),
.B(n_4),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2718),
.Y(n_3176)
);

OAI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2453),
.A2(n_4),
.B(n_6),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_2762),
.B(n_7),
.Y(n_3178)
);

AND2x4_ASAP7_75t_L g3179 ( 
.A(n_2742),
.B(n_6),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2745),
.B(n_7),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2456),
.B(n_2459),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2521),
.B(n_8),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_L g3183 ( 
.A1(n_2750),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_3183)
);

OAI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2522),
.A2(n_8),
.B(n_9),
.Y(n_3184)
);

AOI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2752),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2549),
.B(n_12),
.Y(n_3186)
);

NOR3xp33_ASAP7_75t_L g3187 ( 
.A(n_2739),
.B(n_15),
.C(n_14),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2765),
.B(n_13),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2682),
.B(n_13),
.Y(n_3189)
);

CKINVDCx5p33_ASAP7_75t_R g3190 ( 
.A(n_2771),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2404),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2404),
.B(n_13),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2404),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2404),
.B(n_14),
.Y(n_3194)
);

NOR2xp67_ASAP7_75t_L g3195 ( 
.A(n_2405),
.B(n_15),
.Y(n_3195)
);

BUFx2_ASAP7_75t_SL g3196 ( 
.A(n_2771),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2559),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2404),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2404),
.Y(n_3199)
);

NOR2xp67_ASAP7_75t_SL g3200 ( 
.A(n_2555),
.B(n_16),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2404),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_2771),
.Y(n_3202)
);

AOI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_2559),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_2501),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_2480),
.B(n_20),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2404),
.B(n_19),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2404),
.Y(n_3207)
);

HB1xp67_ASAP7_75t_L g3208 ( 
.A(n_2405),
.Y(n_3208)
);

AND2x4_ASAP7_75t_L g3209 ( 
.A(n_2404),
.B(n_19),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2404),
.Y(n_3210)
);

AOI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_2559),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2404),
.Y(n_3212)
);

NOR2xp67_ASAP7_75t_L g3213 ( 
.A(n_2405),
.B(n_21),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2404),
.B(n_21),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2480),
.B(n_24),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_SL g3216 ( 
.A(n_2480),
.B(n_24),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2404),
.B(n_23),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2404),
.B(n_23),
.Y(n_3218)
);

NAND2xp33_ASAP7_75t_L g3219 ( 
.A(n_2543),
.B(n_25),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2404),
.B(n_24),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_2559),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2404),
.B(n_27),
.Y(n_3222)
);

NAND2x1_ASAP7_75t_L g3223 ( 
.A(n_2501),
.B(n_27),
.Y(n_3223)
);

NAND3xp33_ASAP7_75t_SL g3224 ( 
.A(n_2774),
.B(n_28),
.C(n_29),
.Y(n_3224)
);

AND2x6_ASAP7_75t_SL g3225 ( 
.A(n_2532),
.B(n_28),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2404),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2480),
.B(n_29),
.Y(n_3227)
);

NOR2xp33_ASAP7_75t_SL g3228 ( 
.A(n_2555),
.B(n_28),
.Y(n_3228)
);

BUFx3_ASAP7_75t_L g3229 ( 
.A(n_2540),
.Y(n_3229)
);

AOI22xp33_ASAP7_75t_L g3230 ( 
.A1(n_2559),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_3230)
);

NOR2xp67_ASAP7_75t_L g3231 ( 
.A(n_2405),
.B(n_30),
.Y(n_3231)
);

NAND2x1p5_ASAP7_75t_L g3232 ( 
.A(n_2474),
.B(n_31),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2404),
.B(n_32),
.Y(n_3233)
);

AOI22xp33_ASAP7_75t_L g3234 ( 
.A1(n_2559),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_3234)
);

AOI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_2405),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2404),
.Y(n_3236)
);

AOI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_2405),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2404),
.B(n_36),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2404),
.B(n_37),
.Y(n_3239)
);

NOR2xp67_ASAP7_75t_L g3240 ( 
.A(n_2405),
.B(n_38),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2404),
.B(n_38),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_2480),
.B(n_40),
.Y(n_3242)
);

NAND3xp33_ASAP7_75t_SL g3243 ( 
.A(n_2774),
.B(n_39),
.C(n_40),
.Y(n_3243)
);

OAI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_2403),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2404),
.B(n_41),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_2405),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2404),
.B(n_42),
.Y(n_3247)
);

OR2x2_ASAP7_75t_L g3248 ( 
.A(n_2405),
.B(n_42),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_2480),
.B(n_44),
.Y(n_3249)
);

AND2x6_ASAP7_75t_L g3250 ( 
.A(n_2624),
.B(n_43),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_2489),
.A2(n_43),
.B(n_44),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2404),
.B(n_43),
.Y(n_3252)
);

OR2x6_ASAP7_75t_L g3253 ( 
.A(n_2436),
.B(n_44),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2404),
.B(n_45),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2404),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_SL g3256 ( 
.A(n_2480),
.B(n_46),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2404),
.Y(n_3257)
);

AND2x6_ASAP7_75t_SL g3258 ( 
.A(n_2532),
.B(n_45),
.Y(n_3258)
);

NOR2xp33_ASAP7_75t_L g3259 ( 
.A(n_2550),
.B(n_45),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_2559),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_3260)
);

NOR2xp67_ASAP7_75t_L g3261 ( 
.A(n_2405),
.B(n_46),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2404),
.B(n_47),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2404),
.B(n_47),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2404),
.B(n_48),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2404),
.B(n_48),
.Y(n_3265)
);

NOR2x1_ASAP7_75t_L g3266 ( 
.A(n_2436),
.B(n_50),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2404),
.B(n_50),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2404),
.B(n_50),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_2403),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_R g3270 ( 
.A(n_2771),
.B(n_52),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_2559),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_2540),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2404),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_L g3274 ( 
.A(n_2550),
.B(n_54),
.Y(n_3274)
);

AOI22xp33_ASAP7_75t_L g3275 ( 
.A1(n_2559),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3275)
);

INVx4_ASAP7_75t_L g3276 ( 
.A(n_2555),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_2480),
.B(n_56),
.Y(n_3277)
);

O2A1O1Ixp33_ASAP7_75t_L g3278 ( 
.A1(n_2411),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2404),
.B(n_57),
.Y(n_3279)
);

AND2x4_ASAP7_75t_L g3280 ( 
.A(n_2404),
.B(n_58),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2404),
.B(n_58),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2404),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2550),
.B(n_58),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2404),
.B(n_59),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2404),
.B(n_59),
.Y(n_3285)
);

NOR3x1_ASAP7_75t_L g3286 ( 
.A(n_2405),
.B(n_59),
.C(n_60),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2404),
.B(n_60),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2404),
.B(n_60),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2404),
.B(n_61),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2404),
.B(n_61),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2404),
.Y(n_3291)
);

INVx2_ASAP7_75t_SL g3292 ( 
.A(n_2405),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2404),
.B(n_62),
.Y(n_3293)
);

INVx2_ASAP7_75t_SL g3294 ( 
.A(n_2405),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2404),
.B(n_62),
.Y(n_3295)
);

INVx3_ASAP7_75t_L g3296 ( 
.A(n_2759),
.Y(n_3296)
);

AOI22xp33_ASAP7_75t_L g3297 ( 
.A1(n_2559),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2404),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2404),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2404),
.Y(n_3300)
);

AND2x6_ASAP7_75t_SL g3301 ( 
.A(n_2532),
.B(n_63),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2404),
.B(n_63),
.Y(n_3302)
);

INVx4_ASAP7_75t_L g3303 ( 
.A(n_2555),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_2759),
.Y(n_3304)
);

AO22x1_ASAP7_75t_L g3305 ( 
.A1(n_2649),
.A2(n_66),
.B1(n_67),
.B2(n_65),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2404),
.B(n_64),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2404),
.B(n_65),
.Y(n_3307)
);

NOR2xp67_ASAP7_75t_L g3308 ( 
.A(n_2405),
.B(n_65),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2404),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_2404),
.Y(n_3310)
);

AND2x4_ASAP7_75t_SL g3311 ( 
.A(n_2540),
.B(n_66),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_2559),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_3312)
);

BUFx8_ASAP7_75t_L g3313 ( 
.A(n_2493),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2404),
.B(n_67),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_2480),
.B(n_69),
.Y(n_3315)
);

NAND3xp33_ASAP7_75t_SL g3316 ( 
.A(n_2774),
.B(n_68),
.C(n_69),
.Y(n_3316)
);

AND2x6_ASAP7_75t_L g3317 ( 
.A(n_2624),
.B(n_70),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_SL g3318 ( 
.A(n_2480),
.B(n_71),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_2403),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_2404),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2404),
.B(n_70),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2404),
.Y(n_3322)
);

INVx5_ASAP7_75t_L g3323 ( 
.A(n_2671),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2404),
.B(n_71),
.Y(n_3324)
);

NOR2xp67_ASAP7_75t_L g3325 ( 
.A(n_2405),
.B(n_72),
.Y(n_3325)
);

BUFx6f_ASAP7_75t_L g3326 ( 
.A(n_2501),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2404),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2404),
.B(n_73),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_2489),
.A2(n_73),
.B(n_74),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_2404),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2404),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_2550),
.B(n_73),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2404),
.B(n_74),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2404),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_2404),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2404),
.B(n_75),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_2404),
.B(n_75),
.Y(n_3337)
);

BUFx3_ASAP7_75t_L g3338 ( 
.A(n_2540),
.Y(n_3338)
);

OR2x2_ASAP7_75t_L g3339 ( 
.A(n_2405),
.B(n_76),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2404),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2404),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_2405),
.B(n_76),
.Y(n_3342)
);

AOI22xp33_ASAP7_75t_L g3343 ( 
.A1(n_2559),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_2550),
.B(n_77),
.Y(n_3344)
);

AOI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_2405),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_3345)
);

NAND2x1_ASAP7_75t_L g3346 ( 
.A(n_2501),
.B(n_79),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_2559),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_2404),
.B(n_80),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_2404),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2404),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2404),
.B(n_81),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2404),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_2404),
.B(n_81),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2404),
.B(n_82),
.Y(n_3354)
);

OR2x2_ASAP7_75t_L g3355 ( 
.A(n_2405),
.B(n_82),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2404),
.B(n_83),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_2559),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_3357)
);

INVx2_ASAP7_75t_SL g3358 ( 
.A(n_2405),
.Y(n_3358)
);

NOR2xp33_ASAP7_75t_L g3359 ( 
.A(n_2550),
.B(n_84),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_2405),
.B(n_84),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_2404),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2404),
.B(n_85),
.Y(n_3362)
);

INVxp33_ASAP7_75t_L g3363 ( 
.A(n_2425),
.Y(n_3363)
);

OR2x2_ASAP7_75t_L g3364 ( 
.A(n_2405),
.B(n_86),
.Y(n_3364)
);

NAND2xp33_ASAP7_75t_L g3365 ( 
.A(n_2543),
.B(n_88),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2404),
.B(n_87),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_2404),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_2404),
.B(n_87),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2550),
.B(n_87),
.Y(n_3369)
);

INVxp67_ASAP7_75t_L g3370 ( 
.A(n_2405),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_2404),
.B(n_88),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2550),
.B(n_88),
.Y(n_3372)
);

INVx2_ASAP7_75t_SL g3373 ( 
.A(n_2405),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2404),
.B(n_89),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2404),
.B(n_89),
.Y(n_3375)
);

BUFx12f_ASAP7_75t_L g3376 ( 
.A(n_2406),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2404),
.B(n_89),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_2405),
.B(n_90),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_2405),
.B(n_90),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2404),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_2559),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_3381)
);

O2A1O1Ixp5_ASAP7_75t_L g3382 ( 
.A1(n_2494),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2404),
.B(n_91),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_L g3384 ( 
.A(n_2550),
.B(n_94),
.Y(n_3384)
);

OR2x6_ASAP7_75t_L g3385 ( 
.A(n_2436),
.B(n_94),
.Y(n_3385)
);

INVxp67_ASAP7_75t_SL g3386 ( 
.A(n_2405),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_2480),
.B(n_96),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2404),
.B(n_95),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_2404),
.B(n_95),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_2550),
.B(n_95),
.Y(n_3390)
);

OAI22xp33_ASAP7_75t_SL g3391 ( 
.A1(n_2774),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_2480),
.B(n_97),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2404),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_SL g3394 ( 
.A(n_2480),
.B(n_97),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_2404),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_2550),
.B(n_96),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2404),
.B(n_98),
.Y(n_3397)
);

BUFx6f_ASAP7_75t_SL g3398 ( 
.A(n_2436),
.Y(n_3398)
);

AOI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_2405),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_3399)
);

AOI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_2405),
.A2(n_102),
.B1(n_99),
.B2(n_101),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2404),
.B(n_101),
.Y(n_3401)
);

AOI22xp5_ASAP7_75t_L g3402 ( 
.A1(n_2405),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2404),
.B(n_103),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2404),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_2404),
.B(n_103),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2404),
.B(n_105),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2404),
.B(n_105),
.Y(n_3407)
);

OAI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_2489),
.A2(n_106),
.B(n_107),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2404),
.B(n_106),
.Y(n_3409)
);

INVx3_ASAP7_75t_L g3410 ( 
.A(n_2759),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_2559),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_3411)
);

NOR3xp33_ASAP7_75t_SL g3412 ( 
.A(n_2665),
.B(n_107),
.C(n_108),
.Y(n_3412)
);

AND2x6_ASAP7_75t_SL g3413 ( 
.A(n_2532),
.B(n_108),
.Y(n_3413)
);

O2A1O1Ixp33_ASAP7_75t_L g3414 ( 
.A1(n_2411),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_3414)
);

INVx3_ASAP7_75t_L g3415 ( 
.A(n_2759),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2404),
.Y(n_3416)
);

OR2x2_ASAP7_75t_L g3417 ( 
.A(n_2405),
.B(n_109),
.Y(n_3417)
);

BUFx3_ASAP7_75t_L g3418 ( 
.A(n_2540),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2404),
.B(n_110),
.Y(n_3419)
);

O2A1O1Ixp33_ASAP7_75t_L g3420 ( 
.A1(n_2411),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2404),
.B(n_111),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_2480),
.B(n_113),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_2480),
.B(n_113),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2404),
.Y(n_3424)
);

OR2x2_ASAP7_75t_L g3425 ( 
.A(n_2405),
.B(n_112),
.Y(n_3425)
);

AO221x1_ASAP7_75t_L g3426 ( 
.A1(n_2774),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.C(n_115),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2404),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2404),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2404),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_2404),
.B(n_114),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_2550),
.B(n_114),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2404),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2404),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_2550),
.B(n_115),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2404),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2404),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_2405),
.B(n_116),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_2404),
.B(n_116),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2404),
.B(n_116),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_SL g3440 ( 
.A(n_2555),
.B(n_118),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_2559),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_2480),
.B(n_119),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2404),
.Y(n_3443)
);

NAND2xp33_ASAP7_75t_SL g3444 ( 
.A(n_2592),
.B(n_118),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_2404),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_2480),
.B(n_120),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_2404),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_2404),
.Y(n_3448)
);

CKINVDCx5p33_ASAP7_75t_R g3449 ( 
.A(n_2771),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_2791),
.B(n_119),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_2794),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_2791),
.B(n_120),
.Y(n_3452)
);

INVxp67_ASAP7_75t_L g3453 ( 
.A(n_3208),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_3076),
.B(n_121),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_2795),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3436),
.Y(n_3456)
);

BUFx6f_ASAP7_75t_L g3457 ( 
.A(n_3127),
.Y(n_3457)
);

AOI22x1_ASAP7_75t_SL g3458 ( 
.A1(n_2919),
.A2(n_2899),
.B1(n_3202),
.B2(n_3190),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3447),
.Y(n_3459)
);

INVx3_ASAP7_75t_L g3460 ( 
.A(n_2842),
.Y(n_3460)
);

INVxp67_ASAP7_75t_L g3461 ( 
.A(n_2875),
.Y(n_3461)
);

CKINVDCx20_ASAP7_75t_R g3462 ( 
.A(n_2802),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_2941),
.B(n_121),
.Y(n_3463)
);

BUFx3_ASAP7_75t_L g3464 ( 
.A(n_3229),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3198),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_2863),
.B(n_121),
.Y(n_3466)
);

OR2x2_ASAP7_75t_L g3467 ( 
.A(n_2993),
.B(n_122),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3130),
.B(n_1015),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3199),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3201),
.Y(n_3470)
);

INVx5_ASAP7_75t_L g3471 ( 
.A(n_3253),
.Y(n_3471)
);

INVx4_ASAP7_75t_L g3472 ( 
.A(n_2866),
.Y(n_3472)
);

BUFx2_ASAP7_75t_L g3473 ( 
.A(n_3179),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3236),
.Y(n_3474)
);

BUFx2_ASAP7_75t_L g3475 ( 
.A(n_3179),
.Y(n_3475)
);

INVx5_ASAP7_75t_L g3476 ( 
.A(n_3253),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2792),
.B(n_122),
.Y(n_3477)
);

AND2x4_ASAP7_75t_L g3478 ( 
.A(n_2842),
.B(n_122),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_2793),
.B(n_123),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3191),
.B(n_123),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_3127),
.Y(n_3481)
);

BUFx3_ASAP7_75t_L g3482 ( 
.A(n_3272),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3273),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3193),
.B(n_123),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3300),
.Y(n_3485)
);

BUFx2_ASAP7_75t_L g3486 ( 
.A(n_2875),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3309),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3310),
.Y(n_3488)
);

INVx5_ASAP7_75t_L g3489 ( 
.A(n_3253),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3207),
.B(n_124),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3320),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_2802),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3330),
.Y(n_3493)
);

INVx2_ASAP7_75t_SL g3494 ( 
.A(n_2866),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3210),
.B(n_124),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3433),
.Y(n_3496)
);

INVx8_ASAP7_75t_L g3497 ( 
.A(n_2866),
.Y(n_3497)
);

INVx3_ASAP7_75t_L g3498 ( 
.A(n_2843),
.Y(n_3498)
);

INVxp67_ASAP7_75t_L g3499 ( 
.A(n_2875),
.Y(n_3499)
);

AND2x4_ASAP7_75t_L g3500 ( 
.A(n_2845),
.B(n_125),
.Y(n_3500)
);

BUFx3_ASAP7_75t_L g3501 ( 
.A(n_3338),
.Y(n_3501)
);

NAND2xp33_ASAP7_75t_L g3502 ( 
.A(n_3016),
.B(n_126),
.Y(n_3502)
);

OR2x6_ASAP7_75t_L g3503 ( 
.A(n_3385),
.B(n_126),
.Y(n_3503)
);

OR2x6_ASAP7_75t_L g3504 ( 
.A(n_3385),
.B(n_126),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3370),
.Y(n_3505)
);

NAND3xp33_ASAP7_75t_SL g3506 ( 
.A(n_3270),
.B(n_2838),
.C(n_2948),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3212),
.B(n_127),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3226),
.B(n_127),
.Y(n_3508)
);

INVx2_ASAP7_75t_SL g3509 ( 
.A(n_2988),
.Y(n_3509)
);

NAND2xp33_ASAP7_75t_SL g3510 ( 
.A(n_3200),
.B(n_128),
.Y(n_3510)
);

AND2x4_ASAP7_75t_L g3511 ( 
.A(n_3335),
.B(n_128),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3043),
.B(n_128),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3340),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_R g3514 ( 
.A(n_3449),
.B(n_129),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_2850),
.B(n_129),
.Y(n_3515)
);

AND2x4_ASAP7_75t_L g3516 ( 
.A(n_3361),
.B(n_129),
.Y(n_3516)
);

INVx4_ASAP7_75t_L g3517 ( 
.A(n_3385),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3255),
.B(n_130),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_SL g3519 ( 
.A(n_3130),
.B(n_1016),
.Y(n_3519)
);

AND2x4_ASAP7_75t_L g3520 ( 
.A(n_3367),
.B(n_3393),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3257),
.B(n_130),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3395),
.Y(n_3522)
);

INVx2_ASAP7_75t_SL g3523 ( 
.A(n_2988),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3427),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3282),
.B(n_131),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3291),
.Y(n_3526)
);

INVx4_ASAP7_75t_L g3527 ( 
.A(n_2843),
.Y(n_3527)
);

AOI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_2819),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_3528)
);

NOR3xp33_ASAP7_75t_SL g3529 ( 
.A(n_2931),
.B(n_131),
.C(n_132),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_SL g3530 ( 
.A(n_2838),
.B(n_1016),
.Y(n_3530)
);

AND3x1_ASAP7_75t_SL g3531 ( 
.A(n_2943),
.B(n_133),
.C(n_135),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3298),
.Y(n_3532)
);

INVx1_ASAP7_75t_SL g3533 ( 
.A(n_2805),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3418),
.Y(n_3534)
);

BUFx2_ASAP7_75t_L g3535 ( 
.A(n_3016),
.Y(n_3535)
);

BUFx2_ASAP7_75t_L g3536 ( 
.A(n_3016),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3299),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3322),
.B(n_3327),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3331),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_2975),
.Y(n_3540)
);

OAI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_2948),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_3541)
);

AND2x4_ASAP7_75t_L g3542 ( 
.A(n_3334),
.B(n_135),
.Y(n_3542)
);

BUFx6f_ASAP7_75t_L g3543 ( 
.A(n_3127),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3341),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3349),
.B(n_136),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3350),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3352),
.Y(n_3547)
);

NOR3xp33_ASAP7_75t_SL g3548 ( 
.A(n_3122),
.B(n_136),
.C(n_137),
.Y(n_3548)
);

AOI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_2897),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3380),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3404),
.B(n_138),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3416),
.Y(n_3552)
);

AOI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_2918),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3424),
.Y(n_3554)
);

AND2x4_ASAP7_75t_L g3555 ( 
.A(n_3428),
.B(n_140),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3429),
.Y(n_3556)
);

A2O1A1Ixp33_ASAP7_75t_L g3557 ( 
.A1(n_2965),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_3557)
);

BUFx2_ASAP7_75t_L g3558 ( 
.A(n_3209),
.Y(n_3558)
);

AND3x1_ASAP7_75t_SL g3559 ( 
.A(n_3225),
.B(n_141),
.C(n_142),
.Y(n_3559)
);

INVx2_ASAP7_75t_SL g3560 ( 
.A(n_3313),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_3313),
.Y(n_3561)
);

NOR3xp33_ASAP7_75t_SL g3562 ( 
.A(n_3098),
.B(n_141),
.C(n_142),
.Y(n_3562)
);

BUFx3_ASAP7_75t_L g3563 ( 
.A(n_2909),
.Y(n_3563)
);

CKINVDCx14_ASAP7_75t_R g3564 ( 
.A(n_3376),
.Y(n_3564)
);

NOR3xp33_ASAP7_75t_SL g3565 ( 
.A(n_2829),
.B(n_143),
.C(n_144),
.Y(n_3565)
);

NOR3xp33_ASAP7_75t_SL g3566 ( 
.A(n_3099),
.B(n_143),
.C(n_144),
.Y(n_3566)
);

INVx5_ASAP7_75t_L g3567 ( 
.A(n_2851),
.Y(n_3567)
);

INVx4_ASAP7_75t_SL g3568 ( 
.A(n_3398),
.Y(n_3568)
);

INVx4_ASAP7_75t_L g3569 ( 
.A(n_3398),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_R g3570 ( 
.A(n_3137),
.B(n_144),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_2997),
.Y(n_3571)
);

BUFx2_ASAP7_75t_L g3572 ( 
.A(n_3209),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3432),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3435),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3443),
.Y(n_3575)
);

INVx4_ASAP7_75t_L g3576 ( 
.A(n_2874),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_2867),
.B(n_2869),
.Y(n_3577)
);

A2O1A1Ixp33_ASAP7_75t_L g3578 ( 
.A1(n_2853),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3445),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3448),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_2855),
.Y(n_3581)
);

INVx3_ASAP7_75t_L g3582 ( 
.A(n_2874),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3025),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3192),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_2884),
.Y(n_3585)
);

INVx3_ASAP7_75t_L g3586 ( 
.A(n_2939),
.Y(n_3586)
);

AND2x4_ASAP7_75t_L g3587 ( 
.A(n_3148),
.B(n_145),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_2894),
.Y(n_3588)
);

CKINVDCx20_ASAP7_75t_R g3589 ( 
.A(n_3311),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3192),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_2900),
.Y(n_3591)
);

INVx4_ASAP7_75t_L g3592 ( 
.A(n_2939),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_2978),
.B(n_148),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_SL g3594 ( 
.A(n_3228),
.B(n_3440),
.Y(n_3594)
);

BUFx6f_ASAP7_75t_L g3595 ( 
.A(n_3069),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_2980),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_3596)
);

CKINVDCx5p33_ASAP7_75t_R g3597 ( 
.A(n_3196),
.Y(n_3597)
);

AOI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_2914),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3044),
.B(n_149),
.Y(n_3599)
);

AND2x4_ASAP7_75t_L g3600 ( 
.A(n_3148),
.B(n_150),
.Y(n_3600)
);

OR2x6_ASAP7_75t_L g3601 ( 
.A(n_3232),
.B(n_151),
.Y(n_3601)
);

BUFx3_ASAP7_75t_L g3602 ( 
.A(n_2882),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_2800),
.B(n_151),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_2807),
.B(n_152),
.Y(n_3604)
);

BUFx12f_ASAP7_75t_L g3605 ( 
.A(n_3258),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_3301),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3194),
.Y(n_3607)
);

BUFx4f_ASAP7_75t_SL g3608 ( 
.A(n_2815),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3194),
.Y(n_3609)
);

BUFx2_ASAP7_75t_L g3610 ( 
.A(n_3280),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_2809),
.B(n_152),
.Y(n_3611)
);

INVx5_ASAP7_75t_L g3612 ( 
.A(n_3250),
.Y(n_3612)
);

BUFx6f_ASAP7_75t_L g3613 ( 
.A(n_3069),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_3148),
.B(n_152),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3009),
.B(n_153),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_3413),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3206),
.Y(n_3617)
);

INVx4_ASAP7_75t_L g3618 ( 
.A(n_2974),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_2857),
.B(n_153),
.Y(n_3619)
);

BUFx2_ASAP7_75t_L g3620 ( 
.A(n_3280),
.Y(n_3620)
);

INVx3_ASAP7_75t_L g3621 ( 
.A(n_2974),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_2912),
.Y(n_3622)
);

AOI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_2852),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_3623)
);

BUFx3_ASAP7_75t_L g3624 ( 
.A(n_2893),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_3014),
.Y(n_3625)
);

INVx3_ASAP7_75t_L g3626 ( 
.A(n_2974),
.Y(n_3626)
);

INVx5_ASAP7_75t_L g3627 ( 
.A(n_3250),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3206),
.Y(n_3628)
);

CKINVDCx5p33_ASAP7_75t_R g3629 ( 
.A(n_2989),
.Y(n_3629)
);

OR2x6_ASAP7_75t_L g3630 ( 
.A(n_3232),
.B(n_154),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_2817),
.B(n_154),
.Y(n_3631)
);

INVx5_ASAP7_75t_L g3632 ( 
.A(n_3250),
.Y(n_3632)
);

AND2x4_ASAP7_75t_L g3633 ( 
.A(n_2820),
.B(n_155),
.Y(n_3633)
);

AND2x4_ASAP7_75t_L g3634 ( 
.A(n_2826),
.B(n_155),
.Y(n_3634)
);

NOR3xp33_ASAP7_75t_SL g3635 ( 
.A(n_3099),
.B(n_156),
.C(n_157),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3290),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3290),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_2921),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_2935),
.Y(n_3639)
);

AND2x4_ASAP7_75t_L g3640 ( 
.A(n_2827),
.B(n_2830),
.Y(n_3640)
);

AOI22xp33_ASAP7_75t_SL g3641 ( 
.A1(n_3228),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_3641)
);

INVx5_ASAP7_75t_L g3642 ( 
.A(n_3250),
.Y(n_3642)
);

INVx3_ASAP7_75t_L g3643 ( 
.A(n_3276),
.Y(n_3643)
);

CKINVDCx5p33_ASAP7_75t_R g3644 ( 
.A(n_3029),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3409),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3409),
.Y(n_3646)
);

INVx3_ASAP7_75t_L g3647 ( 
.A(n_3276),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_2831),
.B(n_156),
.Y(n_3648)
);

AND3x2_ASAP7_75t_SL g3649 ( 
.A(n_3286),
.B(n_157),
.C(n_158),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_2947),
.B(n_159),
.Y(n_3650)
);

XNOR2xp5_ASAP7_75t_L g3651 ( 
.A(n_3363),
.B(n_159),
.Y(n_3651)
);

BUFx6f_ASAP7_75t_L g3652 ( 
.A(n_3069),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3419),
.Y(n_3653)
);

BUFx2_ASAP7_75t_L g3654 ( 
.A(n_3317),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_2910),
.B(n_159),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_3041),
.B(n_160),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3017),
.B(n_160),
.Y(n_3657)
);

AND2x4_ASAP7_75t_L g3658 ( 
.A(n_2971),
.B(n_2976),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_2944),
.Y(n_3659)
);

BUFx6f_ASAP7_75t_L g3660 ( 
.A(n_3204),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_R g3661 ( 
.A(n_3440),
.B(n_160),
.Y(n_3661)
);

OR2x2_ASAP7_75t_L g3662 ( 
.A(n_3024),
.B(n_161),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3419),
.Y(n_3663)
);

NOR2xp67_ASAP7_75t_L g3664 ( 
.A(n_3000),
.B(n_2824),
.Y(n_3664)
);

BUFx6f_ASAP7_75t_L g3665 ( 
.A(n_3204),
.Y(n_3665)
);

OR2x6_ASAP7_75t_L g3666 ( 
.A(n_3303),
.B(n_161),
.Y(n_3666)
);

AO22x1_ASAP7_75t_L g3667 ( 
.A1(n_3317),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_3667)
);

BUFx6f_ASAP7_75t_L g3668 ( 
.A(n_3204),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3421),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_2798),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_SL g3671 ( 
.A(n_2928),
.B(n_1017),
.Y(n_3671)
);

INVx3_ASAP7_75t_L g3672 ( 
.A(n_3303),
.Y(n_3672)
);

INVx2_ASAP7_75t_SL g3673 ( 
.A(n_2906),
.Y(n_3673)
);

INVx3_ASAP7_75t_L g3674 ( 
.A(n_3042),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3421),
.Y(n_3675)
);

HB1xp67_ASAP7_75t_L g3676 ( 
.A(n_3246),
.Y(n_3676)
);

OR2x6_ASAP7_75t_L g3677 ( 
.A(n_2954),
.B(n_162),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_2871),
.B(n_162),
.Y(n_3678)
);

BUFx6f_ASAP7_75t_L g3679 ( 
.A(n_3326),
.Y(n_3679)
);

BUFx2_ASAP7_75t_L g3680 ( 
.A(n_3317),
.Y(n_3680)
);

CKINVDCx5p33_ASAP7_75t_R g3681 ( 
.A(n_3056),
.Y(n_3681)
);

BUFx12f_ASAP7_75t_L g3682 ( 
.A(n_2956),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_2839),
.B(n_2904),
.Y(n_3683)
);

INVx4_ASAP7_75t_L g3684 ( 
.A(n_2813),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_2806),
.Y(n_3685)
);

AOI211xp5_ASAP7_75t_L g3686 ( 
.A1(n_3305),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_2888),
.B(n_164),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_2983),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3005),
.Y(n_3689)
);

AO22x1_ASAP7_75t_L g3690 ( 
.A1(n_3317),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_3117),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_2961),
.B(n_166),
.Y(n_3692)
);

AOI221xp5_ASAP7_75t_L g3693 ( 
.A1(n_2892),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.C(n_169),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_2959),
.Y(n_3694)
);

HB1xp67_ASAP7_75t_L g3695 ( 
.A(n_3292),
.Y(n_3695)
);

INVx4_ASAP7_75t_L g3696 ( 
.A(n_2813),
.Y(n_3696)
);

BUFx3_ASAP7_75t_L g3697 ( 
.A(n_3294),
.Y(n_3697)
);

CKINVDCx5p33_ASAP7_75t_R g3698 ( 
.A(n_2982),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3093),
.B(n_167),
.Y(n_3699)
);

NAND2x1p5_ASAP7_75t_L g3700 ( 
.A(n_2812),
.B(n_168),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_2841),
.Y(n_3701)
);

INVx4_ASAP7_75t_L g3702 ( 
.A(n_2812),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_2932),
.B(n_1018),
.Y(n_3703)
);

AND2x4_ASAP7_75t_L g3704 ( 
.A(n_2861),
.B(n_168),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_SL g3705 ( 
.A(n_3195),
.B(n_1018),
.Y(n_3705)
);

AOI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_2883),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_3706)
);

NOR2xp33_ASAP7_75t_L g3707 ( 
.A(n_3067),
.B(n_3062),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3035),
.B(n_169),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_2879),
.Y(n_3709)
);

BUFx3_ASAP7_75t_L g3710 ( 
.A(n_3358),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_2811),
.Y(n_3711)
);

AND2x4_ASAP7_75t_L g3712 ( 
.A(n_2895),
.B(n_170),
.Y(n_3712)
);

AOI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3096),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_3713)
);

INVx3_ASAP7_75t_L g3714 ( 
.A(n_3100),
.Y(n_3714)
);

CKINVDCx5p33_ASAP7_75t_R g3715 ( 
.A(n_2984),
.Y(n_3715)
);

BUFx2_ASAP7_75t_L g3716 ( 
.A(n_2812),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3123),
.B(n_171),
.Y(n_3717)
);

INVx4_ASAP7_75t_L g3718 ( 
.A(n_2847),
.Y(n_3718)
);

AND2x6_ASAP7_75t_L g3719 ( 
.A(n_3175),
.B(n_3326),
.Y(n_3719)
);

AND3x1_ASAP7_75t_SL g3720 ( 
.A(n_2877),
.B(n_172),
.C(n_173),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_2828),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_2992),
.B(n_173),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3022),
.B(n_2878),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_2896),
.Y(n_3724)
);

OAI22xp5_ASAP7_75t_SL g3725 ( 
.A1(n_2933),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_3725)
);

AND3x1_ASAP7_75t_L g3726 ( 
.A(n_3412),
.B(n_174),
.C(n_175),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_2902),
.Y(n_3727)
);

INVx4_ASAP7_75t_L g3728 ( 
.A(n_2847),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_2917),
.Y(n_3729)
);

AND2x4_ASAP7_75t_L g3730 ( 
.A(n_2927),
.B(n_174),
.Y(n_3730)
);

AOI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3151),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_2994),
.B(n_176),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_SL g3733 ( 
.A(n_3213),
.B(n_1019),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_SL g3734 ( 
.A(n_3231),
.B(n_1019),
.Y(n_3734)
);

NOR2x1p5_ASAP7_75t_SL g3735 ( 
.A(n_2929),
.B(n_1020),
.Y(n_3735)
);

CKINVDCx5p33_ASAP7_75t_R g3736 ( 
.A(n_3373),
.Y(n_3736)
);

INVx2_ASAP7_75t_SL g3737 ( 
.A(n_3132),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_2938),
.Y(n_3738)
);

OR2x6_ASAP7_75t_L g3739 ( 
.A(n_2876),
.B(n_176),
.Y(n_3739)
);

HB1xp67_ASAP7_75t_L g3740 ( 
.A(n_3175),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_2949),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_2960),
.Y(n_3742)
);

BUFx3_ASAP7_75t_L g3743 ( 
.A(n_2905),
.Y(n_3743)
);

INVx2_ASAP7_75t_SL g3744 ( 
.A(n_3248),
.Y(n_3744)
);

INVxp33_ASAP7_75t_L g3745 ( 
.A(n_2973),
.Y(n_3745)
);

BUFx2_ASAP7_75t_L g3746 ( 
.A(n_2847),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3188),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_2814),
.B(n_177),
.Y(n_3748)
);

CKINVDCx5p33_ASAP7_75t_R g3749 ( 
.A(n_3031),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3188),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_2854),
.Y(n_3751)
);

INVx4_ASAP7_75t_L g3752 ( 
.A(n_2942),
.Y(n_3752)
);

INVx4_ASAP7_75t_L g3753 ( 
.A(n_2942),
.Y(n_3753)
);

AOI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_2968),
.A2(n_3028),
.B1(n_2977),
.B2(n_2995),
.Y(n_3754)
);

AOI22xp33_ASAP7_75t_L g3755 ( 
.A1(n_3259),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3048),
.Y(n_3756)
);

OR2x6_ASAP7_75t_L g3757 ( 
.A(n_3240),
.B(n_178),
.Y(n_3757)
);

NOR3xp33_ASAP7_75t_SL g3758 ( 
.A(n_3224),
.B(n_178),
.C(n_179),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_2814),
.B(n_180),
.Y(n_3759)
);

HB1xp67_ASAP7_75t_L g3760 ( 
.A(n_2797),
.Y(n_3760)
);

INVx2_ASAP7_75t_SL g3761 ( 
.A(n_3339),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_2818),
.B(n_180),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_2818),
.B(n_180),
.Y(n_3763)
);

HB1xp67_ASAP7_75t_L g3764 ( 
.A(n_3386),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3049),
.Y(n_3765)
);

NOR3xp33_ASAP7_75t_SL g3766 ( 
.A(n_3243),
.B(n_181),
.C(n_182),
.Y(n_3766)
);

INVxp67_ASAP7_75t_SL g3767 ( 
.A(n_3219),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3079),
.B(n_181),
.Y(n_3768)
);

NOR3xp33_ASAP7_75t_SL g3769 ( 
.A(n_3316),
.B(n_181),
.C(n_182),
.Y(n_3769)
);

NOR2xp33_ASAP7_75t_L g3770 ( 
.A(n_3090),
.B(n_182),
.Y(n_3770)
);

BUFx4f_ASAP7_75t_L g3771 ( 
.A(n_3355),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_2823),
.B(n_183),
.Y(n_3772)
);

BUFx2_ASAP7_75t_L g3773 ( 
.A(n_2942),
.Y(n_3773)
);

HB1xp67_ASAP7_75t_L g3774 ( 
.A(n_3180),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3078),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_2891),
.B(n_3002),
.Y(n_3776)
);

INVx3_ASAP7_75t_L g3777 ( 
.A(n_3081),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3083),
.Y(n_3778)
);

AOI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_2987),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_2823),
.B(n_184),
.Y(n_3780)
);

AND3x1_ASAP7_75t_SL g3781 ( 
.A(n_2966),
.B(n_185),
.C(n_186),
.Y(n_3781)
);

INVxp67_ASAP7_75t_L g3782 ( 
.A(n_3364),
.Y(n_3782)
);

OR2x6_ASAP7_75t_L g3783 ( 
.A(n_3261),
.B(n_185),
.Y(n_3783)
);

NOR2x1p5_ASAP7_75t_L g3784 ( 
.A(n_2946),
.B(n_186),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3053),
.Y(n_3785)
);

BUFx6f_ASAP7_75t_L g3786 ( 
.A(n_3326),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3058),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_2825),
.B(n_186),
.Y(n_3788)
);

BUFx3_ASAP7_75t_L g3789 ( 
.A(n_3342),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_2825),
.B(n_187),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3095),
.Y(n_3791)
);

NOR2xp67_ASAP7_75t_L g3792 ( 
.A(n_3323),
.B(n_187),
.Y(n_3792)
);

AND2x4_ASAP7_75t_L g3793 ( 
.A(n_3075),
.B(n_188),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3084),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_2835),
.B(n_189),
.Y(n_3795)
);

BUFx6f_ASAP7_75t_L g3796 ( 
.A(n_3323),
.Y(n_3796)
);

NOR3xp33_ASAP7_75t_SL g3797 ( 
.A(n_2985),
.B(n_189),
.C(n_190),
.Y(n_3797)
);

NOR3xp33_ASAP7_75t_SL g3798 ( 
.A(n_3205),
.B(n_189),
.C(n_190),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3087),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3103),
.Y(n_3800)
);

NOR2xp67_ASAP7_75t_L g3801 ( 
.A(n_3323),
.B(n_191),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3110),
.Y(n_3802)
);

INVx3_ASAP7_75t_L g3803 ( 
.A(n_3112),
.Y(n_3803)
);

BUFx6f_ASAP7_75t_L g3804 ( 
.A(n_2964),
.Y(n_3804)
);

BUFx12f_ASAP7_75t_L g3805 ( 
.A(n_3417),
.Y(n_3805)
);

BUFx6f_ASAP7_75t_L g3806 ( 
.A(n_2964),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3141),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3146),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3106),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3152),
.Y(n_3810)
);

AND2x4_ASAP7_75t_L g3811 ( 
.A(n_3108),
.B(n_191),
.Y(n_3811)
);

AND2x4_ASAP7_75t_L g3812 ( 
.A(n_3109),
.B(n_3114),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3065),
.Y(n_3813)
);

BUFx3_ASAP7_75t_L g3814 ( 
.A(n_3360),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3119),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_SL g3816 ( 
.A(n_3308),
.B(n_1020),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3071),
.Y(n_3817)
);

OR2x2_ASAP7_75t_L g3818 ( 
.A(n_3027),
.B(n_192),
.Y(n_3818)
);

CKINVDCx8_ASAP7_75t_R g3819 ( 
.A(n_3157),
.Y(n_3819)
);

AOI21xp33_ASAP7_75t_L g3820 ( 
.A1(n_3063),
.A2(n_192),
.B(n_193),
.Y(n_3820)
);

AND2x4_ASAP7_75t_L g3821 ( 
.A(n_3120),
.B(n_192),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_2881),
.B(n_193),
.Y(n_3822)
);

NOR2xp33_ASAP7_75t_R g3823 ( 
.A(n_3444),
.B(n_195),
.Y(n_3823)
);

OR2x6_ASAP7_75t_L g3824 ( 
.A(n_3325),
.B(n_195),
.Y(n_3824)
);

AND2x4_ASAP7_75t_L g3825 ( 
.A(n_3147),
.B(n_196),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3214),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_2998),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_2835),
.B(n_196),
.Y(n_3828)
);

OR2x2_ASAP7_75t_L g3829 ( 
.A(n_3030),
.B(n_2799),
.Y(n_3829)
);

OR2x6_ASAP7_75t_L g3830 ( 
.A(n_3164),
.B(n_196),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_3140),
.B(n_1021),
.Y(n_3831)
);

AOI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_2980),
.A2(n_197),
.B(n_198),
.Y(n_3832)
);

NAND2x1_ASAP7_75t_L g3833 ( 
.A(n_3142),
.B(n_2937),
.Y(n_3833)
);

BUFx4f_ASAP7_75t_L g3834 ( 
.A(n_3425),
.Y(n_3834)
);

BUFx3_ASAP7_75t_L g3835 ( 
.A(n_3378),
.Y(n_3835)
);

BUFx3_ASAP7_75t_L g3836 ( 
.A(n_3379),
.Y(n_3836)
);

INVx1_ASAP7_75t_SL g3837 ( 
.A(n_3437),
.Y(n_3837)
);

BUFx3_ASAP7_75t_L g3838 ( 
.A(n_2908),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3140),
.B(n_1022),
.Y(n_3839)
);

HB1xp67_ASAP7_75t_L g3840 ( 
.A(n_3162),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2837),
.B(n_197),
.Y(n_3841)
);

BUFx3_ASAP7_75t_L g3842 ( 
.A(n_2908),
.Y(n_3842)
);

AND2x4_ASAP7_75t_L g3843 ( 
.A(n_3155),
.B(n_197),
.Y(n_3843)
);

OR2x6_ASAP7_75t_L g3844 ( 
.A(n_3157),
.B(n_198),
.Y(n_3844)
);

BUFx3_ASAP7_75t_L g3845 ( 
.A(n_3296),
.Y(n_3845)
);

AOI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3036),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3217),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_2911),
.B(n_199),
.Y(n_3848)
);

NOR2x1p5_ASAP7_75t_L g3849 ( 
.A(n_2801),
.B(n_199),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3218),
.Y(n_3850)
);

INVx3_ASAP7_75t_SL g3851 ( 
.A(n_3157),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_2837),
.B(n_201),
.Y(n_3852)
);

CKINVDCx8_ASAP7_75t_R g3853 ( 
.A(n_3142),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_3274),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_3854)
);

NAND2x1p5_ASAP7_75t_L g3855 ( 
.A(n_3296),
.B(n_201),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3220),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_SL g3857 ( 
.A(n_3050),
.B(n_1022),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3050),
.B(n_1023),
.Y(n_3858)
);

BUFx3_ASAP7_75t_L g3859 ( 
.A(n_3304),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_2926),
.B(n_202),
.Y(n_3860)
);

CKINVDCx5p33_ASAP7_75t_R g3861 ( 
.A(n_3082),
.Y(n_3861)
);

BUFx2_ASAP7_75t_L g3862 ( 
.A(n_3142),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3222),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_2945),
.B(n_203),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3015),
.Y(n_3865)
);

BUFx2_ASAP7_75t_L g3866 ( 
.A(n_3142),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_L g3867 ( 
.A1(n_3283),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_3867)
);

NOR3xp33_ASAP7_75t_SL g3868 ( 
.A(n_3215),
.B(n_3227),
.C(n_3216),
.Y(n_3868)
);

NOR2x1_ASAP7_75t_L g3869 ( 
.A(n_3266),
.B(n_204),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3010),
.B(n_204),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_2952),
.B(n_205),
.Y(n_3871)
);

OAI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3020),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_3872)
);

A2O1A1Ixp33_ASAP7_75t_L g3873 ( 
.A1(n_3278),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_3873)
);

INVxp67_ASAP7_75t_L g3874 ( 
.A(n_2832),
.Y(n_3874)
);

BUFx4f_ASAP7_75t_SL g3875 ( 
.A(n_2816),
.Y(n_3875)
);

NAND2xp33_ASAP7_75t_SL g3876 ( 
.A(n_3244),
.B(n_209),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3233),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3073),
.Y(n_3878)
);

INVx5_ASAP7_75t_L g3879 ( 
.A(n_2821),
.Y(n_3879)
);

BUFx3_ASAP7_75t_L g3880 ( 
.A(n_3304),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_2889),
.B(n_209),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3125),
.B(n_209),
.Y(n_3882)
);

INVx3_ASAP7_75t_L g3883 ( 
.A(n_3410),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3238),
.Y(n_3884)
);

INVx2_ASAP7_75t_SL g3885 ( 
.A(n_3165),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_2930),
.B(n_210),
.Y(n_3886)
);

NOR2xp33_ASAP7_75t_L g3887 ( 
.A(n_2925),
.B(n_211),
.Y(n_3887)
);

INVx5_ASAP7_75t_L g3888 ( 
.A(n_2821),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3077),
.Y(n_3889)
);

BUFx6f_ASAP7_75t_SL g3890 ( 
.A(n_3156),
.Y(n_3890)
);

HB1xp67_ASAP7_75t_L g3891 ( 
.A(n_3144),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3170),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3239),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3172),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_2864),
.B(n_211),
.Y(n_3895)
);

AOI22xp5_ASAP7_75t_L g3896 ( 
.A1(n_2804),
.A2(n_3034),
.B1(n_2844),
.B2(n_2856),
.Y(n_3896)
);

INVx3_ASAP7_75t_L g3897 ( 
.A(n_3410),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3189),
.Y(n_3898)
);

AND2x4_ASAP7_75t_L g3899 ( 
.A(n_3138),
.B(n_212),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_2846),
.B(n_212),
.Y(n_3900)
);

BUFx2_ASAP7_75t_L g3901 ( 
.A(n_3129),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3415),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3241),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_2865),
.B(n_212),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3245),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3176),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_2955),
.B(n_213),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3247),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3252),
.Y(n_3909)
);

AND2x4_ASAP7_75t_L g3910 ( 
.A(n_3145),
.B(n_213),
.Y(n_3910)
);

BUFx4f_ASAP7_75t_SL g3911 ( 
.A(n_3013),
.Y(n_3911)
);

AOI211xp5_ASAP7_75t_L g3912 ( 
.A1(n_3332),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_3912)
);

INVxp67_ASAP7_75t_SL g3913 ( 
.A(n_3365),
.Y(n_3913)
);

BUFx2_ASAP7_75t_L g3914 ( 
.A(n_3129),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3254),
.Y(n_3915)
);

OR2x6_ASAP7_75t_L g3916 ( 
.A(n_3244),
.B(n_215),
.Y(n_3916)
);

CKINVDCx5p33_ASAP7_75t_R g3917 ( 
.A(n_3344),
.Y(n_3917)
);

INVx4_ASAP7_75t_L g3918 ( 
.A(n_3415),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3359),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3163),
.Y(n_3920)
);

INVx2_ASAP7_75t_SL g3921 ( 
.A(n_3150),
.Y(n_3921)
);

NOR3xp33_ASAP7_75t_SL g3922 ( 
.A(n_3242),
.B(n_216),
.C(n_217),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3166),
.Y(n_3923)
);

BUFx6f_ASAP7_75t_L g3924 ( 
.A(n_3223),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_2969),
.B(n_216),
.Y(n_3925)
);

AND2x4_ASAP7_75t_L g3926 ( 
.A(n_3091),
.B(n_217),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_2859),
.B(n_218),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3262),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_2862),
.B(n_218),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3263),
.Y(n_3930)
);

INVx4_ASAP7_75t_L g3931 ( 
.A(n_3097),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3264),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_R g3933 ( 
.A(n_2937),
.B(n_219),
.Y(n_3933)
);

CKINVDCx16_ASAP7_75t_R g3934 ( 
.A(n_3269),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_SL g3935 ( 
.A(n_3020),
.B(n_1023),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_2868),
.B(n_219),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3171),
.Y(n_3937)
);

AND2x2_ASAP7_75t_SL g3938 ( 
.A(n_3060),
.B(n_220),
.Y(n_3938)
);

OAI221xp5_ASAP7_75t_L g3939 ( 
.A1(n_2870),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.C(n_223),
.Y(n_3939)
);

BUFx4f_ASAP7_75t_L g3940 ( 
.A(n_2821),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3265),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3118),
.B(n_2967),
.Y(n_3942)
);

BUFx6f_ASAP7_75t_L g3943 ( 
.A(n_3346),
.Y(n_3943)
);

OAI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_3197),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_3944)
);

HB1xp67_ASAP7_75t_L g3945 ( 
.A(n_3189),
.Y(n_3945)
);

INVx4_ASAP7_75t_L g3946 ( 
.A(n_2821),
.Y(n_3946)
);

INVx2_ASAP7_75t_L g3947 ( 
.A(n_3382),
.Y(n_3947)
);

AND2x4_ASAP7_75t_L g3948 ( 
.A(n_2890),
.B(n_222),
.Y(n_3948)
);

AOI22xp5_ASAP7_75t_L g3949 ( 
.A1(n_3369),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_2970),
.B(n_223),
.Y(n_3950)
);

HB1xp67_ASAP7_75t_L g3951 ( 
.A(n_3153),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_R g3952 ( 
.A(n_2979),
.B(n_2972),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_R g3953 ( 
.A(n_2979),
.B(n_224),
.Y(n_3953)
);

BUFx2_ASAP7_75t_L g3954 ( 
.A(n_3177),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3267),
.Y(n_3955)
);

CKINVDCx5p33_ASAP7_75t_R g3956 ( 
.A(n_3372),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3131),
.B(n_224),
.Y(n_3957)
);

BUFx12f_ASAP7_75t_L g3958 ( 
.A(n_2979),
.Y(n_3958)
);

HB1xp67_ASAP7_75t_L g3959 ( 
.A(n_3153),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3182),
.Y(n_3960)
);

NOR2x1_ASAP7_75t_L g3961 ( 
.A(n_3269),
.B(n_225),
.Y(n_3961)
);

NOR2xp33_ASAP7_75t_L g3962 ( 
.A(n_2950),
.B(n_225),
.Y(n_3962)
);

BUFx3_ASAP7_75t_L g3963 ( 
.A(n_3384),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3268),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_2834),
.B(n_1024),
.Y(n_3965)
);

HB1xp67_ASAP7_75t_L g3966 ( 
.A(n_3102),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3279),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3149),
.B(n_226),
.Y(n_3968)
);

AND2x6_ASAP7_75t_SL g3969 ( 
.A(n_3390),
.B(n_226),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3182),
.Y(n_3970)
);

AOI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_3396),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_3971)
);

OAI21x1_ASAP7_75t_L g3972 ( 
.A1(n_2920),
.A2(n_227),
.B(n_228),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_L g3973 ( 
.A(n_2963),
.B(n_229),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_2885),
.B(n_229),
.Y(n_3974)
);

INVx4_ASAP7_75t_L g3975 ( 
.A(n_2979),
.Y(n_3975)
);

BUFx3_ASAP7_75t_L g3976 ( 
.A(n_3431),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_2886),
.B(n_230),
.Y(n_3977)
);

BUFx6f_ASAP7_75t_L g3978 ( 
.A(n_3158),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_2887),
.B(n_230),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_2986),
.B(n_3032),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3434),
.B(n_230),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3186),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_2834),
.B(n_1025),
.Y(n_3983)
);

INVx2_ASAP7_75t_SL g3984 ( 
.A(n_2822),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3186),
.Y(n_3985)
);

BUFx6f_ASAP7_75t_L g3986 ( 
.A(n_3158),
.Y(n_3986)
);

AND2x4_ASAP7_75t_L g3987 ( 
.A(n_3051),
.B(n_231),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_2923),
.Y(n_3988)
);

INVx3_ASAP7_75t_L g3989 ( 
.A(n_3154),
.Y(n_3989)
);

OR2x6_ASAP7_75t_SL g3990 ( 
.A(n_3319),
.B(n_231),
.Y(n_3990)
);

AND2x4_ASAP7_75t_L g3991 ( 
.A(n_3054),
.B(n_231),
.Y(n_3991)
);

HB1xp67_ASAP7_75t_L g3992 ( 
.A(n_3104),
.Y(n_3992)
);

AOI22xp5_ASAP7_75t_L g3993 ( 
.A1(n_3001),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_2873),
.B(n_232),
.Y(n_3994)
);

INVx6_ASAP7_75t_L g3995 ( 
.A(n_3158),
.Y(n_3995)
);

AND2x4_ASAP7_75t_L g3996 ( 
.A(n_3281),
.B(n_232),
.Y(n_3996)
);

NOR3xp33_ASAP7_75t_SL g3997 ( 
.A(n_3249),
.B(n_233),
.C(n_234),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_2860),
.B(n_234),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3284),
.Y(n_3999)
);

O2A1O1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_3256),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_2848),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3018),
.Y(n_4002)
);

AOI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_2962),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3285),
.Y(n_4004)
);

HB1xp67_ASAP7_75t_L g4005 ( 
.A(n_3115),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_2922),
.B(n_235),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_2810),
.B(n_236),
.Y(n_4007)
);

BUFx6f_ASAP7_75t_L g4008 ( 
.A(n_3181),
.Y(n_4008)
);

AND2x4_ASAP7_75t_L g4009 ( 
.A(n_3287),
.B(n_237),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3288),
.Y(n_4010)
);

BUFx3_ASAP7_75t_L g4011 ( 
.A(n_3289),
.Y(n_4011)
);

OR2x2_ASAP7_75t_SL g4012 ( 
.A(n_3007),
.B(n_238),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_2898),
.B(n_238),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_3293),
.Y(n_4014)
);

CKINVDCx16_ASAP7_75t_R g4015 ( 
.A(n_3319),
.Y(n_4015)
);

INVx5_ASAP7_75t_L g4016 ( 
.A(n_2929),
.Y(n_4016)
);

OAI22xp5_ASAP7_75t_L g4017 ( 
.A1(n_3203),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_4017)
);

INVx3_ASAP7_75t_L g4018 ( 
.A(n_2929),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3295),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3302),
.Y(n_4020)
);

NOR2xp33_ASAP7_75t_L g4021 ( 
.A(n_2849),
.B(n_239),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3767),
.A2(n_3168),
.B(n_3161),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3577),
.B(n_3094),
.Y(n_4023)
);

OAI21x1_ASAP7_75t_L g4024 ( 
.A1(n_4001),
.A2(n_3173),
.B(n_3161),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3526),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_3583),
.B(n_3211),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3913),
.A2(n_3173),
.B(n_2957),
.Y(n_4027)
);

AND2x4_ASAP7_75t_L g4028 ( 
.A(n_3471),
.B(n_3177),
.Y(n_4028)
);

OAI21x1_ASAP7_75t_SL g4029 ( 
.A1(n_3946),
.A2(n_3408),
.B(n_3184),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3934),
.A2(n_3441),
.B1(n_3411),
.B2(n_3221),
.Y(n_4030)
);

OAI21x1_ASAP7_75t_L g4031 ( 
.A1(n_4018),
.A2(n_3181),
.B(n_3160),
.Y(n_4031)
);

OAI21x1_ASAP7_75t_SL g4032 ( 
.A1(n_3975),
.A2(n_3408),
.B(n_3184),
.Y(n_4032)
);

AOI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3844),
.A2(n_3187),
.B1(n_3074),
.B2(n_3277),
.Y(n_4033)
);

OAI21xp33_ASAP7_75t_L g4034 ( 
.A1(n_3661),
.A2(n_3844),
.B(n_3504),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3707),
.B(n_3230),
.Y(n_4035)
);

INVx6_ASAP7_75t_SL g4036 ( 
.A(n_3503),
.Y(n_4036)
);

AOI21x1_ASAP7_75t_SL g4037 ( 
.A1(n_3587),
.A2(n_3116),
.B(n_3306),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3980),
.B(n_3234),
.Y(n_4038)
);

OAI21x1_ASAP7_75t_L g4039 ( 
.A1(n_3947),
.A2(n_3160),
.B(n_3159),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3587),
.B(n_2858),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_3502),
.A2(n_2957),
.B(n_3057),
.Y(n_4041)
);

OAI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_4015),
.A2(n_3271),
.B1(n_3275),
.B2(n_3260),
.Y(n_4042)
);

INVx4_ASAP7_75t_L g4043 ( 
.A(n_3471),
.Y(n_4043)
);

OAI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3942),
.A2(n_3101),
.B(n_3037),
.Y(n_4044)
);

AOI21xp33_ASAP7_75t_L g4045 ( 
.A1(n_3754),
.A2(n_3420),
.B(n_3414),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3988),
.A2(n_3935),
.B(n_3940),
.Y(n_4046)
);

AND2x2_ASAP7_75t_SL g4047 ( 
.A(n_3517),
.B(n_3297),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3683),
.B(n_3312),
.Y(n_4048)
);

AOI21xp5_ASAP7_75t_L g4049 ( 
.A1(n_3876),
.A2(n_3159),
.B(n_3111),
.Y(n_4049)
);

INVx1_ASAP7_75t_SL g4050 ( 
.A(n_3851),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_4002),
.A2(n_3111),
.B(n_3007),
.Y(n_4051)
);

OAI21x1_ASAP7_75t_SL g4052 ( 
.A1(n_3961),
.A2(n_3329),
.B(n_3251),
.Y(n_4052)
);

AO31x2_ASAP7_75t_L g4053 ( 
.A1(n_3954),
.A2(n_2808),
.A3(n_2999),
.B(n_2833),
.Y(n_4053)
);

AOI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3916),
.A2(n_3021),
.B(n_3105),
.Y(n_4054)
);

OAI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3848),
.A2(n_3040),
.B(n_2903),
.Y(n_4055)
);

OAI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3972),
.A2(n_3128),
.B(n_3178),
.Y(n_4056)
);

NOR2xp33_ASAP7_75t_SL g4057 ( 
.A(n_3819),
.B(n_3391),
.Y(n_4057)
);

AOI21xp5_ASAP7_75t_L g4058 ( 
.A1(n_3916),
.A2(n_3107),
.B(n_2836),
.Y(n_4058)
);

OAI21x1_ASAP7_75t_L g4059 ( 
.A1(n_3833),
.A2(n_3169),
.B(n_3008),
.Y(n_4059)
);

OAI21x1_ASAP7_75t_L g4060 ( 
.A1(n_3989),
.A2(n_2953),
.B(n_3307),
.Y(n_4060)
);

INVx1_ASAP7_75t_SL g4061 ( 
.A(n_3589),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3776),
.B(n_3343),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_3600),
.B(n_3614),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3532),
.Y(n_4064)
);

BUFx6f_ASAP7_75t_L g4065 ( 
.A(n_3457),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3960),
.A2(n_3321),
.B(n_3314),
.Y(n_4066)
);

OAI21x1_ASAP7_75t_L g4067 ( 
.A1(n_3970),
.A2(n_3328),
.B(n_3324),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_3600),
.B(n_3086),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3594),
.A2(n_3055),
.B(n_2958),
.Y(n_4069)
);

AOI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3747),
.A2(n_3336),
.B(n_3333),
.Y(n_4070)
);

BUFx12f_ASAP7_75t_L g4071 ( 
.A(n_3492),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_SL g4072 ( 
.A(n_3471),
.B(n_3391),
.Y(n_4072)
);

AO31x2_ASAP7_75t_L g4073 ( 
.A1(n_3954),
.A2(n_3124),
.A3(n_3113),
.B(n_3337),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3723),
.B(n_3347),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3829),
.B(n_3357),
.Y(n_4075)
);

AND2x4_ASAP7_75t_L g4076 ( 
.A(n_3476),
.B(n_3348),
.Y(n_4076)
);

OAI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3900),
.A2(n_3136),
.B(n_3085),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3476),
.B(n_2929),
.Y(n_4078)
);

NAND3xp33_ASAP7_75t_SL g4079 ( 
.A(n_3570),
.B(n_2936),
.C(n_3235),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3476),
.B(n_2929),
.Y(n_4080)
);

OAI21x1_ASAP7_75t_L g4081 ( 
.A1(n_3982),
.A2(n_3353),
.B(n_3351),
.Y(n_4081)
);

HB1xp67_ASAP7_75t_L g4082 ( 
.A(n_3503),
.Y(n_4082)
);

INVx8_ASAP7_75t_L g4083 ( 
.A(n_3497),
.Y(n_4083)
);

OAI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_3929),
.A2(n_2991),
.B(n_3126),
.Y(n_4084)
);

INVx5_ASAP7_75t_L g4085 ( 
.A(n_3504),
.Y(n_4085)
);

INVx6_ASAP7_75t_L g4086 ( 
.A(n_3568),
.Y(n_4086)
);

OAI21x1_ASAP7_75t_L g4087 ( 
.A1(n_3985),
.A2(n_3356),
.B(n_3354),
.Y(n_4087)
);

AOI21xp33_ASAP7_75t_L g4088 ( 
.A1(n_3891),
.A2(n_3366),
.B(n_3362),
.Y(n_4088)
);

AOI21x1_ASAP7_75t_L g4089 ( 
.A1(n_3862),
.A2(n_2880),
.B(n_3133),
.Y(n_4089)
);

AOI21xp5_ASAP7_75t_L g4090 ( 
.A1(n_3750),
.A2(n_3371),
.B(n_3368),
.Y(n_4090)
);

OAI21x1_ASAP7_75t_L g4091 ( 
.A1(n_3878),
.A2(n_3375),
.B(n_3374),
.Y(n_4091)
);

INVx3_ASAP7_75t_L g4092 ( 
.A(n_3684),
.Y(n_4092)
);

INVx2_ASAP7_75t_SL g4093 ( 
.A(n_3497),
.Y(n_4093)
);

AOI21xp5_ASAP7_75t_L g4094 ( 
.A1(n_3901),
.A2(n_3383),
.B(n_3377),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_3745),
.B(n_2872),
.Y(n_4095)
);

AO31x2_ASAP7_75t_L g4096 ( 
.A1(n_3654),
.A2(n_3388),
.A3(n_3397),
.B(n_3389),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3584),
.B(n_3381),
.Y(n_4097)
);

AO31x2_ASAP7_75t_L g4098 ( 
.A1(n_3654),
.A2(n_3401),
.A3(n_3405),
.B(n_3403),
.Y(n_4098)
);

OAI21xp5_ASAP7_75t_L g4099 ( 
.A1(n_3936),
.A2(n_2901),
.B(n_3315),
.Y(n_4099)
);

OAI21x1_ASAP7_75t_L g4100 ( 
.A1(n_3889),
.A2(n_3407),
.B(n_3406),
.Y(n_4100)
);

INVx3_ASAP7_75t_L g4101 ( 
.A(n_3696),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_3614),
.B(n_3426),
.Y(n_4102)
);

INVx4_ASAP7_75t_L g4103 ( 
.A(n_3489),
.Y(n_4103)
);

OAI21xp5_ASAP7_75t_L g4104 ( 
.A1(n_3831),
.A2(n_3387),
.B(n_3318),
.Y(n_4104)
);

O2A1O1Ixp5_ASAP7_75t_L g4105 ( 
.A1(n_3965),
.A2(n_3392),
.B(n_3422),
.C(n_3394),
.Y(n_4105)
);

OAI21x1_ASAP7_75t_L g4106 ( 
.A1(n_3590),
.A2(n_3438),
.B(n_3430),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_SL g4107 ( 
.A(n_3489),
.B(n_2990),
.Y(n_4107)
);

OA22x2_ASAP7_75t_L g4108 ( 
.A1(n_3601),
.A2(n_3345),
.B1(n_3399),
.B2(n_3237),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3839),
.A2(n_3442),
.B(n_3423),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3901),
.A2(n_3439),
.B(n_3072),
.Y(n_4110)
);

AOI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3914),
.A2(n_3070),
.B(n_3134),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3607),
.B(n_2803),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3537),
.Y(n_4113)
);

OAI21x1_ASAP7_75t_L g4114 ( 
.A1(n_3609),
.A2(n_2990),
.B(n_3080),
.Y(n_4114)
);

BUFx4f_ASAP7_75t_L g4115 ( 
.A(n_3677),
.Y(n_4115)
);

AO31x2_ASAP7_75t_L g4116 ( 
.A1(n_3680),
.A2(n_3092),
.A3(n_3139),
.B(n_3135),
.Y(n_4116)
);

OAI22x1_ASAP7_75t_L g4117 ( 
.A1(n_3784),
.A2(n_3402),
.B1(n_3400),
.B2(n_3185),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3539),
.Y(n_4118)
);

OAI21x1_ASAP7_75t_L g4119 ( 
.A1(n_3617),
.A2(n_3636),
.B(n_3628),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3637),
.B(n_2796),
.Y(n_4120)
);

BUFx8_ASAP7_75t_L g4121 ( 
.A(n_3560),
.Y(n_4121)
);

AND2x4_ASAP7_75t_L g4122 ( 
.A(n_3489),
.B(n_3088),
.Y(n_4122)
);

AOI221xp5_ASAP7_75t_L g4123 ( 
.A1(n_3512),
.A2(n_3045),
.B1(n_2981),
.B2(n_3019),
.C(n_3033),
.Y(n_4123)
);

OAI21x1_ASAP7_75t_SL g4124 ( 
.A1(n_3872),
.A2(n_3174),
.B(n_3183),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3645),
.B(n_3068),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_3914),
.A2(n_3143),
.B(n_3121),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3646),
.B(n_3052),
.Y(n_4127)
);

AOI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_3653),
.A2(n_3061),
.B(n_3059),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3544),
.Y(n_4129)
);

OA22x2_ASAP7_75t_L g4130 ( 
.A1(n_3601),
.A2(n_3446),
.B1(n_3006),
.B2(n_2840),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3663),
.B(n_3064),
.Y(n_4131)
);

A2O1A1Ixp33_ASAP7_75t_L g4132 ( 
.A1(n_3510),
.A2(n_3635),
.B(n_3566),
.C(n_3565),
.Y(n_4132)
);

AOI221x1_ASAP7_75t_L g4133 ( 
.A1(n_3832),
.A2(n_3039),
.B1(n_3038),
.B2(n_2924),
.C(n_2934),
.Y(n_4133)
);

A2O1A1Ixp33_ASAP7_75t_L g4134 ( 
.A1(n_3686),
.A2(n_3167),
.B(n_2951),
.C(n_2940),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3669),
.B(n_3023),
.Y(n_4135)
);

AO22x1_ASAP7_75t_L g4136 ( 
.A1(n_3612),
.A2(n_2990),
.B1(n_3089),
.B2(n_2916),
.Y(n_4136)
);

AO21x2_ASAP7_75t_L g4137 ( 
.A1(n_3952),
.A2(n_2915),
.B(n_3046),
.Y(n_4137)
);

OAI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3886),
.A2(n_3004),
.B(n_3003),
.Y(n_4138)
);

CKINVDCx6p67_ASAP7_75t_R g4139 ( 
.A(n_3462),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_SL g4140 ( 
.A(n_3953),
.B(n_2990),
.Y(n_4140)
);

AOI221xp5_ASAP7_75t_L g4141 ( 
.A1(n_4021),
.A2(n_3047),
.B1(n_2996),
.B2(n_3012),
.C(n_3011),
.Y(n_4141)
);

INVx2_ASAP7_75t_SL g4142 ( 
.A(n_3527),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_3675),
.A2(n_3026),
.B(n_2913),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3546),
.Y(n_4144)
);

INVxp67_ASAP7_75t_L g4145 ( 
.A(n_3677),
.Y(n_4145)
);

NAND2x1p5_ASAP7_75t_L g4146 ( 
.A(n_3576),
.B(n_2907),
.Y(n_4146)
);

OAI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3990),
.A2(n_3630),
.B1(n_3572),
.B2(n_3610),
.Y(n_4147)
);

CKINVDCx20_ASAP7_75t_R g4148 ( 
.A(n_3561),
.Y(n_4148)
);

INVx3_ASAP7_75t_L g4149 ( 
.A(n_3457),
.Y(n_4149)
);

AND2x4_ASAP7_75t_L g4150 ( 
.A(n_3630),
.B(n_240),
.Y(n_4150)
);

BUFx6f_ASAP7_75t_L g4151 ( 
.A(n_3457),
.Y(n_4151)
);

BUFx2_ASAP7_75t_L g4152 ( 
.A(n_3460),
.Y(n_4152)
);

OAI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_3983),
.A2(n_3896),
.B(n_4013),
.Y(n_4153)
);

A2O1A1Ixp33_ASAP7_75t_L g4154 ( 
.A1(n_3758),
.A2(n_3066),
.B(n_2990),
.C(n_242),
.Y(n_4154)
);

OAI21x1_ASAP7_75t_L g4155 ( 
.A1(n_3700),
.A2(n_242),
.B(n_241),
.Y(n_4155)
);

INVxp67_ASAP7_75t_L g4156 ( 
.A(n_3890),
.Y(n_4156)
);

INVx4_ASAP7_75t_L g4157 ( 
.A(n_3481),
.Y(n_4157)
);

OAI21x1_ASAP7_75t_L g4158 ( 
.A1(n_3621),
.A2(n_242),
.B(n_241),
.Y(n_4158)
);

BUFx3_ASAP7_75t_L g4159 ( 
.A(n_3464),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_3451),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3547),
.B(n_240),
.Y(n_4161)
);

AO21x1_ASAP7_75t_L g4162 ( 
.A1(n_3541),
.A2(n_243),
.B(n_244),
.Y(n_4162)
);

INVx3_ASAP7_75t_L g4163 ( 
.A(n_3481),
.Y(n_4163)
);

OAI21x1_ASAP7_75t_L g4164 ( 
.A1(n_3626),
.A2(n_245),
.B(n_244),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3550),
.B(n_243),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_3455),
.Y(n_4166)
);

AOI221xp5_ASAP7_75t_SL g4167 ( 
.A1(n_3725),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.C(n_246),
.Y(n_4167)
);

OAI21x1_ASAP7_75t_L g4168 ( 
.A1(n_3571),
.A2(n_247),
.B(n_246),
.Y(n_4168)
);

NOR2x1_ASAP7_75t_SL g4169 ( 
.A(n_3830),
.B(n_245),
.Y(n_4169)
);

NAND2x1p5_ASAP7_75t_L g4170 ( 
.A(n_3592),
.B(n_246),
.Y(n_4170)
);

INVx2_ASAP7_75t_SL g4171 ( 
.A(n_3481),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3465),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_3558),
.A2(n_247),
.B(n_248),
.Y(n_4173)
);

OAI21x1_ASAP7_75t_L g4174 ( 
.A1(n_3813),
.A2(n_3827),
.B(n_3817),
.Y(n_4174)
);

INVx3_ASAP7_75t_L g4175 ( 
.A(n_3543),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3552),
.B(n_247),
.Y(n_4176)
);

BUFx2_ASAP7_75t_SL g4177 ( 
.A(n_3612),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3554),
.B(n_249),
.Y(n_4178)
);

OA21x2_ASAP7_75t_L g4179 ( 
.A1(n_3680),
.A2(n_3873),
.B(n_4014),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3556),
.B(n_249),
.Y(n_4180)
);

AOI21xp5_ASAP7_75t_L g4181 ( 
.A1(n_3558),
.A2(n_249),
.B(n_250),
.Y(n_4181)
);

AO31x2_ASAP7_75t_L g4182 ( 
.A1(n_3596),
.A2(n_252),
.A3(n_250),
.B(n_251),
.Y(n_4182)
);

A2O1A1Ixp33_ASAP7_75t_L g4183 ( 
.A1(n_3766),
.A2(n_253),
.B(n_250),
.C(n_251),
.Y(n_4183)
);

A2O1A1Ixp33_ASAP7_75t_L g4184 ( 
.A1(n_3769),
.A2(n_254),
.B(n_251),
.C(n_253),
.Y(n_4184)
);

OA22x2_ASAP7_75t_L g4185 ( 
.A1(n_3666),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3572),
.A2(n_255),
.B(n_256),
.Y(n_4186)
);

BUFx6f_ASAP7_75t_L g4187 ( 
.A(n_3543),
.Y(n_4187)
);

OAI21x1_ASAP7_75t_L g4188 ( 
.A1(n_3865),
.A2(n_258),
.B(n_256),
.Y(n_4188)
);

AOI21xp5_ASAP7_75t_L g4189 ( 
.A1(n_3610),
.A2(n_255),
.B(n_259),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_3678),
.B(n_259),
.Y(n_4190)
);

NAND2x1p5_ASAP7_75t_L g4191 ( 
.A(n_3472),
.B(n_260),
.Y(n_4191)
);

AO21x1_ASAP7_75t_L g4192 ( 
.A1(n_3511),
.A2(n_261),
.B(n_262),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3573),
.B(n_3574),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_3620),
.A2(n_261),
.B(n_262),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3575),
.B(n_261),
.Y(n_4195)
);

OAI21x1_ASAP7_75t_L g4196 ( 
.A1(n_3581),
.A2(n_3588),
.B(n_3585),
.Y(n_4196)
);

OAI21x1_ASAP7_75t_L g4197 ( 
.A1(n_3591),
.A2(n_265),
.B(n_264),
.Y(n_4197)
);

NAND3x1_ASAP7_75t_L g4198 ( 
.A(n_3869),
.B(n_263),
.C(n_264),
.Y(n_4198)
);

INVx2_ASAP7_75t_SL g4199 ( 
.A(n_3543),
.Y(n_4199)
);

OAI21x1_ASAP7_75t_L g4200 ( 
.A1(n_3622),
.A2(n_266),
.B(n_265),
.Y(n_4200)
);

AOI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3938),
.A2(n_267),
.B1(n_263),
.B2(n_266),
.Y(n_4201)
);

BUFx12f_ASAP7_75t_L g4202 ( 
.A(n_3597),
.Y(n_4202)
);

OAI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3994),
.A2(n_263),
.B(n_267),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3579),
.B(n_267),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_3469),
.Y(n_4205)
);

AOI21xp5_ASAP7_75t_L g4206 ( 
.A1(n_3620),
.A2(n_268),
.B(n_269),
.Y(n_4206)
);

AOI21xp5_ASAP7_75t_L g4207 ( 
.A1(n_3826),
.A2(n_268),
.B(n_269),
.Y(n_4207)
);

O2A1O1Ixp5_ASAP7_75t_L g4208 ( 
.A1(n_3857),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_4208)
);

CKINVDCx5p33_ASAP7_75t_R g4209 ( 
.A(n_3458),
.Y(n_4209)
);

A2O1A1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_3797),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_4210)
);

HB1xp67_ASAP7_75t_L g4211 ( 
.A(n_3760),
.Y(n_4211)
);

OAI21x1_ASAP7_75t_L g4212 ( 
.A1(n_3638),
.A2(n_273),
.B(n_272),
.Y(n_4212)
);

AOI21x1_ASAP7_75t_L g4213 ( 
.A1(n_3862),
.A2(n_1027),
.B(n_1026),
.Y(n_4213)
);

OAI21xp5_ASAP7_75t_SL g4214 ( 
.A1(n_3506),
.A2(n_279),
.B(n_271),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3580),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_3688),
.B(n_272),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_3847),
.A2(n_273),
.B(n_274),
.Y(n_4217)
);

OAI21x1_ASAP7_75t_SL g4218 ( 
.A1(n_3618),
.A2(n_274),
.B(n_275),
.Y(n_4218)
);

AND3x4_ASAP7_75t_L g4219 ( 
.A(n_3562),
.B(n_275),
.C(n_276),
.Y(n_4219)
);

HB1xp67_ASAP7_75t_L g4220 ( 
.A(n_3764),
.Y(n_4220)
);

OAI21x1_ASAP7_75t_L g4221 ( 
.A1(n_3639),
.A2(n_278),
.B(n_277),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3689),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_3861),
.B(n_276),
.Y(n_4223)
);

OAI21x1_ASAP7_75t_L g4224 ( 
.A1(n_3659),
.A2(n_278),
.B(n_277),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_3640),
.B(n_276),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_3640),
.B(n_277),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3658),
.B(n_279),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3658),
.B(n_279),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_3722),
.B(n_3466),
.Y(n_4229)
);

OAI21x1_ASAP7_75t_L g4230 ( 
.A1(n_3483),
.A2(n_282),
.B(n_281),
.Y(n_4230)
);

OAI21x1_ASAP7_75t_L g4231 ( 
.A1(n_3488),
.A2(n_282),
.B(n_281),
.Y(n_4231)
);

BUFx6f_ASAP7_75t_L g4232 ( 
.A(n_3613),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_3513),
.Y(n_4233)
);

OAI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4007),
.A2(n_280),
.B(n_281),
.Y(n_4234)
);

OAI21xp5_ASAP7_75t_L g4235 ( 
.A1(n_3557),
.A2(n_280),
.B(n_282),
.Y(n_4235)
);

OAI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_3578),
.A2(n_280),
.B(n_283),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_3612),
.B(n_283),
.Y(n_4237)
);

A2O1A1Ixp33_ASAP7_75t_L g4238 ( 
.A1(n_3798),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_4238)
);

OAI21x1_ASAP7_75t_L g4239 ( 
.A1(n_3524),
.A2(n_287),
.B(n_286),
.Y(n_4239)
);

OAI21x1_ASAP7_75t_L g4240 ( 
.A1(n_3540),
.A2(n_287),
.B(n_286),
.Y(n_4240)
);

OAI21x1_ASAP7_75t_L g4241 ( 
.A1(n_3670),
.A2(n_288),
.B(n_287),
.Y(n_4241)
);

BUFx3_ASAP7_75t_L g4242 ( 
.A(n_3482),
.Y(n_4242)
);

OAI21x1_ASAP7_75t_L g4243 ( 
.A1(n_3711),
.A2(n_290),
.B(n_288),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_3721),
.Y(n_4244)
);

OAI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_3473),
.A2(n_290),
.B1(n_284),
.B2(n_288),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3751),
.Y(n_4246)
);

OAI21x1_ASAP7_75t_L g4247 ( 
.A1(n_3775),
.A2(n_292),
.B(n_291),
.Y(n_4247)
);

OAI21x1_ASAP7_75t_L g4248 ( 
.A1(n_3778),
.A2(n_292),
.B(n_291),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_3538),
.B(n_290),
.Y(n_4249)
);

CKINVDCx5p33_ASAP7_75t_R g4250 ( 
.A(n_3564),
.Y(n_4250)
);

OAI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3748),
.A2(n_291),
.B(n_293),
.Y(n_4251)
);

NAND3xp33_ASAP7_75t_L g4252 ( 
.A(n_3529),
.B(n_293),
.C(n_294),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_3593),
.B(n_295),
.Y(n_4253)
);

OAI21x1_ASAP7_75t_L g4254 ( 
.A1(n_3791),
.A2(n_297),
.B(n_296),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_3837),
.B(n_295),
.Y(n_4255)
);

OAI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_3759),
.A2(n_295),
.B(n_296),
.Y(n_4256)
);

INVx6_ASAP7_75t_L g4257 ( 
.A(n_3568),
.Y(n_4257)
);

INVx2_ASAP7_75t_SL g4258 ( 
.A(n_3498),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_SL g4259 ( 
.A(n_3627),
.B(n_297),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_3850),
.B(n_3856),
.Y(n_4260)
);

BUFx3_ASAP7_75t_L g4261 ( 
.A(n_3501),
.Y(n_4261)
);

OAI21x1_ASAP7_75t_L g4262 ( 
.A1(n_3800),
.A2(n_299),
.B(n_298),
.Y(n_4262)
);

AOI221xp5_ASAP7_75t_L g4263 ( 
.A1(n_3454),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.C(n_300),
.Y(n_4263)
);

OA21x2_ASAP7_75t_L g4264 ( 
.A1(n_3863),
.A2(n_3884),
.B(n_3877),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3701),
.Y(n_4265)
);

NAND2x1p5_ASAP7_75t_L g4266 ( 
.A(n_3567),
.B(n_298),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3893),
.B(n_299),
.Y(n_4267)
);

AOI21xp5_ASAP7_75t_L g4268 ( 
.A1(n_3903),
.A2(n_300),
.B(n_301),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3905),
.B(n_301),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_3709),
.Y(n_4270)
);

OAI22x1_ASAP7_75t_L g4271 ( 
.A1(n_3567),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_4271)
);

OAI22xp5_ASAP7_75t_L g4272 ( 
.A1(n_3473),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_4272)
);

OAI21x1_ASAP7_75t_L g4273 ( 
.A1(n_3802),
.A2(n_305),
.B(n_304),
.Y(n_4273)
);

HB1xp67_ASAP7_75t_L g4274 ( 
.A(n_3520),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_3807),
.Y(n_4275)
);

INVx2_ASAP7_75t_SL g4276 ( 
.A(n_3582),
.Y(n_4276)
);

AOI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_3908),
.A2(n_302),
.B(n_304),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_3619),
.B(n_305),
.Y(n_4278)
);

INVx3_ASAP7_75t_L g4279 ( 
.A(n_3719),
.Y(n_4279)
);

A2O1A1Ixp33_ASAP7_75t_L g4280 ( 
.A1(n_3922),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_3909),
.B(n_306),
.Y(n_4281)
);

OAI21x1_ASAP7_75t_L g4282 ( 
.A1(n_3808),
.A2(n_308),
.B(n_307),
.Y(n_4282)
);

INVx1_ASAP7_75t_SL g4283 ( 
.A(n_3736),
.Y(n_4283)
);

AOI21xp33_ASAP7_75t_L g4284 ( 
.A1(n_3898),
.A2(n_306),
.B(n_307),
.Y(n_4284)
);

OAI21x1_ASAP7_75t_L g4285 ( 
.A1(n_3810),
.A2(n_311),
.B(n_310),
.Y(n_4285)
);

AOI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_3615),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_4286)
);

AOI21x1_ASAP7_75t_L g4287 ( 
.A1(n_3866),
.A2(n_3945),
.B(n_3951),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3915),
.B(n_309),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_3928),
.A2(n_311),
.B(n_312),
.Y(n_4289)
);

AOI21x1_ASAP7_75t_L g4290 ( 
.A1(n_3866),
.A2(n_1028),
.B(n_1026),
.Y(n_4290)
);

AO21x1_ASAP7_75t_L g4291 ( 
.A1(n_3511),
.A2(n_312),
.B(n_313),
.Y(n_4291)
);

AOI21xp33_ASAP7_75t_L g4292 ( 
.A1(n_3762),
.A2(n_312),
.B(n_313),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_3930),
.B(n_313),
.Y(n_4293)
);

NAND2x1p5_ASAP7_75t_L g4294 ( 
.A(n_3567),
.B(n_314),
.Y(n_4294)
);

OAI21x1_ASAP7_75t_L g4295 ( 
.A1(n_3920),
.A2(n_316),
.B(n_315),
.Y(n_4295)
);

OAI21x1_ASAP7_75t_SL g4296 ( 
.A1(n_4000),
.A2(n_3718),
.B(n_3702),
.Y(n_4296)
);

AOI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_3932),
.A2(n_314),
.B(n_315),
.Y(n_4297)
);

NAND2x1_ASAP7_75t_L g4298 ( 
.A(n_3719),
.B(n_315),
.Y(n_4298)
);

AOI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_3941),
.A2(n_316),
.B(n_317),
.Y(n_4299)
);

OAI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_3763),
.A2(n_317),
.B(n_318),
.Y(n_4300)
);

A2O1A1Ixp33_ASAP7_75t_L g4301 ( 
.A1(n_3997),
.A2(n_320),
.B(n_317),
.C(n_319),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_3955),
.B(n_320),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_3724),
.Y(n_4303)
);

AOI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_3964),
.A2(n_320),
.B(n_321),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_3967),
.A2(n_321),
.B(n_322),
.Y(n_4305)
);

OAI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_3772),
.A2(n_322),
.B(n_323),
.Y(n_4306)
);

OA21x2_ASAP7_75t_L g4307 ( 
.A1(n_3999),
.A2(n_322),
.B(n_323),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3923),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_3727),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_3729),
.Y(n_4310)
);

OA21x2_ASAP7_75t_L g4311 ( 
.A1(n_4004),
.A2(n_323),
.B(n_324),
.Y(n_4311)
);

OAI21x1_ASAP7_75t_L g4312 ( 
.A1(n_3937),
.A2(n_327),
.B(n_326),
.Y(n_4312)
);

OAI22xp5_ASAP7_75t_L g4313 ( 
.A1(n_3475),
.A2(n_3830),
.B1(n_3783),
.B2(n_3824),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_3892),
.Y(n_4314)
);

AOI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_4010),
.A2(n_325),
.B(n_326),
.Y(n_4315)
);

NOR2xp33_ASAP7_75t_L g4316 ( 
.A(n_3911),
.B(n_325),
.Y(n_4316)
);

BUFx8_ASAP7_75t_L g4317 ( 
.A(n_3605),
.Y(n_4317)
);

AOI21xp5_ASAP7_75t_L g4318 ( 
.A1(n_4019),
.A2(n_327),
.B(n_328),
.Y(n_4318)
);

A2O1A1Ixp33_ASAP7_75t_L g4319 ( 
.A1(n_3912),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_4319)
);

BUFx8_ASAP7_75t_SL g4320 ( 
.A(n_3534),
.Y(n_4320)
);

AOI21xp5_ASAP7_75t_SL g4321 ( 
.A1(n_3516),
.A2(n_328),
.B(n_329),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_3894),
.Y(n_4322)
);

A2O1A1Ixp33_ASAP7_75t_L g4323 ( 
.A1(n_3735),
.A2(n_331),
.B(n_329),
.C(n_330),
.Y(n_4323)
);

AOI211x1_ASAP7_75t_L g4324 ( 
.A1(n_3667),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_4324)
);

AND2x4_ASAP7_75t_L g4325 ( 
.A(n_3627),
.B(n_331),
.Y(n_4325)
);

INVx2_ASAP7_75t_SL g4326 ( 
.A(n_3586),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_3906),
.Y(n_4327)
);

OAI21x1_ASAP7_75t_L g4328 ( 
.A1(n_3456),
.A2(n_334),
.B(n_333),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_3459),
.Y(n_4329)
);

OAI21x1_ASAP7_75t_L g4330 ( 
.A1(n_3470),
.A2(n_334),
.B(n_333),
.Y(n_4330)
);

OAI22xp5_ASAP7_75t_L g4331 ( 
.A1(n_3475),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4020),
.B(n_335),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_3738),
.B(n_335),
.Y(n_4333)
);

NAND2xp33_ASAP7_75t_L g4334 ( 
.A(n_3719),
.B(n_335),
.Y(n_4334)
);

AOI21x1_ASAP7_75t_L g4335 ( 
.A1(n_3959),
.A2(n_1029),
.B(n_1028),
.Y(n_4335)
);

OAI21x1_ASAP7_75t_L g4336 ( 
.A1(n_3474),
.A2(n_338),
.B(n_337),
.Y(n_4336)
);

OAI21x1_ASAP7_75t_L g4337 ( 
.A1(n_3485),
.A2(n_338),
.B(n_337),
.Y(n_4337)
);

OAI21x1_ASAP7_75t_L g4338 ( 
.A1(n_3487),
.A2(n_340),
.B(n_339),
.Y(n_4338)
);

OA21x2_ASAP7_75t_L g4339 ( 
.A1(n_3780),
.A2(n_336),
.B(n_339),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_3741),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_3804),
.A2(n_336),
.B(n_340),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_3804),
.A2(n_336),
.B(n_341),
.Y(n_4342)
);

AND2x4_ASAP7_75t_L g4343 ( 
.A(n_3627),
.B(n_341),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_3742),
.B(n_3756),
.Y(n_4344)
);

OAI21x1_ASAP7_75t_L g4345 ( 
.A1(n_3491),
.A2(n_344),
.B(n_343),
.Y(n_4345)
);

OAI21x1_ASAP7_75t_L g4346 ( 
.A1(n_3493),
.A2(n_345),
.B(n_344),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_3765),
.B(n_342),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3785),
.B(n_3787),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_3788),
.A2(n_342),
.B(n_344),
.Y(n_4349)
);

NOR2x1_ASAP7_75t_L g4350 ( 
.A(n_3666),
.B(n_345),
.Y(n_4350)
);

OAI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_3790),
.A2(n_346),
.B(n_347),
.Y(n_4351)
);

CKINVDCx8_ASAP7_75t_R g4352 ( 
.A(n_3625),
.Y(n_4352)
);

AOI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_3804),
.A2(n_3806),
.B(n_3519),
.Y(n_4353)
);

INVx2_ASAP7_75t_SL g4354 ( 
.A(n_3478),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_3806),
.A2(n_346),
.B(n_347),
.Y(n_4355)
);

INVx2_ASAP7_75t_SL g4356 ( 
.A(n_3478),
.Y(n_4356)
);

OAI21xp5_ASAP7_75t_L g4357 ( 
.A1(n_3795),
.A2(n_346),
.B(n_348),
.Y(n_4357)
);

OAI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3828),
.A2(n_348),
.B(n_349),
.Y(n_4358)
);

AO31x2_ASAP7_75t_L g4359 ( 
.A1(n_3944),
.A2(n_352),
.A3(n_350),
.B(n_351),
.Y(n_4359)
);

OAI21xp5_ASAP7_75t_L g4360 ( 
.A1(n_3841),
.A2(n_350),
.B(n_351),
.Y(n_4360)
);

AOI22xp5_ASAP7_75t_L g4361 ( 
.A1(n_3917),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_4361)
);

INVx3_ASAP7_75t_L g4362 ( 
.A(n_3853),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_SL g4363 ( 
.A(n_3632),
.B(n_352),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_SL g4364 ( 
.A1(n_3516),
.A2(n_353),
.B(n_354),
.Y(n_4364)
);

INVx3_ASAP7_75t_L g4365 ( 
.A(n_3728),
.Y(n_4365)
);

AOI21x1_ASAP7_75t_L g4366 ( 
.A1(n_3716),
.A2(n_1031),
.B(n_1030),
.Y(n_4366)
);

INVx1_ASAP7_75t_SL g4367 ( 
.A(n_3875),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_3794),
.B(n_353),
.Y(n_4368)
);

OAI21x1_ASAP7_75t_L g4369 ( 
.A1(n_3496),
.A2(n_356),
.B(n_355),
.Y(n_4369)
);

AOI21xp5_ASAP7_75t_L g4370 ( 
.A1(n_3806),
.A2(n_354),
.B(n_355),
.Y(n_4370)
);

NAND2xp33_ASAP7_75t_L g4371 ( 
.A(n_3823),
.B(n_356),
.Y(n_4371)
);

OAI22x1_ASAP7_75t_L g4372 ( 
.A1(n_3849),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_4372)
);

OAI21x1_ASAP7_75t_L g4373 ( 
.A1(n_3522),
.A2(n_359),
.B(n_358),
.Y(n_4373)
);

OAI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_3852),
.A2(n_357),
.B(n_359),
.Y(n_4374)
);

AND2x4_ASAP7_75t_L g4375 ( 
.A(n_3632),
.B(n_357),
.Y(n_4375)
);

BUFx6f_ASAP7_75t_L g4376 ( 
.A(n_3613),
.Y(n_4376)
);

NOR2x1_ASAP7_75t_L g4377 ( 
.A(n_3757),
.B(n_359),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_3799),
.B(n_3809),
.Y(n_4378)
);

AND2x4_ASAP7_75t_L g4379 ( 
.A(n_3632),
.B(n_360),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3815),
.Y(n_4380)
);

OAI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_3732),
.A2(n_360),
.B(n_361),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_4011),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_4382)
);

INVx2_ASAP7_75t_SL g4383 ( 
.A(n_3674),
.Y(n_4383)
);

BUFx3_ASAP7_75t_L g4384 ( 
.A(n_3563),
.Y(n_4384)
);

AOI21xp5_ASAP7_75t_L g4385 ( 
.A1(n_3468),
.A2(n_361),
.B(n_362),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_3520),
.Y(n_4386)
);

INVxp67_ASAP7_75t_L g4387 ( 
.A(n_3505),
.Y(n_4387)
);

AOI31xp33_ASAP7_75t_L g4388 ( 
.A1(n_3641),
.A2(n_364),
.A3(n_362),
.B(n_363),
.Y(n_4388)
);

NAND3x1_ASAP7_75t_L g4389 ( 
.A(n_3713),
.B(n_363),
.C(n_364),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_4008),
.A2(n_363),
.B(n_365),
.Y(n_4390)
);

OR2x6_ASAP7_75t_L g4391 ( 
.A(n_3757),
.B(n_365),
.Y(n_4391)
);

OAI21x1_ASAP7_75t_L g4392 ( 
.A1(n_3883),
.A2(n_367),
.B(n_366),
.Y(n_4392)
);

AOI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_4008),
.A2(n_365),
.B(n_366),
.Y(n_4393)
);

INVx3_ASAP7_75t_L g4394 ( 
.A(n_3752),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_3774),
.B(n_367),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_4008),
.A2(n_368),
.B(n_369),
.Y(n_4396)
);

OAI21xp5_ASAP7_75t_L g4397 ( 
.A1(n_3927),
.A2(n_368),
.B(n_369),
.Y(n_4397)
);

AO31x2_ASAP7_75t_L g4398 ( 
.A1(n_4017),
.A2(n_371),
.A3(n_369),
.B(n_370),
.Y(n_4398)
);

AOI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_3450),
.A2(n_370),
.B(n_371),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_3812),
.Y(n_4400)
);

NAND2x1p5_ASAP7_75t_L g4401 ( 
.A(n_3535),
.B(n_370),
.Y(n_4401)
);

AOI21xp5_ASAP7_75t_SL g4402 ( 
.A1(n_3783),
.A2(n_371),
.B(n_372),
.Y(n_4402)
);

A2O1A1Ixp33_ASAP7_75t_L g4403 ( 
.A1(n_3693),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_4403)
);

BUFx3_ASAP7_75t_L g4404 ( 
.A(n_3608),
.Y(n_4404)
);

OAI21x1_ASAP7_75t_L g4405 ( 
.A1(n_3897),
.A2(n_375),
.B(n_374),
.Y(n_4405)
);

OAI21x1_ASAP7_75t_L g4406 ( 
.A1(n_3902),
.A2(n_375),
.B(n_374),
.Y(n_4406)
);

AO31x2_ASAP7_75t_L g4407 ( 
.A1(n_3452),
.A2(n_376),
.A3(n_373),
.B(n_375),
.Y(n_4407)
);

O2A1O1Ixp5_ASAP7_75t_L g4408 ( 
.A1(n_3858),
.A2(n_377),
.B(n_373),
.C(n_376),
.Y(n_4408)
);

AOI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_3956),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_4409)
);

AO31x2_ASAP7_75t_L g4410 ( 
.A1(n_3692),
.A2(n_379),
.A3(n_377),
.B(n_378),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_3740),
.A2(n_379),
.B(n_380),
.Y(n_4411)
);

O2A1O1Ixp5_ASAP7_75t_L g4412 ( 
.A1(n_3705),
.A2(n_382),
.B(n_380),
.C(n_381),
.Y(n_4412)
);

OAI21x1_ASAP7_75t_L g4413 ( 
.A1(n_3792),
.A2(n_383),
.B(n_382),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_3907),
.B(n_381),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_3950),
.B(n_381),
.Y(n_4415)
);

A2O1A1Ixp33_ASAP7_75t_L g4416 ( 
.A1(n_3779),
.A2(n_384),
.B(n_382),
.C(n_383),
.Y(n_4416)
);

OAI21x1_ASAP7_75t_L g4417 ( 
.A1(n_3801),
.A2(n_385),
.B(n_384),
.Y(n_4417)
);

OAI21x1_ASAP7_75t_L g4418 ( 
.A1(n_3777),
.A2(n_386),
.B(n_385),
.Y(n_4418)
);

OAI21xp5_ASAP7_75t_L g4419 ( 
.A1(n_3974),
.A2(n_383),
.B(n_385),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_3812),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4006),
.B(n_386),
.Y(n_4421)
);

OAI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_3977),
.A2(n_386),
.B(n_387),
.Y(n_4422)
);

AND2x6_ASAP7_75t_L g4423 ( 
.A(n_3796),
.B(n_387),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_L g4424 ( 
.A(n_3874),
.B(n_388),
.Y(n_4424)
);

INVx2_ASAP7_75t_SL g4425 ( 
.A(n_3714),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_3998),
.B(n_388),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_3656),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_3803),
.Y(n_4428)
);

OAI21x1_ASAP7_75t_L g4429 ( 
.A1(n_3855),
.A2(n_392),
.B(n_391),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_3895),
.B(n_3904),
.Y(n_4430)
);

HB1xp67_ASAP7_75t_L g4431 ( 
.A(n_3789),
.Y(n_4431)
);

AOI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_3879),
.A2(n_390),
.B(n_391),
.Y(n_4432)
);

AO31x2_ASAP7_75t_L g4433 ( 
.A1(n_3860),
.A2(n_393),
.A3(n_391),
.B(n_392),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_3642),
.B(n_392),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_3768),
.B(n_393),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_3770),
.B(n_394),
.Y(n_4436)
);

OAI21xp33_ASAP7_75t_SL g4437 ( 
.A1(n_3824),
.A2(n_394),
.B(n_395),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_3879),
.A2(n_394),
.B(n_396),
.Y(n_4438)
);

AO21x2_ASAP7_75t_L g4439 ( 
.A1(n_3733),
.A2(n_3816),
.B(n_3734),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3656),
.Y(n_4440)
);

NOR3xp33_ASAP7_75t_L g4441 ( 
.A(n_3650),
.B(n_396),
.C(n_397),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_3699),
.B(n_397),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_3744),
.B(n_397),
.Y(n_4443)
);

AND2x2_ASAP7_75t_SL g4444 ( 
.A(n_3486),
.B(n_398),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_3595),
.Y(n_4445)
);

OAI21x1_ASAP7_75t_L g4446 ( 
.A1(n_3871),
.A2(n_400),
.B(n_399),
.Y(n_4446)
);

CKINVDCx6p67_ASAP7_75t_R g4447 ( 
.A(n_3682),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_3477),
.A2(n_401),
.B(n_399),
.Y(n_4448)
);

OAI21x1_ASAP7_75t_L g4449 ( 
.A1(n_3479),
.A2(n_401),
.B(n_399),
.Y(n_4449)
);

AND2x4_ASAP7_75t_L g4450 ( 
.A(n_3642),
.B(n_398),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_3500),
.B(n_398),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_3595),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_3704),
.Y(n_4453)
);

OR2x2_ASAP7_75t_L g4454 ( 
.A(n_3467),
.B(n_402),
.Y(n_4454)
);

AOI21xp5_ASAP7_75t_L g4455 ( 
.A1(n_3879),
.A2(n_402),
.B(n_403),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_3652),
.Y(n_4456)
);

OAI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_3979),
.A2(n_403),
.B(n_404),
.Y(n_4457)
);

AOI21x1_ASAP7_75t_L g4458 ( 
.A1(n_3716),
.A2(n_1031),
.B(n_1030),
.Y(n_4458)
);

OAI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_3981),
.A2(n_403),
.B(n_404),
.Y(n_4459)
);

OAI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_3962),
.A2(n_404),
.B(n_405),
.Y(n_4460)
);

BUFx6f_ASAP7_75t_L g4461 ( 
.A(n_3613),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_3480),
.A2(n_407),
.B(n_406),
.Y(n_4462)
);

AOI21xp33_ASAP7_75t_L g4463 ( 
.A1(n_3963),
.A2(n_405),
.B(n_406),
.Y(n_4463)
);

OAI21x1_ASAP7_75t_L g4464 ( 
.A1(n_3484),
.A2(n_408),
.B(n_407),
.Y(n_4464)
);

AOI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_3888),
.A2(n_3665),
.B(n_3660),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_3652),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_3888),
.A2(n_405),
.B(n_407),
.Y(n_4467)
);

AOI21x1_ASAP7_75t_L g4468 ( 
.A1(n_3746),
.A2(n_3773),
.B(n_3690),
.Y(n_4468)
);

AOI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_3888),
.A2(n_408),
.B(n_409),
.Y(n_4469)
);

A2O1A1Ixp33_ASAP7_75t_L g4470 ( 
.A1(n_3846),
.A2(n_411),
.B(n_408),
.C(n_409),
.Y(n_4470)
);

OAI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_3739),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_4471)
);

AO21x1_ASAP7_75t_L g4472 ( 
.A1(n_3899),
.A2(n_413),
.B(n_414),
.Y(n_4472)
);

OA22x2_ASAP7_75t_L g4473 ( 
.A1(n_3739),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_4473)
);

BUFx12f_ASAP7_75t_L g4474 ( 
.A(n_3569),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_3704),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_3500),
.B(n_3542),
.Y(n_4476)
);

OAI21x1_ASAP7_75t_L g4477 ( 
.A1(n_3490),
.A2(n_416),
.B(n_415),
.Y(n_4477)
);

AOI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_3660),
.A2(n_414),
.B(n_416),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_3899),
.Y(n_4479)
);

AO31x2_ASAP7_75t_L g4480 ( 
.A1(n_3599),
.A2(n_419),
.A3(n_417),
.B(n_418),
.Y(n_4480)
);

AO31x2_ASAP7_75t_L g4481 ( 
.A1(n_3655),
.A2(n_421),
.A3(n_418),
.B(n_420),
.Y(n_4481)
);

OAI21x1_ASAP7_75t_L g4482 ( 
.A1(n_3495),
.A2(n_422),
.B(n_421),
.Y(n_4482)
);

AO31x2_ASAP7_75t_L g4483 ( 
.A1(n_3507),
.A2(n_422),
.A3(n_418),
.B(n_421),
.Y(n_4483)
);

OAI21x1_ASAP7_75t_L g4484 ( 
.A1(n_3508),
.A2(n_425),
.B(n_424),
.Y(n_4484)
);

OAI21x1_ASAP7_75t_L g4485 ( 
.A1(n_3518),
.A2(n_426),
.B(n_424),
.Y(n_4485)
);

OAI21x1_ASAP7_75t_L g4486 ( 
.A1(n_3521),
.A2(n_426),
.B(n_424),
.Y(n_4486)
);

A2O1A1Ixp33_ASAP7_75t_L g4487 ( 
.A1(n_3973),
.A2(n_427),
.B(n_423),
.C(n_426),
.Y(n_4487)
);

A2O1A1Ixp33_ASAP7_75t_L g4488 ( 
.A1(n_3553),
.A2(n_3993),
.B(n_3881),
.C(n_3948),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_SL g4489 ( 
.A(n_3642),
.B(n_427),
.Y(n_4489)
);

OR2x2_ASAP7_75t_L g4490 ( 
.A(n_3761),
.B(n_427),
.Y(n_4490)
);

INVx3_ASAP7_75t_L g4491 ( 
.A(n_3753),
.Y(n_4491)
);

A2O1A1Ixp33_ASAP7_75t_L g4492 ( 
.A1(n_3948),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_3515),
.B(n_428),
.Y(n_4493)
);

INVxp67_ASAP7_75t_L g4494 ( 
.A(n_3676),
.Y(n_4494)
);

OAI21x1_ASAP7_75t_L g4495 ( 
.A1(n_3525),
.A2(n_431),
.B(n_429),
.Y(n_4495)
);

AOI21x1_ASAP7_75t_L g4496 ( 
.A1(n_3746),
.A2(n_1033),
.B(n_1032),
.Y(n_4496)
);

OAI21xp5_ASAP7_75t_L g4497 ( 
.A1(n_3868),
.A2(n_428),
.B(n_429),
.Y(n_4497)
);

AOI21xp5_ASAP7_75t_L g4498 ( 
.A1(n_3660),
.A2(n_431),
.B(n_432),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_3885),
.B(n_431),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_3840),
.B(n_432),
.Y(n_4500)
);

A2O1A1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_3463),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_4501)
);

AOI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_3665),
.A2(n_433),
.B(n_434),
.Y(n_4502)
);

OAI21xp33_ASAP7_75t_L g4503 ( 
.A1(n_3933),
.A2(n_3598),
.B(n_3528),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3782),
.B(n_434),
.Y(n_4504)
);

OAI21xp33_ASAP7_75t_SL g4505 ( 
.A1(n_3530),
.A2(n_435),
.B(n_436),
.Y(n_4505)
);

AOI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_3665),
.A2(n_435),
.B(n_436),
.Y(n_4506)
);

AOI21xp33_ASAP7_75t_L g4507 ( 
.A1(n_3976),
.A2(n_3921),
.B(n_3499),
.Y(n_4507)
);

BUFx12f_ASAP7_75t_L g4508 ( 
.A(n_3644),
.Y(n_4508)
);

OR2x6_ASAP7_75t_L g4509 ( 
.A(n_3486),
.B(n_436),
.Y(n_4509)
);

OAI21x1_ASAP7_75t_L g4510 ( 
.A1(n_3545),
.A2(n_439),
.B(n_438),
.Y(n_4510)
);

A2O1A1Ixp33_ASAP7_75t_L g4511 ( 
.A1(n_3887),
.A2(n_440),
.B(n_437),
.C(n_439),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_3910),
.Y(n_4512)
);

INVxp67_ASAP7_75t_SL g4513 ( 
.A(n_3966),
.Y(n_4513)
);

INVx1_ASAP7_75t_SL g4514 ( 
.A(n_3694),
.Y(n_4514)
);

AOI21xp33_ASAP7_75t_L g4515 ( 
.A1(n_3461),
.A2(n_437),
.B(n_439),
.Y(n_4515)
);

OAI21x1_ASAP7_75t_L g4516 ( 
.A1(n_3551),
.A2(n_442),
.B(n_441),
.Y(n_4516)
);

AOI21xp5_ASAP7_75t_L g4517 ( 
.A1(n_3668),
.A2(n_437),
.B(n_441),
.Y(n_4517)
);

AOI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_3668),
.A2(n_441),
.B(n_442),
.Y(n_4518)
);

AO31x2_ASAP7_75t_L g4519 ( 
.A1(n_3603),
.A2(n_444),
.A3(n_442),
.B(n_443),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_3992),
.B(n_443),
.Y(n_4520)
);

AND3x4_ASAP7_75t_L g4521 ( 
.A(n_3664),
.B(n_443),
.C(n_444),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_SL g4522 ( 
.A(n_3958),
.B(n_444),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4005),
.B(n_445),
.Y(n_4523)
);

BUFx12f_ASAP7_75t_L g4524 ( 
.A(n_3681),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3712),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_3882),
.B(n_445),
.Y(n_4526)
);

OAI21x1_ASAP7_75t_L g4527 ( 
.A1(n_3604),
.A2(n_448),
.B(n_447),
.Y(n_4527)
);

A2O1A1Ixp33_ASAP7_75t_L g4528 ( 
.A1(n_3926),
.A2(n_3939),
.B(n_3549),
.C(n_3706),
.Y(n_4528)
);

BUFx2_ASAP7_75t_L g4529 ( 
.A(n_3494),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3712),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_3910),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_SL g4532 ( 
.A1(n_3931),
.A2(n_446),
.B(n_448),
.Y(n_4532)
);

AOI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_3668),
.A2(n_446),
.B(n_448),
.Y(n_4533)
);

OAI21x1_ASAP7_75t_SL g4534 ( 
.A1(n_4003),
.A2(n_449),
.B(n_450),
.Y(n_4534)
);

O2A1O1Ixp5_ASAP7_75t_L g4535 ( 
.A1(n_3771),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_4535)
);

OAI21x1_ASAP7_75t_L g4536 ( 
.A1(n_3611),
.A2(n_453),
.B(n_452),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_3818),
.B(n_451),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3814),
.B(n_452),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_3835),
.B(n_453),
.Y(n_4539)
);

OAI21x1_ASAP7_75t_L g4540 ( 
.A1(n_3631),
.A2(n_455),
.B(n_454),
.Y(n_4540)
);

AOI21xp5_ASAP7_75t_L g4541 ( 
.A1(n_3679),
.A2(n_3786),
.B(n_4016),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_3836),
.B(n_453),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_3925),
.B(n_454),
.Y(n_4543)
);

A2O1A1Ixp33_ASAP7_75t_L g4544 ( 
.A1(n_3926),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_SL g4545 ( 
.A(n_3749),
.B(n_3834),
.Y(n_4545)
);

NOR2xp33_ASAP7_75t_SL g4546 ( 
.A(n_3691),
.B(n_457),
.Y(n_4546)
);

OAI22xp5_ASAP7_75t_L g4547 ( 
.A1(n_3542),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_4547)
);

BUFx10_ASAP7_75t_L g4548 ( 
.A(n_3698),
.Y(n_4548)
);

OAI21xp5_ASAP7_75t_L g4549 ( 
.A1(n_3717),
.A2(n_458),
.B(n_459),
.Y(n_4549)
);

OAI21x1_ASAP7_75t_L g4550 ( 
.A1(n_3648),
.A2(n_460),
.B(n_459),
.Y(n_4550)
);

A2O1A1Ixp33_ASAP7_75t_L g4551 ( 
.A1(n_3548),
.A2(n_461),
.B(n_458),
.C(n_460),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_3996),
.B(n_461),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_3679),
.Y(n_4553)
);

BUFx4f_ASAP7_75t_L g4554 ( 
.A(n_3555),
.Y(n_4554)
);

AOI21xp5_ASAP7_75t_L g4555 ( 
.A1(n_3679),
.A2(n_462),
.B(n_463),
.Y(n_4555)
);

AO21x2_ASAP7_75t_L g4556 ( 
.A1(n_3820),
.A2(n_462),
.B(n_463),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_3786),
.A2(n_464),
.B(n_465),
.Y(n_4557)
);

HB1xp67_ASAP7_75t_L g4558 ( 
.A(n_3453),
.Y(n_4558)
);

OAI21x1_ASAP7_75t_SL g4559 ( 
.A1(n_3918),
.A2(n_464),
.B(n_465),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_3996),
.B(n_464),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3730),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_3786),
.A2(n_465),
.B(n_466),
.Y(n_4562)
);

BUFx6f_ASAP7_75t_L g4563 ( 
.A(n_3796),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4009),
.B(n_466),
.Y(n_4564)
);

INVx2_ASAP7_75t_SL g4565 ( 
.A(n_3697),
.Y(n_4565)
);

OAI22xp5_ASAP7_75t_L g4566 ( 
.A1(n_3555),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_4566)
);

OAI21x1_ASAP7_75t_L g4567 ( 
.A1(n_3643),
.A2(n_469),
.B(n_468),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_L g4568 ( 
.A1(n_3647),
.A2(n_470),
.B(n_469),
.Y(n_4568)
);

AOI21xp33_ASAP7_75t_L g4569 ( 
.A1(n_3984),
.A2(n_467),
.B(n_470),
.Y(n_4569)
);

AOI21xp5_ASAP7_75t_L g4570 ( 
.A1(n_4016),
.A2(n_467),
.B(n_471),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4009),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_4016),
.A2(n_472),
.B(n_473),
.Y(n_4572)
);

NOR2xp33_ASAP7_75t_L g4573 ( 
.A(n_3533),
.B(n_472),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_3730),
.Y(n_4574)
);

NAND2x1_ASAP7_75t_L g4575 ( 
.A(n_3773),
.B(n_472),
.Y(n_4575)
);

INVx1_ASAP7_75t_SL g4576 ( 
.A(n_3710),
.Y(n_4576)
);

CKINVDCx5p33_ASAP7_75t_R g4577 ( 
.A(n_3514),
.Y(n_4577)
);

AOI21x1_ASAP7_75t_L g4578 ( 
.A1(n_3535),
.A2(n_1034),
.B(n_1033),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_3864),
.B(n_473),
.Y(n_4579)
);

OAI21x1_ASAP7_75t_L g4580 ( 
.A1(n_3672),
.A2(n_476),
.B(n_474),
.Y(n_4580)
);

AO31x2_ASAP7_75t_L g4581 ( 
.A1(n_3957),
.A2(n_477),
.A3(n_473),
.B(n_474),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_3870),
.B(n_3968),
.Y(n_4582)
);

OAI21x1_ASAP7_75t_L g4583 ( 
.A1(n_3708),
.A2(n_478),
.B(n_477),
.Y(n_4583)
);

OAI21x1_ASAP7_75t_L g4584 ( 
.A1(n_3978),
.A2(n_478),
.B(n_477),
.Y(n_4584)
);

NOR2x1_ASAP7_75t_SL g4585 ( 
.A(n_3978),
.B(n_478),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_3987),
.B(n_474),
.Y(n_4586)
);

INVx3_ASAP7_75t_L g4587 ( 
.A(n_4083),
.Y(n_4587)
);

AOI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_4034),
.A2(n_3726),
.B1(n_3531),
.B2(n_3781),
.Y(n_4588)
);

INVx5_ASAP7_75t_L g4589 ( 
.A(n_4083),
.Y(n_4589)
);

OAI21x1_ASAP7_75t_L g4590 ( 
.A1(n_4039),
.A2(n_3703),
.B(n_3671),
.Y(n_4590)
);

AND2x4_ASAP7_75t_L g4591 ( 
.A(n_4085),
.B(n_3633),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4229),
.B(n_3633),
.Y(n_4592)
);

AO31x2_ASAP7_75t_L g4593 ( 
.A1(n_4022),
.A2(n_3822),
.A3(n_3536),
.B(n_3657),
.Y(n_4593)
);

AO31x2_ASAP7_75t_L g4594 ( 
.A1(n_4049),
.A2(n_3536),
.A3(n_4012),
.B(n_3720),
.Y(n_4594)
);

CKINVDCx5p33_ASAP7_75t_R g4595 ( 
.A(n_4139),
.Y(n_4595)
);

AND2x4_ASAP7_75t_L g4596 ( 
.A(n_4085),
.B(n_3634),
.Y(n_4596)
);

NAND2xp5_ASAP7_75t_L g4597 ( 
.A(n_4260),
.B(n_3634),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4025),
.Y(n_4598)
);

BUFx2_ASAP7_75t_L g4599 ( 
.A(n_4036),
.Y(n_4599)
);

INVx2_ASAP7_75t_SL g4600 ( 
.A(n_4121),
.Y(n_4600)
);

INVx2_ASAP7_75t_SL g4601 ( 
.A(n_4121),
.Y(n_4601)
);

AOI21xp5_ASAP7_75t_L g4602 ( 
.A1(n_4027),
.A2(n_3986),
.B(n_3978),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_4160),
.Y(n_4603)
);

A2O1A1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_4371),
.A2(n_3843),
.B(n_3793),
.C(n_3821),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4064),
.B(n_3843),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_4071),
.Y(n_4606)
);

INVx4_ASAP7_75t_L g4607 ( 
.A(n_4404),
.Y(n_4607)
);

AND2x4_ASAP7_75t_L g4608 ( 
.A(n_4085),
.B(n_3793),
.Y(n_4608)
);

OAI21x1_ASAP7_75t_L g4609 ( 
.A1(n_4024),
.A2(n_3854),
.B(n_3755),
.Y(n_4609)
);

INVx3_ASAP7_75t_L g4610 ( 
.A(n_4157),
.Y(n_4610)
);

NOR2x1_ASAP7_75t_SL g4611 ( 
.A(n_4391),
.B(n_3737),
.Y(n_4611)
);

AOI22xp5_ASAP7_75t_L g4612 ( 
.A1(n_4391),
.A2(n_3559),
.B1(n_3687),
.B2(n_3987),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4113),
.B(n_3811),
.Y(n_4613)
);

O2A1O1Ixp33_ASAP7_75t_SL g4614 ( 
.A1(n_4210),
.A2(n_3731),
.B(n_3971),
.C(n_3949),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4118),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4166),
.Y(n_4616)
);

A2O1A1Ixp33_ASAP7_75t_L g4617 ( 
.A1(n_4554),
.A2(n_3821),
.B(n_3825),
.C(n_3811),
.Y(n_4617)
);

OAI21x1_ASAP7_75t_L g4618 ( 
.A1(n_4031),
.A2(n_3919),
.B(n_3867),
.Y(n_4618)
);

CKINVDCx5p33_ASAP7_75t_R g4619 ( 
.A(n_4317),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4129),
.Y(n_4620)
);

AOI21xp5_ASAP7_75t_L g4621 ( 
.A1(n_4051),
.A2(n_3986),
.B(n_3943),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4144),
.Y(n_4622)
);

AND2x4_ASAP7_75t_L g4623 ( 
.A(n_4157),
.B(n_3825),
.Y(n_4623)
);

CKINVDCx20_ASAP7_75t_R g4624 ( 
.A(n_4148),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4190),
.B(n_3662),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4215),
.Y(n_4626)
);

AOI22xp33_ASAP7_75t_L g4627 ( 
.A1(n_4503),
.A2(n_3805),
.B1(n_3991),
.B2(n_3623),
.Y(n_4627)
);

AOI221xp5_ASAP7_75t_SL g4628 ( 
.A1(n_4388),
.A2(n_3651),
.B1(n_3649),
.B2(n_3969),
.C(n_3943),
.Y(n_4628)
);

OR2x2_ASAP7_75t_L g4629 ( 
.A(n_4211),
.B(n_3695),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4222),
.B(n_3991),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4265),
.Y(n_4631)
);

OAI21x1_ASAP7_75t_L g4632 ( 
.A1(n_4465),
.A2(n_3986),
.B(n_3995),
.Y(n_4632)
);

AOI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4136),
.A2(n_3924),
.B(n_3842),
.Y(n_4633)
);

BUFx10_ASAP7_75t_L g4634 ( 
.A(n_4086),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4270),
.B(n_3673),
.Y(n_4635)
);

OAI21x1_ASAP7_75t_L g4636 ( 
.A1(n_4541),
.A2(n_3995),
.B(n_3924),
.Y(n_4636)
);

OAI21xp5_ASAP7_75t_L g4637 ( 
.A1(n_4535),
.A2(n_3715),
.B(n_3629),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4303),
.B(n_3602),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4309),
.Y(n_4639)
);

NAND2xp33_ASAP7_75t_SL g4640 ( 
.A(n_4313),
.B(n_3606),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4310),
.Y(n_4641)
);

AOI22xp33_ASAP7_75t_L g4642 ( 
.A1(n_4108),
.A2(n_3624),
.B1(n_3743),
.B2(n_3616),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4172),
.Y(n_4643)
);

INVx3_ASAP7_75t_L g4644 ( 
.A(n_4036),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_4317),
.Y(n_4645)
);

OAI22xp5_ASAP7_75t_L g4646 ( 
.A1(n_4115),
.A2(n_3685),
.B1(n_3845),
.B2(n_3838),
.Y(n_4646)
);

INVx4_ASAP7_75t_SL g4647 ( 
.A(n_4423),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4340),
.B(n_4380),
.Y(n_4648)
);

AO31x2_ASAP7_75t_L g4649 ( 
.A1(n_4133),
.A2(n_3880),
.A3(n_3859),
.B(n_481),
.Y(n_4649)
);

INVx3_ASAP7_75t_SL g4650 ( 
.A(n_4447),
.Y(n_4650)
);

AO21x1_ASAP7_75t_L g4651 ( 
.A1(n_4057),
.A2(n_479),
.B(n_480),
.Y(n_4651)
);

NOR3xp33_ASAP7_75t_L g4652 ( 
.A(n_4079),
.B(n_3523),
.C(n_3509),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4193),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4314),
.B(n_479),
.Y(n_4654)
);

OAI21x1_ASAP7_75t_L g4655 ( 
.A1(n_4037),
.A2(n_1053),
.B(n_1042),
.Y(n_4655)
);

AO31x2_ASAP7_75t_L g4656 ( 
.A1(n_4046),
.A2(n_481),
.A3(n_479),
.B(n_480),
.Y(n_4656)
);

OAI22xp5_ASAP7_75t_L g4657 ( 
.A1(n_4201),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_4657)
);

OAI22xp5_ASAP7_75t_L g4658 ( 
.A1(n_4444),
.A2(n_485),
.B1(n_482),
.B2(n_484),
.Y(n_4658)
);

A2O1A1Ixp33_ASAP7_75t_L g4659 ( 
.A1(n_4214),
.A2(n_486),
.B(n_484),
.C(n_485),
.Y(n_4659)
);

BUFx6f_ASAP7_75t_L g4660 ( 
.A(n_4065),
.Y(n_4660)
);

NOR2xp33_ASAP7_75t_L g4661 ( 
.A(n_4082),
.B(n_485),
.Y(n_4661)
);

AOI21xp5_ASAP7_75t_L g4662 ( 
.A1(n_4136),
.A2(n_486),
.B(n_487),
.Y(n_4662)
);

INVx3_ASAP7_75t_L g4663 ( 
.A(n_4142),
.Y(n_4663)
);

AOI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4126),
.A2(n_486),
.B(n_487),
.Y(n_4664)
);

OAI21x1_ASAP7_75t_L g4665 ( 
.A1(n_4060),
.A2(n_1051),
.B(n_1041),
.Y(n_4665)
);

AND2x4_ASAP7_75t_L g4666 ( 
.A(n_4150),
.B(n_4092),
.Y(n_4666)
);

NOR2xp33_ASAP7_75t_L g4667 ( 
.A(n_4145),
.B(n_487),
.Y(n_4667)
);

AOI21xp5_ASAP7_75t_L g4668 ( 
.A1(n_4094),
.A2(n_488),
.B(n_489),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4344),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4322),
.B(n_488),
.Y(n_4670)
);

AOI21xp5_ASAP7_75t_L g4671 ( 
.A1(n_4041),
.A2(n_489),
.B(n_490),
.Y(n_4671)
);

INVx3_ASAP7_75t_L g4672 ( 
.A(n_4548),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4348),
.Y(n_4673)
);

BUFx2_ASAP7_75t_L g4674 ( 
.A(n_4220),
.Y(n_4674)
);

AO31x2_ASAP7_75t_L g4675 ( 
.A1(n_4585),
.A2(n_4353),
.A3(n_4132),
.B(n_4323),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4327),
.B(n_489),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4378),
.B(n_4062),
.Y(n_4677)
);

CKINVDCx20_ASAP7_75t_R g4678 ( 
.A(n_4320),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_4063),
.B(n_490),
.Y(n_4679)
);

AO21x2_ASAP7_75t_L g4680 ( 
.A1(n_4072),
.A2(n_490),
.B(n_491),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4110),
.A2(n_491),
.B(n_492),
.Y(n_4681)
);

AOI21xp5_ASAP7_75t_L g4682 ( 
.A1(n_4029),
.A2(n_491),
.B(n_493),
.Y(n_4682)
);

A2O1A1Ixp33_ASAP7_75t_L g4683 ( 
.A1(n_4437),
.A2(n_495),
.B(n_493),
.C(n_494),
.Y(n_4683)
);

CKINVDCx5p33_ASAP7_75t_R g4684 ( 
.A(n_4250),
.Y(n_4684)
);

OAI21x1_ASAP7_75t_L g4685 ( 
.A1(n_4114),
.A2(n_1051),
.B(n_1040),
.Y(n_4685)
);

AOI221x1_ASAP7_75t_L g4686 ( 
.A1(n_4271),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.C(n_497),
.Y(n_4686)
);

NOR2xp33_ASAP7_75t_L g4687 ( 
.A(n_4061),
.B(n_4367),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4329),
.Y(n_4688)
);

CKINVDCx11_ASAP7_75t_R g4689 ( 
.A(n_4352),
.Y(n_4689)
);

OAI21x1_ASAP7_75t_L g4690 ( 
.A1(n_4059),
.A2(n_1055),
.B(n_1042),
.Y(n_4690)
);

OAI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4412),
.A2(n_494),
.B(n_496),
.Y(n_4691)
);

AO32x2_ASAP7_75t_L g4692 ( 
.A1(n_4147),
.A2(n_498),
.A3(n_496),
.B1(n_497),
.B2(n_499),
.Y(n_4692)
);

NAND3x1_ASAP7_75t_L g4693 ( 
.A(n_4350),
.B(n_497),
.C(n_498),
.Y(n_4693)
);

AOI21xp5_ASAP7_75t_L g4694 ( 
.A1(n_4032),
.A2(n_498),
.B(n_499),
.Y(n_4694)
);

OA21x2_ASAP7_75t_L g4695 ( 
.A1(n_4091),
.A2(n_499),
.B(n_500),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4205),
.Y(n_4696)
);

OAI22xp5_ASAP7_75t_L g4697 ( 
.A1(n_4509),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_4697)
);

INVxp67_ASAP7_75t_L g4698 ( 
.A(n_4431),
.Y(n_4698)
);

O2A1O1Ixp33_ASAP7_75t_L g4699 ( 
.A1(n_4084),
.A2(n_502),
.B(n_500),
.C(n_501),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4476),
.B(n_503),
.Y(n_4700)
);

NOR2xp33_ASAP7_75t_L g4701 ( 
.A(n_4095),
.B(n_503),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4264),
.Y(n_4702)
);

NOR2x1_ASAP7_75t_SL g4703 ( 
.A(n_4177),
.B(n_504),
.Y(n_4703)
);

OAI21xp33_ASAP7_75t_L g4704 ( 
.A1(n_4150),
.A2(n_504),
.B(n_505),
.Y(n_4704)
);

AOI21xp5_ASAP7_75t_L g4705 ( 
.A1(n_4111),
.A2(n_504),
.B(n_505),
.Y(n_4705)
);

OAI21x1_ASAP7_75t_L g4706 ( 
.A1(n_4100),
.A2(n_1046),
.B(n_1036),
.Y(n_4706)
);

AO21x2_ASAP7_75t_L g4707 ( 
.A1(n_4089),
.A2(n_506),
.B(n_507),
.Y(n_4707)
);

NOR2xp67_ASAP7_75t_L g4708 ( 
.A(n_4092),
.B(n_506),
.Y(n_4708)
);

BUFx3_ASAP7_75t_L g4709 ( 
.A(n_4159),
.Y(n_4709)
);

O2A1O1Ixp33_ASAP7_75t_L g4710 ( 
.A1(n_4055),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_4710)
);

A2O1A1Ixp33_ASAP7_75t_L g4711 ( 
.A1(n_4334),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_4711)
);

O2A1O1Ixp33_ASAP7_75t_L g4712 ( 
.A1(n_4238),
.A2(n_510),
.B(n_508),
.C(n_509),
.Y(n_4712)
);

OAI21x1_ASAP7_75t_L g4713 ( 
.A1(n_4066),
.A2(n_1058),
.B(n_1043),
.Y(n_4713)
);

NAND2xp5_ASAP7_75t_L g4714 ( 
.A(n_4513),
.B(n_509),
.Y(n_4714)
);

O2A1O1Ixp33_ASAP7_75t_L g4715 ( 
.A1(n_4280),
.A2(n_513),
.B(n_511),
.C(n_512),
.Y(n_4715)
);

NAND2x1p5_ASAP7_75t_L g4716 ( 
.A(n_4093),
.B(n_511),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4264),
.Y(n_4717)
);

AO31x2_ASAP7_75t_L g4718 ( 
.A1(n_4585),
.A2(n_4553),
.A3(n_4192),
.B(n_4291),
.Y(n_4718)
);

BUFx6f_ASAP7_75t_L g4719 ( 
.A(n_4065),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4233),
.Y(n_4720)
);

AND2x4_ASAP7_75t_L g4721 ( 
.A(n_4101),
.B(n_513),
.Y(n_4721)
);

AO31x2_ASAP7_75t_L g4722 ( 
.A1(n_4162),
.A2(n_515),
.A3(n_512),
.B(n_514),
.Y(n_4722)
);

NAND3x1_ASAP7_75t_L g4723 ( 
.A(n_4377),
.B(n_514),
.C(n_515),
.Y(n_4723)
);

A2O1A1Ixp33_ASAP7_75t_L g4724 ( 
.A1(n_4301),
.A2(n_517),
.B(n_514),
.C(n_516),
.Y(n_4724)
);

AOI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4070),
.A2(n_516),
.B(n_517),
.Y(n_4725)
);

OAI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4105),
.A2(n_516),
.B(n_517),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4244),
.Y(n_4727)
);

A2O1A1Ixp33_ASAP7_75t_L g4728 ( 
.A1(n_4319),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4074),
.B(n_518),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4246),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4275),
.Y(n_4731)
);

CKINVDCx5p33_ASAP7_75t_R g4732 ( 
.A(n_4209),
.Y(n_4732)
);

INVx8_ASAP7_75t_L g4733 ( 
.A(n_4474),
.Y(n_4733)
);

CKINVDCx5p33_ASAP7_75t_R g4734 ( 
.A(n_4508),
.Y(n_4734)
);

AOI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4030),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4308),
.Y(n_4736)
);

BUFx6f_ASAP7_75t_L g4737 ( 
.A(n_4065),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4119),
.Y(n_4738)
);

AOI21xp5_ASAP7_75t_L g4739 ( 
.A1(n_4090),
.A2(n_520),
.B(n_521),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4038),
.B(n_522),
.Y(n_4740)
);

BUFx6f_ASAP7_75t_L g4741 ( 
.A(n_4151),
.Y(n_4741)
);

AOI21x1_ASAP7_75t_L g4742 ( 
.A1(n_4468),
.A2(n_4287),
.B(n_4213),
.Y(n_4742)
);

OA21x2_ASAP7_75t_L g4743 ( 
.A1(n_4067),
.A2(n_522),
.B(n_523),
.Y(n_4743)
);

BUFx10_ASAP7_75t_L g4744 ( 
.A(n_4086),
.Y(n_4744)
);

AOI21xp5_ASAP7_75t_L g4745 ( 
.A1(n_4140),
.A2(n_522),
.B(n_523),
.Y(n_4745)
);

OAI21xp33_ASAP7_75t_L g4746 ( 
.A1(n_4185),
.A2(n_523),
.B(n_524),
.Y(n_4746)
);

OAI21x1_ASAP7_75t_L g4747 ( 
.A1(n_4081),
.A2(n_1056),
.B(n_1039),
.Y(n_4747)
);

AOI22xp33_ASAP7_75t_L g4748 ( 
.A1(n_4042),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_4748)
);

AOI221x1_ASAP7_75t_L g4749 ( 
.A1(n_4402),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.C(n_527),
.Y(n_4749)
);

OAI21x1_ASAP7_75t_L g4750 ( 
.A1(n_4087),
.A2(n_1059),
.B(n_1044),
.Y(n_4750)
);

OR2x2_ASAP7_75t_L g4751 ( 
.A(n_4454),
.B(n_525),
.Y(n_4751)
);

AOI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_4052),
.A2(n_528),
.B(n_529),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4196),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4274),
.B(n_528),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4407),
.Y(n_4755)
);

A2O1A1Ixp33_ASAP7_75t_L g4756 ( 
.A1(n_4058),
.A2(n_531),
.B(n_528),
.C(n_529),
.Y(n_4756)
);

AOI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4128),
.A2(n_529),
.B(n_531),
.Y(n_4757)
);

HB1xp67_ASAP7_75t_L g4758 ( 
.A(n_4386),
.Y(n_4758)
);

OAI21xp5_ASAP7_75t_L g4759 ( 
.A1(n_4208),
.A2(n_531),
.B(n_532),
.Y(n_4759)
);

OAI21x1_ASAP7_75t_L g4760 ( 
.A1(n_4078),
.A2(n_4107),
.B(n_4080),
.Y(n_4760)
);

OR2x2_ASAP7_75t_L g4761 ( 
.A(n_4430),
.B(n_532),
.Y(n_4761)
);

A2O1A1Ixp33_ASAP7_75t_L g4762 ( 
.A1(n_4054),
.A2(n_534),
.B(n_532),
.C(n_533),
.Y(n_4762)
);

OAI21x1_ASAP7_75t_L g4763 ( 
.A1(n_4106),
.A2(n_1056),
.B(n_1039),
.Y(n_4763)
);

CKINVDCx11_ASAP7_75t_R g4764 ( 
.A(n_4548),
.Y(n_4764)
);

INVx1_ASAP7_75t_SL g4765 ( 
.A(n_4514),
.Y(n_4765)
);

O2A1O1Ixp33_ASAP7_75t_L g4766 ( 
.A1(n_4551),
.A2(n_535),
.B(n_533),
.C(n_534),
.Y(n_4766)
);

AOI21x1_ASAP7_75t_L g4767 ( 
.A1(n_4290),
.A2(n_4335),
.B(n_4366),
.Y(n_4767)
);

AOI21xp5_ASAP7_75t_L g4768 ( 
.A1(n_4028),
.A2(n_533),
.B(n_534),
.Y(n_4768)
);

AOI21xp5_ASAP7_75t_L g4769 ( 
.A1(n_4028),
.A2(n_4044),
.B(n_4137),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4407),
.Y(n_4770)
);

A2O1A1Ixp33_ASAP7_75t_L g4771 ( 
.A1(n_4167),
.A2(n_537),
.B(n_535),
.C(n_536),
.Y(n_4771)
);

AOI21x1_ASAP7_75t_SL g4772 ( 
.A1(n_4237),
.A2(n_535),
.B(n_536),
.Y(n_4772)
);

OAI21x1_ASAP7_75t_L g4773 ( 
.A1(n_4056),
.A2(n_1064),
.B(n_1049),
.Y(n_4773)
);

INVx3_ASAP7_75t_L g4774 ( 
.A(n_4101),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_SL g4775 ( 
.A(n_4043),
.B(n_537),
.Y(n_4775)
);

A2O1A1Ixp33_ASAP7_75t_L g4776 ( 
.A1(n_4298),
.A2(n_539),
.B(n_537),
.C(n_538),
.Y(n_4776)
);

INVx5_ASAP7_75t_L g4777 ( 
.A(n_4423),
.Y(n_4777)
);

OAI22x1_ASAP7_75t_L g4778 ( 
.A1(n_4521),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.Y(n_4778)
);

BUFx2_ASAP7_75t_L g4779 ( 
.A(n_4152),
.Y(n_4779)
);

INVx3_ASAP7_75t_SL g4780 ( 
.A(n_4257),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4174),
.Y(n_4781)
);

INVx4_ASAP7_75t_L g4782 ( 
.A(n_4257),
.Y(n_4782)
);

O2A1O1Ixp33_ASAP7_75t_L g4783 ( 
.A1(n_4183),
.A2(n_540),
.B(n_538),
.C(n_539),
.Y(n_4783)
);

O2A1O1Ixp33_ASAP7_75t_L g4784 ( 
.A1(n_4184),
.A2(n_544),
.B(n_541),
.C(n_543),
.Y(n_4784)
);

OAI21x1_ASAP7_75t_L g4785 ( 
.A1(n_4584),
.A2(n_1058),
.B(n_1040),
.Y(n_4785)
);

O2A1O1Ixp33_ASAP7_75t_L g4786 ( 
.A1(n_4138),
.A2(n_544),
.B(n_541),
.C(n_543),
.Y(n_4786)
);

O2A1O1Ixp5_ASAP7_75t_L g4787 ( 
.A1(n_4045),
.A2(n_544),
.B(n_541),
.C(n_543),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4407),
.Y(n_4788)
);

AOI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4153),
.A2(n_545),
.B(n_546),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_4328),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4102),
.B(n_545),
.Y(n_4791)
);

CKINVDCx5p33_ASAP7_75t_R g4792 ( 
.A(n_4524),
.Y(n_4792)
);

HB1xp67_ASAP7_75t_L g4793 ( 
.A(n_4558),
.Y(n_4793)
);

OR2x2_ASAP7_75t_L g4794 ( 
.A(n_4023),
.B(n_545),
.Y(n_4794)
);

INVx3_ASAP7_75t_SL g4795 ( 
.A(n_4577),
.Y(n_4795)
);

INVx3_ASAP7_75t_SL g4796 ( 
.A(n_4050),
.Y(n_4796)
);

BUFx8_ASAP7_75t_L g4797 ( 
.A(n_4202),
.Y(n_4797)
);

OAI21x1_ASAP7_75t_L g4798 ( 
.A1(n_4168),
.A2(n_1067),
.B(n_1050),
.Y(n_4798)
);

OAI22x1_ASAP7_75t_L g4799 ( 
.A1(n_4170),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_4799)
);

NOR2xp33_ASAP7_75t_L g4800 ( 
.A(n_4283),
.B(n_546),
.Y(n_4800)
);

AOI22xp5_ASAP7_75t_L g4801 ( 
.A1(n_4047),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.Y(n_4801)
);

OAI21x1_ASAP7_75t_L g4802 ( 
.A1(n_4188),
.A2(n_1059),
.B(n_1037),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4076),
.A2(n_548),
.B(n_549),
.Y(n_4803)
);

AOI21xp5_ASAP7_75t_L g4804 ( 
.A1(n_4076),
.A2(n_549),
.B(n_550),
.Y(n_4804)
);

AOI21xp5_ASAP7_75t_L g4805 ( 
.A1(n_4179),
.A2(n_550),
.B(n_551),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_4330),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_4179),
.A2(n_550),
.B(n_551),
.Y(n_4807)
);

BUFx10_ASAP7_75t_L g4808 ( 
.A(n_4423),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4433),
.Y(n_4809)
);

AND2x4_ASAP7_75t_L g4810 ( 
.A(n_4169),
.B(n_553),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4433),
.Y(n_4811)
);

O2A1O1Ixp33_ASAP7_75t_L g4812 ( 
.A1(n_4077),
.A2(n_554),
.B(n_552),
.C(n_553),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_4336),
.Y(n_4813)
);

AOI21xp5_ASAP7_75t_L g4814 ( 
.A1(n_4125),
.A2(n_552),
.B(n_553),
.Y(n_4814)
);

OAI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4408),
.A2(n_552),
.B(n_554),
.Y(n_4815)
);

OAI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_4509),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_4816)
);

BUFx6f_ASAP7_75t_L g4817 ( 
.A(n_4151),
.Y(n_4817)
);

INVx5_ASAP7_75t_L g4818 ( 
.A(n_4423),
.Y(n_4818)
);

CKINVDCx11_ASAP7_75t_R g4819 ( 
.A(n_4242),
.Y(n_4819)
);

AOI221x1_ASAP7_75t_L g4820 ( 
.A1(n_4372),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.C(n_558),
.Y(n_4820)
);

INVxp67_ASAP7_75t_SL g4821 ( 
.A(n_4479),
.Y(n_4821)
);

OAI21x1_ASAP7_75t_L g4822 ( 
.A1(n_4197),
.A2(n_1057),
.B(n_1035),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_4253),
.B(n_555),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4075),
.B(n_556),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4433),
.Y(n_4825)
);

AOI21xp5_ASAP7_75t_L g4826 ( 
.A1(n_4127),
.A2(n_557),
.B(n_558),
.Y(n_4826)
);

INVx3_ASAP7_75t_L g4827 ( 
.A(n_4151),
.Y(n_4827)
);

AND2x4_ASAP7_75t_L g4828 ( 
.A(n_4171),
.B(n_560),
.Y(n_4828)
);

AOI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4131),
.A2(n_4134),
.B(n_4528),
.Y(n_4829)
);

AOI21xp5_ASAP7_75t_L g4830 ( 
.A1(n_4088),
.A2(n_559),
.B(n_560),
.Y(n_4830)
);

OR2x2_ASAP7_75t_L g4831 ( 
.A(n_4278),
.B(n_559),
.Y(n_4831)
);

NOR4xp25_ASAP7_75t_L g4832 ( 
.A(n_4198),
.B(n_562),
.C(n_560),
.D(n_561),
.Y(n_4832)
);

OAI21xp5_ASAP7_75t_L g4833 ( 
.A1(n_4488),
.A2(n_561),
.B(n_562),
.Y(n_4833)
);

OAI22x1_ASAP7_75t_L g4834 ( 
.A1(n_4266),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4337),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4481),
.Y(n_4836)
);

AO31x2_ASAP7_75t_L g4837 ( 
.A1(n_4472),
.A2(n_565),
.A3(n_563),
.B(n_564),
.Y(n_4837)
);

BUFx2_ASAP7_75t_L g4838 ( 
.A(n_4232),
.Y(n_4838)
);

INVx2_ASAP7_75t_SL g4839 ( 
.A(n_4261),
.Y(n_4839)
);

CKINVDCx5p33_ASAP7_75t_R g4840 ( 
.A(n_4384),
.Y(n_4840)
);

OAI21x1_ASAP7_75t_L g4841 ( 
.A1(n_4200),
.A2(n_1060),
.B(n_1037),
.Y(n_4841)
);

NOR2xp33_ASAP7_75t_SL g4842 ( 
.A(n_4156),
.B(n_563),
.Y(n_4842)
);

NAND3xp33_ASAP7_75t_SL g4843 ( 
.A(n_4546),
.B(n_564),
.C(n_565),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4481),
.Y(n_4844)
);

AOI21xp5_ASAP7_75t_L g4845 ( 
.A1(n_4445),
.A2(n_566),
.B(n_567),
.Y(n_4845)
);

AOI21xp5_ASAP7_75t_L g4846 ( 
.A1(n_4452),
.A2(n_566),
.B(n_567),
.Y(n_4846)
);

NOR2xp33_ASAP7_75t_L g4847 ( 
.A(n_4576),
.B(n_4223),
.Y(n_4847)
);

AOI221x1_ASAP7_75t_L g4848 ( 
.A1(n_4218),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.C(n_569),
.Y(n_4848)
);

AOI21xp5_ASAP7_75t_L g4849 ( 
.A1(n_4456),
.A2(n_568),
.B(n_569),
.Y(n_4849)
);

BUFx10_ASAP7_75t_L g4850 ( 
.A(n_4187),
.Y(n_4850)
);

A2O1A1Ixp33_ASAP7_75t_L g4851 ( 
.A1(n_4492),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_4851)
);

OR2x2_ASAP7_75t_L g4852 ( 
.A(n_4490),
.B(n_570),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4040),
.B(n_571),
.Y(n_4853)
);

HB1xp67_ASAP7_75t_L g4854 ( 
.A(n_4512),
.Y(n_4854)
);

NOR2xp67_ASAP7_75t_L g4855 ( 
.A(n_4043),
.B(n_571),
.Y(n_4855)
);

OAI21x1_ASAP7_75t_L g4856 ( 
.A1(n_4212),
.A2(n_1065),
.B(n_1043),
.Y(n_4856)
);

OAI21xp5_ASAP7_75t_L g4857 ( 
.A1(n_4154),
.A2(n_572),
.B(n_573),
.Y(n_4857)
);

BUFx12f_ASAP7_75t_L g4858 ( 
.A(n_4294),
.Y(n_4858)
);

A2O1A1Ixp33_ASAP7_75t_L g4859 ( 
.A1(n_4033),
.A2(n_574),
.B(n_572),
.C(n_573),
.Y(n_4859)
);

AOI21xp5_ASAP7_75t_L g4860 ( 
.A1(n_4466),
.A2(n_574),
.B(n_575),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4481),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4048),
.B(n_575),
.Y(n_4862)
);

AOI21xp5_ASAP7_75t_L g4863 ( 
.A1(n_4097),
.A2(n_4363),
.B(n_4259),
.Y(n_4863)
);

AOI21xp5_ASAP7_75t_L g4864 ( 
.A1(n_4434),
.A2(n_575),
.B(n_576),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4400),
.B(n_4427),
.Y(n_4865)
);

AOI21xp5_ASAP7_75t_L g4866 ( 
.A1(n_4489),
.A2(n_576),
.B(n_577),
.Y(n_4866)
);

INVx3_ASAP7_75t_L g4867 ( 
.A(n_4187),
.Y(n_4867)
);

NOR2xp33_ASAP7_75t_L g4868 ( 
.A(n_4316),
.B(n_576),
.Y(n_4868)
);

OR2x2_ASAP7_75t_L g4869 ( 
.A(n_4354),
.B(n_577),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4420),
.Y(n_4870)
);

INVxp67_ASAP7_75t_SL g4871 ( 
.A(n_4531),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4440),
.B(n_577),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4581),
.Y(n_4873)
);

AOI21xp5_ASAP7_75t_L g4874 ( 
.A1(n_4232),
.A2(n_578),
.B(n_579),
.Y(n_4874)
);

BUFx12f_ASAP7_75t_L g4875 ( 
.A(n_4191),
.Y(n_4875)
);

AOI31xp67_ASAP7_75t_L g4876 ( 
.A1(n_4571),
.A2(n_1044),
.A3(n_1045),
.B(n_1038),
.Y(n_4876)
);

AOI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4232),
.A2(n_578),
.B(n_579),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4453),
.B(n_580),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4475),
.B(n_580),
.Y(n_4879)
);

AOI21xp5_ASAP7_75t_L g4880 ( 
.A1(n_4376),
.A2(n_581),
.B(n_582),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4525),
.B(n_4530),
.Y(n_4881)
);

AO31x2_ASAP7_75t_L g4882 ( 
.A1(n_4117),
.A2(n_583),
.A3(n_581),
.B(n_582),
.Y(n_4882)
);

INVx2_ASAP7_75t_SL g4883 ( 
.A(n_4187),
.Y(n_4883)
);

AOI221x1_ASAP7_75t_L g4884 ( 
.A1(n_4321),
.A2(n_584),
.B1(n_582),
.B2(n_583),
.C(n_585),
.Y(n_4884)
);

INVx2_ASAP7_75t_L g4885 ( 
.A(n_4338),
.Y(n_4885)
);

HB1xp67_ASAP7_75t_L g4886 ( 
.A(n_4356),
.Y(n_4886)
);

OAI21x1_ASAP7_75t_L g4887 ( 
.A1(n_4221),
.A2(n_1071),
.B(n_1057),
.Y(n_4887)
);

CKINVDCx5p33_ASAP7_75t_R g4888 ( 
.A(n_4565),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4345),
.Y(n_4889)
);

INVxp67_ASAP7_75t_SL g4890 ( 
.A(n_4376),
.Y(n_4890)
);

AO31x2_ASAP7_75t_L g4891 ( 
.A1(n_4416),
.A2(n_4470),
.A3(n_4403),
.B(n_4103),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4561),
.B(n_583),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4376),
.A2(n_584),
.B(n_585),
.Y(n_4893)
);

INVx3_ASAP7_75t_L g4894 ( 
.A(n_4103),
.Y(n_4894)
);

AOI21xp5_ASAP7_75t_L g4895 ( 
.A1(n_4461),
.A2(n_4069),
.B(n_4143),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4574),
.B(n_584),
.Y(n_4896)
);

AOI221x1_ASAP7_75t_L g4897 ( 
.A1(n_4364),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.C(n_589),
.Y(n_4897)
);

OA21x2_ASAP7_75t_L g4898 ( 
.A1(n_4413),
.A2(n_586),
.B(n_587),
.Y(n_4898)
);

AO21x2_ASAP7_75t_L g4899 ( 
.A1(n_4559),
.A2(n_586),
.B(n_587),
.Y(n_4899)
);

AOI21x1_ASAP7_75t_L g4900 ( 
.A1(n_4458),
.A2(n_4496),
.B(n_4578),
.Y(n_4900)
);

INVx2_ASAP7_75t_SL g4901 ( 
.A(n_4199),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4451),
.B(n_589),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4346),
.Y(n_4903)
);

AO31x2_ASAP7_75t_L g4904 ( 
.A1(n_4432),
.A2(n_591),
.A3(n_589),
.B(n_590),
.Y(n_4904)
);

O2A1O1Ixp33_ASAP7_75t_SL g4905 ( 
.A1(n_4544),
.A2(n_4575),
.B(n_4487),
.C(n_4511),
.Y(n_4905)
);

OAI21x1_ASAP7_75t_L g4906 ( 
.A1(n_4224),
.A2(n_1071),
.B(n_1054),
.Y(n_4906)
);

AO32x2_ASAP7_75t_L g4907 ( 
.A1(n_4471),
.A2(n_592),
.A3(n_590),
.B1(n_591),
.B2(n_593),
.Y(n_4907)
);

OAI22xp5_ASAP7_75t_L g4908 ( 
.A1(n_4473),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_4908)
);

BUFx10_ASAP7_75t_L g4909 ( 
.A(n_4237),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4581),
.Y(n_4910)
);

AOI21xp33_ASAP7_75t_L g4911 ( 
.A1(n_4130),
.A2(n_592),
.B(n_593),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4581),
.Y(n_4912)
);

NAND2x1p5_ASAP7_75t_L g4913 ( 
.A(n_4149),
.B(n_593),
.Y(n_4913)
);

INVx3_ASAP7_75t_L g4914 ( 
.A(n_4149),
.Y(n_4914)
);

NOR2xp67_ASAP7_75t_L g4915 ( 
.A(n_4258),
.B(n_594),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4483),
.Y(n_4916)
);

O2A1O1Ixp33_ASAP7_75t_SL g4917 ( 
.A1(n_4501),
.A2(n_596),
.B(n_594),
.C(n_595),
.Y(n_4917)
);

INVx4_ASAP7_75t_L g4918 ( 
.A(n_4163),
.Y(n_4918)
);

OAI22xp33_ASAP7_75t_L g4919 ( 
.A1(n_4401),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_4919)
);

CKINVDCx20_ASAP7_75t_R g4920 ( 
.A(n_4545),
.Y(n_4920)
);

AOI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4461),
.A2(n_595),
.B(n_597),
.Y(n_4921)
);

OAI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4389),
.A2(n_597),
.B(n_598),
.Y(n_4922)
);

NOR2xp33_ASAP7_75t_L g4923 ( 
.A(n_4068),
.B(n_597),
.Y(n_4923)
);

A2O1A1Ixp33_ASAP7_75t_L g4924 ( 
.A1(n_4429),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4483),
.Y(n_4925)
);

OAI21x1_ASAP7_75t_L g4926 ( 
.A1(n_4230),
.A2(n_1074),
.B(n_1060),
.Y(n_4926)
);

AOI21xp5_ASAP7_75t_L g4927 ( 
.A1(n_4461),
.A2(n_599),
.B(n_600),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4483),
.Y(n_4928)
);

AOI21xp5_ASAP7_75t_L g4929 ( 
.A1(n_4104),
.A2(n_600),
.B(n_601),
.Y(n_4929)
);

BUFx3_ASAP7_75t_L g4930 ( 
.A(n_4529),
.Y(n_4930)
);

O2A1O1Ixp33_ASAP7_75t_L g4931 ( 
.A1(n_4099),
.A2(n_603),
.B(n_601),
.C(n_602),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4387),
.B(n_601),
.Y(n_4932)
);

AOI21xp5_ASAP7_75t_L g4933 ( 
.A1(n_4109),
.A2(n_602),
.B(n_603),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4369),
.Y(n_4934)
);

AOI21x1_ASAP7_75t_L g4935 ( 
.A1(n_4307),
.A2(n_603),
.B(n_604),
.Y(n_4935)
);

INVx4_ASAP7_75t_L g4936 ( 
.A(n_4163),
.Y(n_4936)
);

AOI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4141),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4026),
.A2(n_605),
.B(n_607),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4582),
.B(n_607),
.Y(n_4939)
);

OAI21xp5_ASAP7_75t_SL g4940 ( 
.A1(n_4460),
.A2(n_608),
.B(n_609),
.Y(n_4940)
);

OAI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4235),
.A2(n_608),
.B(n_609),
.Y(n_4941)
);

AOI21xp5_ASAP7_75t_L g4942 ( 
.A1(n_4236),
.A2(n_608),
.B(n_609),
.Y(n_4942)
);

AOI21xp5_ASAP7_75t_L g4943 ( 
.A1(n_4296),
.A2(n_610),
.B(n_611),
.Y(n_4943)
);

INVx2_ASAP7_75t_L g4944 ( 
.A(n_4373),
.Y(n_4944)
);

AO31x2_ASAP7_75t_L g4945 ( 
.A1(n_4438),
.A2(n_612),
.A3(n_610),
.B(n_611),
.Y(n_4945)
);

A2O1A1Ixp33_ASAP7_75t_L g4946 ( 
.A1(n_4497),
.A2(n_612),
.B(n_610),
.C(n_611),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4428),
.B(n_612),
.Y(n_4947)
);

AOI21xp5_ASAP7_75t_L g4948 ( 
.A1(n_4112),
.A2(n_613),
.B(n_614),
.Y(n_4948)
);

O2A1O1Ixp33_ASAP7_75t_SL g4949 ( 
.A1(n_4522),
.A2(n_616),
.B(n_614),
.C(n_615),
.Y(n_4949)
);

AOI21xp5_ASAP7_75t_L g4950 ( 
.A1(n_4120),
.A2(n_615),
.B(n_616),
.Y(n_4950)
);

A2O1A1Ixp33_ASAP7_75t_L g4951 ( 
.A1(n_4155),
.A2(n_618),
.B(n_616),
.C(n_617),
.Y(n_4951)
);

NOR2xp33_ASAP7_75t_L g4952 ( 
.A(n_4494),
.B(n_4421),
.Y(n_4952)
);

AND2x4_ASAP7_75t_L g4953 ( 
.A(n_4175),
.B(n_618),
.Y(n_4953)
);

OR2x2_ASAP7_75t_L g4954 ( 
.A(n_4395),
.B(n_617),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4135),
.B(n_617),
.Y(n_4955)
);

O2A1O1Ixp33_ASAP7_75t_L g4956 ( 
.A1(n_4035),
.A2(n_621),
.B(n_619),
.C(n_620),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_SL g4957 ( 
.A(n_4365),
.B(n_4394),
.Y(n_4957)
);

AOI21x1_ASAP7_75t_L g4958 ( 
.A1(n_4307),
.A2(n_619),
.B(n_621),
.Y(n_4958)
);

AND2x4_ASAP7_75t_L g4959 ( 
.A(n_4175),
.B(n_4279),
.Y(n_4959)
);

AO21x2_ASAP7_75t_L g4960 ( 
.A1(n_4534),
.A2(n_4284),
.B(n_4256),
.Y(n_4960)
);

NOR2x1_ASAP7_75t_R g4961 ( 
.A(n_4177),
.B(n_621),
.Y(n_4961)
);

AO31x2_ASAP7_75t_L g4962 ( 
.A1(n_4455),
.A2(n_624),
.A3(n_622),
.B(n_623),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4339),
.A2(n_625),
.B(n_626),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4339),
.A2(n_625),
.B(n_626),
.Y(n_4964)
);

O2A1O1Ixp33_ASAP7_75t_SL g4965 ( 
.A1(n_4547),
.A2(n_627),
.B(n_625),
.C(n_626),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4519),
.Y(n_4966)
);

INVxp67_ASAP7_75t_SL g4967 ( 
.A(n_4520),
.Y(n_4967)
);

OR2x2_ASAP7_75t_L g4968 ( 
.A(n_4523),
.B(n_627),
.Y(n_4968)
);

NAND3xp33_ASAP7_75t_SL g4969 ( 
.A(n_4219),
.B(n_627),
.C(n_628),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_SL g4970 ( 
.A(n_4365),
.B(n_4394),
.Y(n_4970)
);

OAI21x1_ASAP7_75t_L g4971 ( 
.A1(n_4231),
.A2(n_4240),
.B(n_4239),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4424),
.B(n_629),
.Y(n_4972)
);

AND2x6_ASAP7_75t_L g4973 ( 
.A(n_4325),
.B(n_629),
.Y(n_4973)
);

AOI21x1_ASAP7_75t_L g4974 ( 
.A1(n_4311),
.A2(n_630),
.B(n_632),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4311),
.Y(n_4975)
);

AOI21x1_ASAP7_75t_L g4976 ( 
.A1(n_4325),
.A2(n_630),
.B(n_632),
.Y(n_4976)
);

AO31x2_ASAP7_75t_L g4977 ( 
.A1(n_4467),
.A2(n_633),
.A3(n_630),
.B(n_632),
.Y(n_4977)
);

OAI21x1_ASAP7_75t_L g4978 ( 
.A1(n_4241),
.A2(n_1045),
.B(n_1038),
.Y(n_4978)
);

OAI21xp5_ASAP7_75t_L g4979 ( 
.A1(n_4505),
.A2(n_633),
.B(n_634),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4426),
.B(n_633),
.Y(n_4980)
);

AOI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4123),
.A2(n_4441),
.B1(n_4566),
.B2(n_4286),
.Y(n_4981)
);

INVx1_ASAP7_75t_SL g4982 ( 
.A(n_4383),
.Y(n_4982)
);

AO31x2_ASAP7_75t_L g4983 ( 
.A1(n_4469),
.A2(n_4390),
.A3(n_4396),
.B(n_4393),
.Y(n_4983)
);

OAI21x1_ASAP7_75t_L g4984 ( 
.A1(n_4243),
.A2(n_4248),
.B(n_4247),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_4418),
.Y(n_4985)
);

OAI22xp5_ASAP7_75t_L g4986 ( 
.A1(n_4382),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_4986)
);

AND2x6_ASAP7_75t_SL g4987 ( 
.A(n_4573),
.B(n_635),
.Y(n_4987)
);

OAI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4399),
.A2(n_635),
.B(n_636),
.Y(n_4988)
);

CKINVDCx5p33_ASAP7_75t_R g4989 ( 
.A(n_4425),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4579),
.B(n_637),
.Y(n_4990)
);

AO31x2_ASAP7_75t_L g4991 ( 
.A1(n_4570),
.A2(n_639),
.A3(n_637),
.B(n_638),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4519),
.Y(n_4992)
);

AO22x1_ASAP7_75t_L g4993 ( 
.A1(n_4343),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4519),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4249),
.B(n_639),
.Y(n_4995)
);

INVx1_ASAP7_75t_SL g4996 ( 
.A(n_4276),
.Y(n_4996)
);

AOI21xp5_ASAP7_75t_L g4997 ( 
.A1(n_4124),
.A2(n_4300),
.B(n_4251),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4538),
.B(n_640),
.Y(n_4998)
);

AOI22xp5_ASAP7_75t_L g4999 ( 
.A1(n_4361),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_4999)
);

AOI21xp5_ASAP7_75t_L g5000 ( 
.A1(n_4306),
.A2(n_641),
.B(n_642),
.Y(n_5000)
);

O2A1O1Ixp33_ASAP7_75t_SL g5001 ( 
.A1(n_4463),
.A2(n_644),
.B(n_641),
.C(n_642),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4539),
.B(n_644),
.Y(n_5002)
);

A2O1A1Ixp33_ASAP7_75t_L g5003 ( 
.A1(n_4549),
.A2(n_4459),
.B(n_4351),
.C(n_4357),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4349),
.A2(n_644),
.B(n_645),
.Y(n_5004)
);

OAI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_4385),
.A2(n_645),
.B(n_646),
.Y(n_5005)
);

NAND2xp5_ASAP7_75t_L g5006 ( 
.A(n_4161),
.B(n_646),
.Y(n_5006)
);

OAI21x1_ASAP7_75t_L g5007 ( 
.A1(n_4254),
.A2(n_1054),
.B(n_1049),
.Y(n_5007)
);

OAI21x1_ASAP7_75t_L g5008 ( 
.A1(n_4262),
.A2(n_4282),
.B(n_4273),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4165),
.B(n_4176),
.Y(n_5009)
);

AOI21xp5_ASAP7_75t_L g5010 ( 
.A1(n_4358),
.A2(n_647),
.B(n_648),
.Y(n_5010)
);

OAI21x1_ASAP7_75t_L g5011 ( 
.A1(n_4285),
.A2(n_1066),
.B(n_1061),
.Y(n_5011)
);

AO21x1_ASAP7_75t_L g5012 ( 
.A1(n_4343),
.A2(n_647),
.B(n_649),
.Y(n_5012)
);

AOI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_4360),
.A2(n_649),
.B(n_650),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_L g5014 ( 
.A(n_4178),
.B(n_650),
.Y(n_5014)
);

AO21x1_ASAP7_75t_L g5015 ( 
.A1(n_4375),
.A2(n_650),
.B(n_651),
.Y(n_5015)
);

BUFx3_ASAP7_75t_L g5016 ( 
.A(n_4326),
.Y(n_5016)
);

AOI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_4374),
.A2(n_651),
.B(n_652),
.Y(n_5017)
);

OAI21x1_ASAP7_75t_L g5018 ( 
.A1(n_4295),
.A2(n_4312),
.B(n_4417),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4542),
.B(n_652),
.Y(n_5019)
);

OAI21xp5_ASAP7_75t_L g5020 ( 
.A1(n_4446),
.A2(n_652),
.B(n_653),
.Y(n_5020)
);

OAI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_4448),
.A2(n_653),
.B(n_654),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_L g5022 ( 
.A(n_4180),
.B(n_653),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4480),
.Y(n_5023)
);

A2O1A1Ixp33_ASAP7_75t_L g5024 ( 
.A1(n_4381),
.A2(n_657),
.B(n_655),
.C(n_656),
.Y(n_5024)
);

AOI22xp5_ASAP7_75t_L g5025 ( 
.A1(n_4409),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4480),
.Y(n_5026)
);

NOR2xp67_ASAP7_75t_R g5027 ( 
.A(n_4362),
.B(n_655),
.Y(n_5027)
);

AO31x2_ASAP7_75t_L g5028 ( 
.A1(n_4572),
.A2(n_4272),
.A3(n_4331),
.B(n_4245),
.Y(n_5028)
);

AOI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4439),
.A2(n_656),
.B(n_657),
.Y(n_5029)
);

AOI21x1_ASAP7_75t_L g5030 ( 
.A1(n_4375),
.A2(n_658),
.B(n_659),
.Y(n_5030)
);

CKINVDCx11_ASAP7_75t_R g5031 ( 
.A(n_4563),
.Y(n_5031)
);

OA22x2_ASAP7_75t_L g5032 ( 
.A1(n_4532),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4195),
.B(n_4204),
.Y(n_5033)
);

AOI21xp5_ASAP7_75t_L g5034 ( 
.A1(n_4203),
.A2(n_659),
.B(n_660),
.Y(n_5034)
);

OAI21xp5_ASAP7_75t_L g5035 ( 
.A1(n_4449),
.A2(n_660),
.B(n_661),
.Y(n_5035)
);

INVx2_ASAP7_75t_SL g5036 ( 
.A(n_4563),
.Y(n_5036)
);

BUFx2_ASAP7_75t_L g5037 ( 
.A(n_4563),
.Y(n_5037)
);

NOR2xp33_ASAP7_75t_L g5038 ( 
.A(n_4507),
.B(n_661),
.Y(n_5038)
);

O2A1O1Ixp33_ASAP7_75t_SL g5039 ( 
.A1(n_4515),
.A2(n_4569),
.B(n_4397),
.C(n_4422),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_SL g5040 ( 
.A(n_4491),
.B(n_662),
.Y(n_5040)
);

CKINVDCx5p33_ASAP7_75t_R g5041 ( 
.A(n_4362),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4480),
.Y(n_5042)
);

OAI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4462),
.A2(n_662),
.B(n_663),
.Y(n_5043)
);

AOI22xp5_ASAP7_75t_L g5044 ( 
.A1(n_4263),
.A2(n_665),
.B1(n_662),
.B2(n_664),
.Y(n_5044)
);

INVx2_ASAP7_75t_L g5045 ( 
.A(n_4392),
.Y(n_5045)
);

AO21x2_ASAP7_75t_L g5046 ( 
.A1(n_4234),
.A2(n_664),
.B(n_665),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4216),
.B(n_664),
.Y(n_5047)
);

CKINVDCx5p33_ASAP7_75t_R g5048 ( 
.A(n_4491),
.Y(n_5048)
);

AO31x2_ASAP7_75t_L g5049 ( 
.A1(n_4207),
.A2(n_667),
.A3(n_665),
.B(n_666),
.Y(n_5049)
);

AO32x2_ASAP7_75t_L g5050 ( 
.A1(n_4073),
.A2(n_668),
.A3(n_666),
.B1(n_667),
.B2(n_669),
.Y(n_5050)
);

A2O1A1Ixp33_ASAP7_75t_L g5051 ( 
.A1(n_4419),
.A2(n_668),
.B(n_666),
.C(n_667),
.Y(n_5051)
);

BUFx2_ASAP7_75t_L g5052 ( 
.A(n_4279),
.Y(n_5052)
);

OAI21x1_ASAP7_75t_L g5053 ( 
.A1(n_4405),
.A2(n_1068),
.B(n_1066),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_L g5054 ( 
.A1(n_4406),
.A2(n_1069),
.B(n_1068),
.Y(n_5054)
);

AOI21xp5_ASAP7_75t_L g5055 ( 
.A1(n_4457),
.A2(n_4450),
.B(n_4379),
.Y(n_5055)
);

INVxp67_ASAP7_75t_L g5056 ( 
.A(n_4255),
.Y(n_5056)
);

AO31x2_ASAP7_75t_L g5057 ( 
.A1(n_4217),
.A2(n_670),
.A3(n_668),
.B(n_669),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_SL g5058 ( 
.A(n_4379),
.B(n_669),
.Y(n_5058)
);

INVx3_ASAP7_75t_L g5059 ( 
.A(n_4146),
.Y(n_5059)
);

AOI21xp5_ASAP7_75t_L g5060 ( 
.A1(n_4450),
.A2(n_670),
.B(n_671),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4333),
.Y(n_5061)
);

AND2x4_ASAP7_75t_L g5062 ( 
.A(n_4122),
.B(n_670),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4347),
.B(n_4368),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4598),
.Y(n_5064)
);

INVx8_ASAP7_75t_L g5065 ( 
.A(n_4589),
.Y(n_5065)
);

CKINVDCx6p67_ASAP7_75t_R g5066 ( 
.A(n_4589),
.Y(n_5066)
);

HB1xp67_ASAP7_75t_L g5067 ( 
.A(n_4674),
.Y(n_5067)
);

INVx2_ASAP7_75t_SL g5068 ( 
.A(n_4589),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4677),
.B(n_4073),
.Y(n_5069)
);

AOI22xp33_ASAP7_75t_L g5070 ( 
.A1(n_4973),
.A2(n_4252),
.B1(n_4556),
.B2(n_4292),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_4653),
.B(n_4073),
.Y(n_5071)
);

AOI22xp33_ASAP7_75t_L g5072 ( 
.A1(n_4973),
.A2(n_4969),
.B1(n_5032),
.B2(n_4746),
.Y(n_5072)
);

INVx6_ASAP7_75t_L g5073 ( 
.A(n_4733),
.Y(n_5073)
);

AOI22xp33_ASAP7_75t_L g5074 ( 
.A1(n_4973),
.A2(n_4436),
.B1(n_4435),
.B2(n_4586),
.Y(n_5074)
);

AOI22xp33_ASAP7_75t_L g5075 ( 
.A1(n_4833),
.A2(n_4493),
.B1(n_4442),
.B2(n_4342),
.Y(n_5075)
);

OAI22xp33_ASAP7_75t_L g5076 ( 
.A1(n_4940),
.A2(n_4560),
.B1(n_4564),
.B2(n_4552),
.Y(n_5076)
);

BUFx2_ASAP7_75t_SL g5077 ( 
.A(n_4587),
.Y(n_5077)
);

HB1xp67_ASAP7_75t_L g5078 ( 
.A(n_4793),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_4619),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_4603),
.Y(n_5080)
);

INVx5_ASAP7_75t_L g5081 ( 
.A(n_4733),
.Y(n_5081)
);

BUFx2_ASAP7_75t_SL g5082 ( 
.A(n_4600),
.Y(n_5082)
);

INVx2_ASAP7_75t_SL g5083 ( 
.A(n_4709),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4615),
.Y(n_5084)
);

BUFx12f_ASAP7_75t_L g5085 ( 
.A(n_4764),
.Y(n_5085)
);

CKINVDCx20_ASAP7_75t_R g5086 ( 
.A(n_4678),
.Y(n_5086)
);

INVx2_ASAP7_75t_L g5087 ( 
.A(n_4616),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4620),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4622),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4626),
.Y(n_5090)
);

AOI22xp33_ASAP7_75t_SL g5091 ( 
.A1(n_4611),
.A2(n_4122),
.B1(n_4568),
.B2(n_4567),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4669),
.B(n_4410),
.Y(n_5092)
);

INVx2_ASAP7_75t_L g5093 ( 
.A(n_4643),
.Y(n_5093)
);

AOI22xp33_ASAP7_75t_SL g5094 ( 
.A1(n_4777),
.A2(n_4580),
.B1(n_4226),
.B2(n_4227),
.Y(n_5094)
);

AOI22xp33_ASAP7_75t_L g5095 ( 
.A1(n_4778),
.A2(n_4355),
.B1(n_4370),
.B2(n_4341),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_4696),
.Y(n_5096)
);

AOI22xp33_ASAP7_75t_L g5097 ( 
.A1(n_4704),
.A2(n_4498),
.B1(n_4502),
.B2(n_4478),
.Y(n_5097)
);

OAI22xp33_ASAP7_75t_L g5098 ( 
.A1(n_4588),
.A2(n_4228),
.B1(n_4225),
.B2(n_4173),
.Y(n_5098)
);

BUFx12f_ASAP7_75t_L g5099 ( 
.A(n_4645),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4631),
.Y(n_5100)
);

OAI21xp5_ASAP7_75t_SL g5101 ( 
.A1(n_4612),
.A2(n_4801),
.B(n_5055),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4639),
.Y(n_5102)
);

INVx4_ASAP7_75t_L g5103 ( 
.A(n_4650),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_4641),
.Y(n_5104)
);

OAI22xp33_ASAP7_75t_L g5105 ( 
.A1(n_4777),
.A2(n_4181),
.B1(n_4189),
.B2(n_4186),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4648),
.Y(n_5106)
);

OAI22xp5_ASAP7_75t_L g5107 ( 
.A1(n_4604),
.A2(n_4324),
.B1(n_4194),
.B2(n_4206),
.Y(n_5107)
);

INVx2_ASAP7_75t_SL g5108 ( 
.A(n_4601),
.Y(n_5108)
);

AOI22xp33_ASAP7_75t_L g5109 ( 
.A1(n_4997),
.A2(n_4517),
.B1(n_4518),
.B2(n_4506),
.Y(n_5109)
);

AOI22xp5_ASAP7_75t_L g5110 ( 
.A1(n_4628),
.A2(n_4415),
.B1(n_4414),
.B2(n_4537),
.Y(n_5110)
);

INVxp67_ASAP7_75t_L g5111 ( 
.A(n_4779),
.Y(n_5111)
);

INVx2_ASAP7_75t_SL g5112 ( 
.A(n_5048),
.Y(n_5112)
);

AOI22xp33_ASAP7_75t_SL g5113 ( 
.A1(n_4777),
.A2(n_4158),
.B1(n_4164),
.B2(n_4500),
.Y(n_5113)
);

AOI22xp33_ASAP7_75t_L g5114 ( 
.A1(n_4843),
.A2(n_4533),
.B1(n_4557),
.B2(n_4555),
.Y(n_5114)
);

AOI22xp33_ASAP7_75t_L g5115 ( 
.A1(n_4627),
.A2(n_4562),
.B1(n_4543),
.B2(n_4411),
.Y(n_5115)
);

OR2x2_ASAP7_75t_L g5116 ( 
.A(n_4629),
.B(n_4116),
.Y(n_5116)
);

BUFx4f_ASAP7_75t_SL g5117 ( 
.A(n_4624),
.Y(n_5117)
);

BUFx3_ASAP7_75t_L g5118 ( 
.A(n_4819),
.Y(n_5118)
);

BUFx4f_ASAP7_75t_SL g5119 ( 
.A(n_4797),
.Y(n_5119)
);

BUFx8_ASAP7_75t_L g5120 ( 
.A(n_4599),
.Y(n_5120)
);

BUFx2_ASAP7_75t_L g5121 ( 
.A(n_4930),
.Y(n_5121)
);

BUFx6f_ASAP7_75t_L g5122 ( 
.A(n_5031),
.Y(n_5122)
);

BUFx10_ASAP7_75t_L g5123 ( 
.A(n_4840),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4688),
.Y(n_5124)
);

BUFx12f_ASAP7_75t_L g5125 ( 
.A(n_4689),
.Y(n_5125)
);

BUFx8_ASAP7_75t_L g5126 ( 
.A(n_4858),
.Y(n_5126)
);

INVx2_ASAP7_75t_L g5127 ( 
.A(n_4736),
.Y(n_5127)
);

INVx4_ASAP7_75t_L g5128 ( 
.A(n_4607),
.Y(n_5128)
);

OAI21xp5_ASAP7_75t_SL g5129 ( 
.A1(n_4658),
.A2(n_4277),
.B(n_4268),
.Y(n_5129)
);

CKINVDCx11_ASAP7_75t_R g5130 ( 
.A(n_4796),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_4673),
.Y(n_5131)
);

INVx6_ASAP7_75t_L g5132 ( 
.A(n_4634),
.Y(n_5132)
);

BUFx12f_ASAP7_75t_L g5133 ( 
.A(n_4595),
.Y(n_5133)
);

INVxp33_ASAP7_75t_SL g5134 ( 
.A(n_4961),
.Y(n_5134)
);

BUFx6f_ASAP7_75t_L g5135 ( 
.A(n_5016),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4720),
.Y(n_5136)
);

BUFx8_ASAP7_75t_L g5137 ( 
.A(n_4875),
.Y(n_5137)
);

INVx2_ASAP7_75t_L g5138 ( 
.A(n_4727),
.Y(n_5138)
);

INVx5_ASAP7_75t_L g5139 ( 
.A(n_4744),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_5061),
.B(n_4410),
.Y(n_5140)
);

INVx2_ASAP7_75t_L g5141 ( 
.A(n_4730),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_4731),
.Y(n_5142)
);

AND2x2_ASAP7_75t_L g5143 ( 
.A(n_4592),
.B(n_4116),
.Y(n_5143)
);

CKINVDCx20_ASAP7_75t_R g5144 ( 
.A(n_4606),
.Y(n_5144)
);

INVx2_ASAP7_75t_L g5145 ( 
.A(n_4870),
.Y(n_5145)
);

OAI22xp5_ASAP7_75t_L g5146 ( 
.A1(n_4617),
.A2(n_4297),
.B1(n_4299),
.B2(n_4289),
.Y(n_5146)
);

BUFx3_ASAP7_75t_L g5147 ( 
.A(n_4839),
.Y(n_5147)
);

AOI22xp33_ASAP7_75t_L g5148 ( 
.A1(n_4857),
.A2(n_4526),
.B1(n_4305),
.B2(n_4315),
.Y(n_5148)
);

AOI22xp33_ASAP7_75t_SL g5149 ( 
.A1(n_4818),
.A2(n_4583),
.B1(n_4477),
.B2(n_4482),
.Y(n_5149)
);

OAI22xp33_ASAP7_75t_L g5150 ( 
.A1(n_4818),
.A2(n_4318),
.B1(n_4304),
.B2(n_4267),
.Y(n_5150)
);

AOI22xp33_ASAP7_75t_SL g5151 ( 
.A1(n_4818),
.A2(n_4484),
.B1(n_4485),
.B2(n_4464),
.Y(n_5151)
);

BUFx6f_ASAP7_75t_L g5152 ( 
.A(n_4850),
.Y(n_5152)
);

INVx5_ASAP7_75t_SL g5153 ( 
.A(n_4666),
.Y(n_5153)
);

HB1xp67_ASAP7_75t_L g5154 ( 
.A(n_4758),
.Y(n_5154)
);

CKINVDCx20_ASAP7_75t_R g5155 ( 
.A(n_4684),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4635),
.Y(n_5156)
);

AOI22xp33_ASAP7_75t_L g5157 ( 
.A1(n_4923),
.A2(n_4504),
.B1(n_4269),
.B2(n_4288),
.Y(n_5157)
);

INVx2_ASAP7_75t_L g5158 ( 
.A(n_4702),
.Y(n_5158)
);

BUFx12f_ASAP7_75t_L g5159 ( 
.A(n_4734),
.Y(n_5159)
);

BUFx12f_ASAP7_75t_L g5160 ( 
.A(n_4792),
.Y(n_5160)
);

NAND2x1p5_ASAP7_75t_L g5161 ( 
.A(n_4663),
.B(n_4550),
.Y(n_5161)
);

AOI22xp5_ASAP7_75t_L g5162 ( 
.A1(n_4981),
.A2(n_4281),
.B1(n_4302),
.B2(n_4293),
.Y(n_5162)
);

INVx5_ASAP7_75t_L g5163 ( 
.A(n_4774),
.Y(n_5163)
);

OAI22xp5_ASAP7_75t_SL g5164 ( 
.A1(n_4920),
.A2(n_4499),
.B1(n_4443),
.B2(n_4332),
.Y(n_5164)
);

INVx6_ASAP7_75t_L g5165 ( 
.A(n_4782),
.Y(n_5165)
);

INVx6_ASAP7_75t_L g5166 ( 
.A(n_4909),
.Y(n_5166)
);

BUFx3_ASAP7_75t_L g5167 ( 
.A(n_4888),
.Y(n_5167)
);

INVxp67_ASAP7_75t_L g5168 ( 
.A(n_4915),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_4625),
.B(n_4116),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4881),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_4698),
.Y(n_5171)
);

AOI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_4735),
.A2(n_4816),
.B1(n_4697),
.B2(n_4701),
.Y(n_5172)
);

OAI22xp5_ASAP7_75t_L g5173 ( 
.A1(n_5003),
.A2(n_4182),
.B1(n_4398),
.B2(n_4359),
.Y(n_5173)
);

BUFx4f_ASAP7_75t_L g5174 ( 
.A(n_4780),
.Y(n_5174)
);

INVx2_ASAP7_75t_L g5175 ( 
.A(n_4717),
.Y(n_5175)
);

BUFx10_ASAP7_75t_L g5176 ( 
.A(n_4989),
.Y(n_5176)
);

AOI22xp33_ASAP7_75t_SL g5177 ( 
.A1(n_4703),
.A2(n_4808),
.B1(n_4591),
.B2(n_4608),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_4605),
.Y(n_5178)
);

BUFx4_ASAP7_75t_SL g5179 ( 
.A(n_5041),
.Y(n_5179)
);

AOI22xp33_ASAP7_75t_L g5180 ( 
.A1(n_4829),
.A2(n_4495),
.B1(n_4510),
.B2(n_4486),
.Y(n_5180)
);

CKINVDCx11_ASAP7_75t_R g5181 ( 
.A(n_4795),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_4967),
.B(n_4410),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4613),
.Y(n_5183)
);

BUFx12f_ASAP7_75t_L g5184 ( 
.A(n_4732),
.Y(n_5184)
);

AOI22xp33_ASAP7_75t_L g5185 ( 
.A1(n_5012),
.A2(n_4527),
.B1(n_4536),
.B2(n_4516),
.Y(n_5185)
);

AOI22xp5_ASAP7_75t_L g5186 ( 
.A1(n_4868),
.A2(n_4540),
.B1(n_4182),
.B2(n_4398),
.Y(n_5186)
);

OAI22xp5_ASAP7_75t_L g5187 ( 
.A1(n_4659),
.A2(n_4182),
.B1(n_4398),
.B2(n_4359),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_4630),
.Y(n_5188)
);

INVx6_ASAP7_75t_L g5189 ( 
.A(n_4647),
.Y(n_5189)
);

BUFx10_ASAP7_75t_L g5190 ( 
.A(n_4721),
.Y(n_5190)
);

CKINVDCx11_ASAP7_75t_R g5191 ( 
.A(n_4765),
.Y(n_5191)
);

INVx4_ASAP7_75t_L g5192 ( 
.A(n_4672),
.Y(n_5192)
);

AOI22xp33_ASAP7_75t_L g5193 ( 
.A1(n_5015),
.A2(n_4359),
.B1(n_4053),
.B2(n_4098),
.Y(n_5193)
);

BUFx3_ASAP7_75t_L g5194 ( 
.A(n_4610),
.Y(n_5194)
);

INVxp67_ASAP7_75t_SL g5195 ( 
.A(n_4854),
.Y(n_5195)
);

INVx6_ASAP7_75t_L g5196 ( 
.A(n_4647),
.Y(n_5196)
);

CKINVDCx11_ASAP7_75t_R g5197 ( 
.A(n_4987),
.Y(n_5197)
);

CKINVDCx20_ASAP7_75t_R g5198 ( 
.A(n_4640),
.Y(n_5198)
);

OAI22xp5_ASAP7_75t_L g5199 ( 
.A1(n_4711),
.A2(n_4096),
.B1(n_4098),
.B2(n_4053),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_4638),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4865),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_4886),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4821),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_4838),
.Y(n_5204)
);

INVx6_ASAP7_75t_L g5205 ( 
.A(n_4623),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4871),
.Y(n_5206)
);

BUFx8_ASAP7_75t_L g5207 ( 
.A(n_4810),
.Y(n_5207)
);

OAI22xp33_ASAP7_75t_L g5208 ( 
.A1(n_4842),
.A2(n_4096),
.B1(n_4098),
.B2(n_4053),
.Y(n_5208)
);

AOI22xp33_ASAP7_75t_L g5209 ( 
.A1(n_4911),
.A2(n_4096),
.B1(n_673),
.B2(n_671),
.Y(n_5209)
);

INVx2_ASAP7_75t_SL g5210 ( 
.A(n_4996),
.Y(n_5210)
);

AOI22xp33_ASAP7_75t_SL g5211 ( 
.A1(n_4596),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_5211)
);

AOI22xp33_ASAP7_75t_L g5212 ( 
.A1(n_4922),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_4838),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_4975),
.Y(n_5214)
);

AOI22xp33_ASAP7_75t_SL g5215 ( 
.A1(n_5062),
.A2(n_676),
.B1(n_674),
.B2(n_675),
.Y(n_5215)
);

CKINVDCx11_ASAP7_75t_R g5216 ( 
.A(n_4982),
.Y(n_5216)
);

BUFx8_ASAP7_75t_SL g5217 ( 
.A(n_4644),
.Y(n_5217)
);

BUFx12f_ASAP7_75t_L g5218 ( 
.A(n_4716),
.Y(n_5218)
);

AOI22xp33_ASAP7_75t_SL g5219 ( 
.A1(n_5052),
.A2(n_677),
.B1(n_675),
.B2(n_676),
.Y(n_5219)
);

BUFx12f_ASAP7_75t_L g5220 ( 
.A(n_4831),
.Y(n_5220)
);

AOI22xp5_ASAP7_75t_L g5221 ( 
.A1(n_4652),
.A2(n_4657),
.B1(n_4748),
.B2(n_4919),
.Y(n_5221)
);

AOI22xp33_ASAP7_75t_L g5222 ( 
.A1(n_4941),
.A2(n_678),
.B1(n_675),
.B2(n_677),
.Y(n_5222)
);

BUFx12f_ASAP7_75t_L g5223 ( 
.A(n_4828),
.Y(n_5223)
);

INVx1_ASAP7_75t_SL g5224 ( 
.A(n_5037),
.Y(n_5224)
);

INVx8_ASAP7_75t_L g5225 ( 
.A(n_4959),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4714),
.Y(n_5226)
);

CKINVDCx20_ASAP7_75t_R g5227 ( 
.A(n_4687),
.Y(n_5227)
);

INVx8_ASAP7_75t_L g5228 ( 
.A(n_5059),
.Y(n_5228)
);

INVx2_ASAP7_75t_L g5229 ( 
.A(n_4660),
.Y(n_5229)
);

AOI22xp33_ASAP7_75t_L g5230 ( 
.A1(n_4651),
.A2(n_679),
.B1(n_677),
.B2(n_678),
.Y(n_5230)
);

OAI22xp5_ASAP7_75t_L g5231 ( 
.A1(n_4708),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_4800),
.Y(n_5232)
);

BUFx2_ASAP7_75t_SL g5233 ( 
.A(n_4855),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_4755),
.Y(n_5234)
);

INVx2_ASAP7_75t_L g5235 ( 
.A(n_4660),
.Y(n_5235)
);

OAI22xp33_ASAP7_75t_L g5236 ( 
.A1(n_4884),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_4894),
.Y(n_5237)
);

INVx6_ASAP7_75t_L g5238 ( 
.A(n_4918),
.Y(n_5238)
);

BUFx2_ASAP7_75t_L g5239 ( 
.A(n_4936),
.Y(n_5239)
);

AND2x4_ASAP7_75t_SL g5240 ( 
.A(n_4953),
.B(n_681),
.Y(n_5240)
);

INVx1_ASAP7_75t_SL g5241 ( 
.A(n_4823),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_L g5242 ( 
.A(n_4597),
.B(n_683),
.Y(n_5242)
);

OAI22xp5_ASAP7_75t_L g5243 ( 
.A1(n_4723),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_4719),
.Y(n_5244)
);

AOI22xp33_ASAP7_75t_L g5245 ( 
.A1(n_4960),
.A2(n_686),
.B1(n_683),
.B2(n_685),
.Y(n_5245)
);

INVx5_ASAP7_75t_L g5246 ( 
.A(n_4719),
.Y(n_5246)
);

CKINVDCx11_ASAP7_75t_R g5247 ( 
.A(n_4646),
.Y(n_5247)
);

BUFx6f_ASAP7_75t_L g5248 ( 
.A(n_4737),
.Y(n_5248)
);

INVx8_ASAP7_75t_L g5249 ( 
.A(n_4737),
.Y(n_5249)
);

INVx2_ASAP7_75t_SL g5250 ( 
.A(n_4901),
.Y(n_5250)
);

AOI22xp5_ASAP7_75t_L g5251 ( 
.A1(n_5038),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.Y(n_5251)
);

AOI22xp33_ASAP7_75t_L g5252 ( 
.A1(n_4942),
.A2(n_4799),
.B1(n_4972),
.B2(n_4899),
.Y(n_5252)
);

INVx6_ASAP7_75t_L g5253 ( 
.A(n_4741),
.Y(n_5253)
);

CKINVDCx20_ASAP7_75t_R g5254 ( 
.A(n_4902),
.Y(n_5254)
);

INVx6_ASAP7_75t_SL g5255 ( 
.A(n_4642),
.Y(n_5255)
);

CKINVDCx5p33_ASAP7_75t_R g5256 ( 
.A(n_4847),
.Y(n_5256)
);

OAI22xp5_ASAP7_75t_L g5257 ( 
.A1(n_4693),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.Y(n_5257)
);

BUFx2_ASAP7_75t_L g5258 ( 
.A(n_4741),
.Y(n_5258)
);

CKINVDCx6p67_ASAP7_75t_R g5259 ( 
.A(n_4834),
.Y(n_5259)
);

AOI22xp33_ASAP7_75t_L g5260 ( 
.A1(n_4791),
.A2(n_689),
.B1(n_687),
.B2(n_688),
.Y(n_5260)
);

INVx5_ASAP7_75t_L g5261 ( 
.A(n_4817),
.Y(n_5261)
);

OAI22xp33_ASAP7_75t_L g5262 ( 
.A1(n_4897),
.A2(n_691),
.B1(n_689),
.B2(n_690),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4770),
.Y(n_5263)
);

INVx2_ASAP7_75t_L g5264 ( 
.A(n_4817),
.Y(n_5264)
);

INVx1_ASAP7_75t_SL g5265 ( 
.A(n_4794),
.Y(n_5265)
);

INVx2_ASAP7_75t_L g5266 ( 
.A(n_5036),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_4788),
.Y(n_5267)
);

CKINVDCx20_ASAP7_75t_R g5268 ( 
.A(n_4679),
.Y(n_5268)
);

OAI22xp33_ASAP7_75t_L g5269 ( 
.A1(n_4749),
.A2(n_693),
.B1(n_690),
.B2(n_692),
.Y(n_5269)
);

INVx4_ASAP7_75t_L g5270 ( 
.A(n_4827),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_4883),
.Y(n_5271)
);

AOI22xp33_ASAP7_75t_SL g5272 ( 
.A1(n_4908),
.A2(n_693),
.B1(n_690),
.B2(n_692),
.Y(n_5272)
);

INVx2_ASAP7_75t_SL g5273 ( 
.A(n_4957),
.Y(n_5273)
);

HB1xp67_ASAP7_75t_L g5274 ( 
.A(n_4970),
.Y(n_5274)
);

OAI22xp5_ASAP7_75t_SL g5275 ( 
.A1(n_4832),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_5056),
.B(n_4729),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_4952),
.B(n_694),
.Y(n_5277)
);

AOI22xp33_ASAP7_75t_SL g5278 ( 
.A1(n_4913),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4809),
.Y(n_5279)
);

BUFx12f_ASAP7_75t_L g5280 ( 
.A(n_4751),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4811),
.Y(n_5281)
);

OAI22xp33_ASAP7_75t_L g5282 ( 
.A1(n_4820),
.A2(n_4848),
.B1(n_4686),
.B2(n_5058),
.Y(n_5282)
);

CKINVDCx11_ASAP7_75t_R g5283 ( 
.A(n_5045),
.Y(n_5283)
);

BUFx10_ASAP7_75t_L g5284 ( 
.A(n_4661),
.Y(n_5284)
);

BUFx12f_ASAP7_75t_L g5285 ( 
.A(n_4852),
.Y(n_5285)
);

AOI22xp5_ASAP7_75t_L g5286 ( 
.A1(n_5044),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_5286)
);

BUFx3_ASAP7_75t_L g5287 ( 
.A(n_4867),
.Y(n_5287)
);

OAI22xp33_ASAP7_75t_L g5288 ( 
.A1(n_4768),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4825),
.Y(n_5289)
);

AOI22xp33_ASAP7_75t_L g5290 ( 
.A1(n_4979),
.A2(n_700),
.B1(n_697),
.B2(n_699),
.Y(n_5290)
);

INVxp67_ASAP7_75t_L g5291 ( 
.A(n_4932),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_4836),
.Y(n_5292)
);

INVx2_ASAP7_75t_L g5293 ( 
.A(n_4844),
.Y(n_5293)
);

NAND2x1p5_ASAP7_75t_L g5294 ( 
.A(n_4775),
.B(n_5040),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4861),
.Y(n_5295)
);

BUFx3_ASAP7_75t_L g5296 ( 
.A(n_4914),
.Y(n_5296)
);

AOI22xp33_ASAP7_75t_SL g5297 ( 
.A1(n_4680),
.A2(n_4898),
.B1(n_5046),
.B2(n_4743),
.Y(n_5297)
);

BUFx3_ASAP7_75t_L g5298 ( 
.A(n_4947),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_4916),
.Y(n_5299)
);

OAI22xp5_ASAP7_75t_L g5300 ( 
.A1(n_4683),
.A2(n_701),
.B1(n_699),
.B2(n_700),
.Y(n_5300)
);

INVx1_ASAP7_75t_SL g5301 ( 
.A(n_4869),
.Y(n_5301)
);

OAI22xp33_ASAP7_75t_L g5302 ( 
.A1(n_5060),
.A2(n_4937),
.B1(n_5004),
.B2(n_5000),
.Y(n_5302)
);

AOI22xp33_ASAP7_75t_L g5303 ( 
.A1(n_5034),
.A2(n_704),
.B1(n_699),
.B2(n_702),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4925),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4928),
.Y(n_5305)
);

INVx2_ASAP7_75t_L g5306 ( 
.A(n_4966),
.Y(n_5306)
);

OAI21xp5_ASAP7_75t_SL g5307 ( 
.A1(n_4710),
.A2(n_702),
.B(n_704),
.Y(n_5307)
);

CKINVDCx20_ASAP7_75t_R g5308 ( 
.A(n_4700),
.Y(n_5308)
);

BUFx2_ASAP7_75t_L g5309 ( 
.A(n_4890),
.Y(n_5309)
);

OAI22xp5_ASAP7_75t_L g5310 ( 
.A1(n_4771),
.A2(n_706),
.B1(n_702),
.B2(n_705),
.Y(n_5310)
);

OAI22xp5_ASAP7_75t_L g5311 ( 
.A1(n_4946),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_5311)
);

BUFx3_ASAP7_75t_L g5312 ( 
.A(n_4761),
.Y(n_5312)
);

BUFx10_ASAP7_75t_L g5313 ( 
.A(n_4667),
.Y(n_5313)
);

AOI22xp33_ASAP7_75t_L g5314 ( 
.A1(n_5010),
.A2(n_5017),
.B1(n_5013),
.B2(n_4988),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_4992),
.Y(n_5315)
);

BUFx2_ASAP7_75t_L g5316 ( 
.A(n_4636),
.Y(n_5316)
);

OAI22xp5_ASAP7_75t_L g5317 ( 
.A1(n_5024),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_5317)
);

CKINVDCx6p67_ASAP7_75t_R g5318 ( 
.A(n_4853),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_4994),
.Y(n_5319)
);

BUFx4f_ASAP7_75t_SL g5320 ( 
.A(n_4954),
.Y(n_5320)
);

BUFx6f_ASAP7_75t_L g5321 ( 
.A(n_4632),
.Y(n_5321)
);

BUFx2_ASAP7_75t_SL g5322 ( 
.A(n_4633),
.Y(n_5322)
);

INVxp67_ASAP7_75t_L g5323 ( 
.A(n_4968),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_4637),
.B(n_4760),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5023),
.Y(n_5325)
);

CKINVDCx20_ASAP7_75t_R g5326 ( 
.A(n_4998),
.Y(n_5326)
);

INVx2_ASAP7_75t_SL g5327 ( 
.A(n_5002),
.Y(n_5327)
);

INVx3_ASAP7_75t_L g5328 ( 
.A(n_4976),
.Y(n_5328)
);

NAND2x1p5_ASAP7_75t_L g5329 ( 
.A(n_5030),
.B(n_707),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5026),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5042),
.Y(n_5331)
);

AOI22xp33_ASAP7_75t_L g5332 ( 
.A1(n_4726),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_5332)
);

AOI22xp33_ASAP7_75t_L g5333 ( 
.A1(n_5005),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_5333)
);

BUFx12f_ASAP7_75t_L g5334 ( 
.A(n_5019),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4873),
.Y(n_5335)
);

AOI22xp33_ASAP7_75t_L g5336 ( 
.A1(n_4986),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_4910),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_4912),
.Y(n_5338)
);

INVx6_ASAP7_75t_L g5339 ( 
.A(n_5027),
.Y(n_5339)
);

CKINVDCx5p33_ASAP7_75t_R g5340 ( 
.A(n_4993),
.Y(n_5340)
);

CKINVDCx20_ASAP7_75t_R g5341 ( 
.A(n_4754),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_4654),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4670),
.Y(n_5343)
);

CKINVDCx6p67_ASAP7_75t_R g5344 ( 
.A(n_4955),
.Y(n_5344)
);

INVx2_ASAP7_75t_L g5345 ( 
.A(n_4743),
.Y(n_5345)
);

OAI22xp5_ASAP7_75t_L g5346 ( 
.A1(n_5051),
.A2(n_714),
.B1(n_712),
.B2(n_713),
.Y(n_5346)
);

CKINVDCx20_ASAP7_75t_R g5347 ( 
.A(n_4939),
.Y(n_5347)
);

OAI22xp33_ASAP7_75t_L g5348 ( 
.A1(n_4999),
.A2(n_5025),
.B1(n_4803),
.B2(n_4804),
.Y(n_5348)
);

OAI22xp5_ASAP7_75t_L g5349 ( 
.A1(n_4776),
.A2(n_715),
.B1(n_712),
.B2(n_713),
.Y(n_5349)
);

INVx1_ASAP7_75t_SL g5350 ( 
.A(n_4980),
.Y(n_5350)
);

AOI22xp33_ASAP7_75t_L g5351 ( 
.A1(n_4789),
.A2(n_716),
.B1(n_713),
.B2(n_715),
.Y(n_5351)
);

INVx4_ASAP7_75t_L g5352 ( 
.A(n_4898),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_4676),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5050),
.Y(n_5354)
);

INVx3_ASAP7_75t_L g5355 ( 
.A(n_4675),
.Y(n_5355)
);

CKINVDCx11_ASAP7_75t_R g5356 ( 
.A(n_4985),
.Y(n_5356)
);

BUFx8_ASAP7_75t_L g5357 ( 
.A(n_4692),
.Y(n_5357)
);

BUFx3_ASAP7_75t_L g5358 ( 
.A(n_4990),
.Y(n_5358)
);

AOI22xp33_ASAP7_75t_L g5359 ( 
.A1(n_4682),
.A2(n_717),
.B1(n_715),
.B2(n_716),
.Y(n_5359)
);

HB1xp67_ASAP7_75t_L g5360 ( 
.A(n_4718),
.Y(n_5360)
);

INVx6_ASAP7_75t_L g5361 ( 
.A(n_4772),
.Y(n_5361)
);

CKINVDCx20_ASAP7_75t_R g5362 ( 
.A(n_4862),
.Y(n_5362)
);

INVx6_ASAP7_75t_L g5363 ( 
.A(n_4949),
.Y(n_5363)
);

CKINVDCx5p33_ASAP7_75t_R g5364 ( 
.A(n_4824),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_5050),
.Y(n_5365)
);

INVx6_ASAP7_75t_L g5366 ( 
.A(n_4692),
.Y(n_5366)
);

CKINVDCx20_ASAP7_75t_R g5367 ( 
.A(n_4740),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_4882),
.Y(n_5368)
);

AOI22xp33_ASAP7_75t_L g5369 ( 
.A1(n_4694),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_5369)
);

OAI22xp5_ASAP7_75t_L g5370 ( 
.A1(n_4859),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_5370)
);

INVx6_ASAP7_75t_L g5371 ( 
.A(n_4675),
.Y(n_5371)
);

OAI22xp5_ASAP7_75t_L g5372 ( 
.A1(n_4756),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4882),
.Y(n_5373)
);

INVx2_ASAP7_75t_L g5374 ( 
.A(n_4695),
.Y(n_5374)
);

AOI22xp33_ASAP7_75t_L g5375 ( 
.A1(n_4691),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_5064),
.Y(n_5376)
);

NAND2xp5_ASAP7_75t_L g5377 ( 
.A(n_5169),
.B(n_5009),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_5084),
.Y(n_5378)
);

INVx2_ASAP7_75t_L g5379 ( 
.A(n_5309),
.Y(n_5379)
);

INVx2_ASAP7_75t_L g5380 ( 
.A(n_5203),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5088),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_5206),
.Y(n_5382)
);

AND2x4_ASAP7_75t_L g5383 ( 
.A(n_5195),
.B(n_5239),
.Y(n_5383)
);

INVxp33_ASAP7_75t_L g5384 ( 
.A(n_5130),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5089),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_5080),
.Y(n_5386)
);

NAND2xp5_ASAP7_75t_L g5387 ( 
.A(n_5188),
.B(n_5033),
.Y(n_5387)
);

BUFx2_ASAP7_75t_L g5388 ( 
.A(n_5237),
.Y(n_5388)
);

AND2x2_ASAP7_75t_L g5389 ( 
.A(n_5143),
.B(n_4769),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_5090),
.Y(n_5390)
);

INVx2_ASAP7_75t_L g5391 ( 
.A(n_5087),
.Y(n_5391)
);

CKINVDCx20_ASAP7_75t_R g5392 ( 
.A(n_5119),
.Y(n_5392)
);

INVx2_ASAP7_75t_SL g5393 ( 
.A(n_5081),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_5093),
.Y(n_5394)
);

AND2x2_ASAP7_75t_L g5395 ( 
.A(n_5067),
.B(n_4593),
.Y(n_5395)
);

INVxp67_ASAP7_75t_L g5396 ( 
.A(n_5121),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5096),
.Y(n_5397)
);

OR2x6_ASAP7_75t_L g5398 ( 
.A(n_5065),
.B(n_4662),
.Y(n_5398)
);

BUFx2_ASAP7_75t_L g5399 ( 
.A(n_5238),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_5100),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5102),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5104),
.Y(n_5402)
);

OAI21x1_ASAP7_75t_L g5403 ( 
.A1(n_5328),
.A2(n_4742),
.B(n_4767),
.Y(n_5403)
);

INVx2_ASAP7_75t_SL g5404 ( 
.A(n_5081),
.Y(n_5404)
);

NOR3xp33_ASAP7_75t_SL g5405 ( 
.A(n_5340),
.B(n_4943),
.C(n_4762),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5078),
.Y(n_5406)
);

INVx1_ASAP7_75t_SL g5407 ( 
.A(n_5082),
.Y(n_5407)
);

INVx2_ASAP7_75t_SL g5408 ( 
.A(n_5073),
.Y(n_5408)
);

AOI22xp33_ASAP7_75t_SL g5409 ( 
.A1(n_5357),
.A2(n_4695),
.B1(n_5020),
.B2(n_5021),
.Y(n_5409)
);

AOI21x1_ASAP7_75t_L g5410 ( 
.A1(n_5360),
.A2(n_4900),
.B(n_4935),
.Y(n_5410)
);

INVx3_ASAP7_75t_L g5411 ( 
.A(n_5128),
.Y(n_5411)
);

OAI21x1_ASAP7_75t_L g5412 ( 
.A1(n_5355),
.A2(n_5345),
.B(n_5374),
.Y(n_5412)
);

INVx3_ASAP7_75t_L g5413 ( 
.A(n_5065),
.Y(n_5413)
);

INVx2_ASAP7_75t_SL g5414 ( 
.A(n_5073),
.Y(n_5414)
);

CKINVDCx6p67_ASAP7_75t_R g5415 ( 
.A(n_5103),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5131),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5127),
.Y(n_5417)
);

OAI21x1_ASAP7_75t_L g5418 ( 
.A1(n_5368),
.A2(n_4602),
.B(n_4805),
.Y(n_5418)
);

OAI21xp33_ASAP7_75t_SL g5419 ( 
.A1(n_5134),
.A2(n_4690),
.B(n_5053),
.Y(n_5419)
);

BUFx6f_ASAP7_75t_L g5420 ( 
.A(n_5066),
.Y(n_5420)
);

INVx2_ASAP7_75t_L g5421 ( 
.A(n_5138),
.Y(n_5421)
);

NOR2xp33_ASAP7_75t_L g5422 ( 
.A(n_5197),
.B(n_4995),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5124),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5154),
.Y(n_5424)
);

INVx2_ASAP7_75t_L g5425 ( 
.A(n_5141),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_5145),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_5136),
.Y(n_5427)
);

HB1xp67_ASAP7_75t_L g5428 ( 
.A(n_5224),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_5142),
.Y(n_5429)
);

AND2x2_ASAP7_75t_L g5430 ( 
.A(n_5202),
.B(n_4593),
.Y(n_5430)
);

NOR2x1_ASAP7_75t_SL g5431 ( 
.A(n_5233),
.B(n_4707),
.Y(n_5431)
);

AO21x2_ASAP7_75t_L g5432 ( 
.A1(n_5208),
.A2(n_4807),
.B(n_4958),
.Y(n_5432)
);

HB1xp67_ASAP7_75t_L g5433 ( 
.A(n_5111),
.Y(n_5433)
);

HB1xp67_ASAP7_75t_L g5434 ( 
.A(n_5210),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5106),
.Y(n_5435)
);

OAI21x1_ASAP7_75t_L g5436 ( 
.A1(n_5373),
.A2(n_4621),
.B(n_4974),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5156),
.Y(n_5437)
);

INVx2_ASAP7_75t_SL g5438 ( 
.A(n_5174),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5171),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_5200),
.Y(n_5440)
);

INVx2_ASAP7_75t_L g5441 ( 
.A(n_5158),
.Y(n_5441)
);

INVx2_ASAP7_75t_SL g5442 ( 
.A(n_5147),
.Y(n_5442)
);

INVx2_ASAP7_75t_L g5443 ( 
.A(n_5175),
.Y(n_5443)
);

BUFx6f_ASAP7_75t_L g5444 ( 
.A(n_5152),
.Y(n_5444)
);

OA21x2_ASAP7_75t_L g5445 ( 
.A1(n_5316),
.A2(n_4895),
.B(n_4738),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_L g5446 ( 
.A(n_5178),
.B(n_5063),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_5170),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5201),
.Y(n_5448)
);

INVx2_ASAP7_75t_SL g5449 ( 
.A(n_5135),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5183),
.Y(n_5450)
);

AOI22xp5_ASAP7_75t_L g5451 ( 
.A1(n_5101),
.A2(n_5076),
.B1(n_5072),
.B2(n_5172),
.Y(n_5451)
);

INVx2_ASAP7_75t_L g5452 ( 
.A(n_5204),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5116),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5234),
.Y(n_5454)
);

AND2x2_ASAP7_75t_L g5455 ( 
.A(n_5241),
.B(n_4718),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_5263),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_5267),
.Y(n_5457)
);

HB1xp67_ASAP7_75t_L g5458 ( 
.A(n_5298),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5279),
.Y(n_5459)
);

OAI21x1_ASAP7_75t_L g5460 ( 
.A1(n_5161),
.A2(n_4655),
.B(n_5018),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5281),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5289),
.Y(n_5462)
);

INVx2_ASAP7_75t_L g5463 ( 
.A(n_5213),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5295),
.Y(n_5464)
);

AOI22xp33_ASAP7_75t_L g5465 ( 
.A1(n_5275),
.A2(n_4752),
.B1(n_4933),
.B2(n_4929),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5299),
.Y(n_5466)
);

OAI21x1_ASAP7_75t_L g5467 ( 
.A1(n_5173),
.A2(n_4665),
.B(n_4790),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5304),
.Y(n_5468)
);

AND2x4_ASAP7_75t_L g5469 ( 
.A(n_5324),
.B(n_4753),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_5214),
.Y(n_5470)
);

AO31x2_ASAP7_75t_L g5471 ( 
.A1(n_5199),
.A2(n_4806),
.A3(n_4835),
.B(n_4813),
.Y(n_5471)
);

AND2x2_ASAP7_75t_L g5472 ( 
.A(n_5327),
.B(n_4649),
.Y(n_5472)
);

HB1xp67_ASAP7_75t_L g5473 ( 
.A(n_5250),
.Y(n_5473)
);

OR2x6_ASAP7_75t_L g5474 ( 
.A(n_5189),
.B(n_4963),
.Y(n_5474)
);

NOR2xp67_ASAP7_75t_L g5475 ( 
.A(n_5139),
.B(n_4964),
.Y(n_5475)
);

BUFx2_ASAP7_75t_L g5476 ( 
.A(n_5238),
.Y(n_5476)
);

AND2x2_ASAP7_75t_L g5477 ( 
.A(n_5226),
.B(n_4649),
.Y(n_5477)
);

AND2x4_ASAP7_75t_L g5478 ( 
.A(n_5194),
.B(n_5182),
.Y(n_5478)
);

HB1xp67_ASAP7_75t_L g5479 ( 
.A(n_5274),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5305),
.Y(n_5480)
);

INVxp67_ASAP7_75t_L g5481 ( 
.A(n_5083),
.Y(n_5481)
);

AND2x2_ASAP7_75t_SL g5482 ( 
.A(n_5192),
.B(n_4885),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_5292),
.Y(n_5483)
);

AND2x4_ASAP7_75t_L g5484 ( 
.A(n_5315),
.B(n_4781),
.Y(n_5484)
);

INVx2_ASAP7_75t_L g5485 ( 
.A(n_5293),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5306),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_5319),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_5352),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_5325),
.Y(n_5489)
);

INVx2_ASAP7_75t_SL g5490 ( 
.A(n_5135),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5330),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5331),
.Y(n_5492)
);

OAI21x1_ASAP7_75t_L g5493 ( 
.A1(n_5193),
.A2(n_4903),
.B(n_4889),
.Y(n_5493)
);

OAI21x1_ASAP7_75t_L g5494 ( 
.A1(n_5187),
.A2(n_4944),
.B(n_4934),
.Y(n_5494)
);

OAI22xp33_ASAP7_75t_L g5495 ( 
.A1(n_5259),
.A2(n_5035),
.B1(n_5043),
.B2(n_4863),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5335),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5337),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5338),
.Y(n_5498)
);

NOR2xp33_ASAP7_75t_L g5499 ( 
.A(n_5191),
.B(n_5006),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_5071),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_5271),
.Y(n_5501)
);

INVx2_ASAP7_75t_L g5502 ( 
.A(n_5266),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5140),
.Y(n_5503)
);

INVx3_ASAP7_75t_L g5504 ( 
.A(n_5165),
.Y(n_5504)
);

INVx2_ASAP7_75t_L g5505 ( 
.A(n_5283),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_5092),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5342),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5343),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5353),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5366),
.Y(n_5510)
);

OAI21x1_ASAP7_75t_L g5511 ( 
.A1(n_5329),
.A2(n_4685),
.B(n_4590),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5366),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5356),
.Y(n_5513)
);

INVx3_ASAP7_75t_L g5514 ( 
.A(n_5165),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5354),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5365),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5069),
.Y(n_5517)
);

A2O1A1Ixp33_ASAP7_75t_L g5518 ( 
.A1(n_5307),
.A2(n_4956),
.B(n_4699),
.C(n_4786),
.Y(n_5518)
);

BUFx2_ASAP7_75t_L g5519 ( 
.A(n_5258),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5273),
.Y(n_5520)
);

OR2x6_ASAP7_75t_L g5521 ( 
.A(n_5189),
.B(n_5029),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_5229),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5276),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5235),
.Y(n_5524)
);

AOI21xp5_ASAP7_75t_L g5525 ( 
.A1(n_5150),
.A2(n_5039),
.B(n_4905),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5301),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_5323),
.Y(n_5527)
);

OAI21xp5_ASAP7_75t_L g5528 ( 
.A1(n_5215),
.A2(n_4924),
.B(n_4951),
.Y(n_5528)
);

AND2x2_ASAP7_75t_L g5529 ( 
.A(n_5265),
.B(n_4656),
.Y(n_5529)
);

INVx4_ASAP7_75t_L g5530 ( 
.A(n_5228),
.Y(n_5530)
);

AO31x2_ASAP7_75t_L g5531 ( 
.A1(n_5244),
.A2(n_4830),
.A3(n_4671),
.B(n_4668),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5312),
.B(n_4656),
.Y(n_5532)
);

INVx2_ASAP7_75t_L g5533 ( 
.A(n_5264),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5291),
.Y(n_5534)
);

NAND2xp5_ASAP7_75t_L g5535 ( 
.A(n_5350),
.B(n_4837),
.Y(n_5535)
);

AOI22xp33_ASAP7_75t_L g5536 ( 
.A1(n_5361),
.A2(n_4759),
.B1(n_4815),
.B2(n_4874),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5186),
.Y(n_5537)
);

NAND2xp5_ASAP7_75t_L g5538 ( 
.A(n_5162),
.B(n_4837),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_L g5539 ( 
.A(n_5242),
.B(n_4722),
.Y(n_5539)
);

OR2x2_ASAP7_75t_L g5540 ( 
.A(n_5358),
.B(n_4872),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5296),
.Y(n_5541)
);

HB1xp67_ASAP7_75t_L g5542 ( 
.A(n_5163),
.Y(n_5542)
);

BUFx3_ASAP7_75t_L g5543 ( 
.A(n_5392),
.Y(n_5543)
);

INVx2_ASAP7_75t_L g5544 ( 
.A(n_5388),
.Y(n_5544)
);

INVx2_ASAP7_75t_SL g5545 ( 
.A(n_5411),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5376),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5378),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_5381),
.Y(n_5548)
);

OR2x2_ASAP7_75t_L g5549 ( 
.A(n_5377),
.B(n_5108),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5385),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5390),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5400),
.Y(n_5552)
);

AO21x2_ASAP7_75t_L g5553 ( 
.A1(n_5403),
.A2(n_5282),
.B(n_5168),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5401),
.Y(n_5554)
);

INVx2_ASAP7_75t_L g5555 ( 
.A(n_5388),
.Y(n_5555)
);

OR2x2_ASAP7_75t_L g5556 ( 
.A(n_5453),
.B(n_5153),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5402),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_5415),
.Y(n_5558)
);

INVx2_ASAP7_75t_L g5559 ( 
.A(n_5383),
.Y(n_5559)
);

BUFx6f_ASAP7_75t_L g5560 ( 
.A(n_5420),
.Y(n_5560)
);

HB1xp67_ASAP7_75t_L g5561 ( 
.A(n_5458),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_5383),
.Y(n_5562)
);

HB1xp67_ASAP7_75t_L g5563 ( 
.A(n_5428),
.Y(n_5563)
);

NAND2xp5_ASAP7_75t_L g5564 ( 
.A(n_5517),
.B(n_5252),
.Y(n_5564)
);

AND2x4_ASAP7_75t_L g5565 ( 
.A(n_5510),
.B(n_5321),
.Y(n_5565)
);

HB1xp67_ASAP7_75t_L g5566 ( 
.A(n_5379),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_5470),
.Y(n_5567)
);

NOR2xp33_ASAP7_75t_L g5568 ( 
.A(n_5384),
.B(n_5118),
.Y(n_5568)
);

NAND2x1p5_ASAP7_75t_L g5569 ( 
.A(n_5530),
.B(n_5139),
.Y(n_5569)
);

HB1xp67_ASAP7_75t_L g5570 ( 
.A(n_5479),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5423),
.Y(n_5571)
);

AND2x2_ASAP7_75t_L g5572 ( 
.A(n_5478),
.B(n_5344),
.Y(n_5572)
);

INVx2_ASAP7_75t_L g5573 ( 
.A(n_5519),
.Y(n_5573)
);

HB1xp67_ASAP7_75t_L g5574 ( 
.A(n_5399),
.Y(n_5574)
);

OR2x6_ASAP7_75t_L g5575 ( 
.A(n_5399),
.B(n_5077),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_5519),
.Y(n_5576)
);

INVx3_ASAP7_75t_L g5577 ( 
.A(n_5482),
.Y(n_5577)
);

AND2x2_ASAP7_75t_L g5578 ( 
.A(n_5478),
.B(n_5318),
.Y(n_5578)
);

INVx2_ASAP7_75t_L g5579 ( 
.A(n_5441),
.Y(n_5579)
);

AO21x2_ASAP7_75t_L g5580 ( 
.A1(n_5410),
.A2(n_5277),
.B(n_5269),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5427),
.Y(n_5581)
);

AND2x4_ASAP7_75t_L g5582 ( 
.A(n_5512),
.B(n_5321),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5416),
.Y(n_5583)
);

AND2x2_ASAP7_75t_L g5584 ( 
.A(n_5433),
.B(n_5216),
.Y(n_5584)
);

AO21x2_ASAP7_75t_L g5585 ( 
.A1(n_5410),
.A2(n_5262),
.B(n_5236),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_5426),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5380),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5382),
.Y(n_5588)
);

HB1xp67_ASAP7_75t_L g5589 ( 
.A(n_5476),
.Y(n_5589)
);

INVx3_ASAP7_75t_L g5590 ( 
.A(n_5420),
.Y(n_5590)
);

AO21x2_ASAP7_75t_L g5591 ( 
.A1(n_5535),
.A2(n_5098),
.B(n_5243),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5507),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5508),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_5509),
.Y(n_5594)
);

INVxp67_ASAP7_75t_SL g5595 ( 
.A(n_5434),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5443),
.Y(n_5596)
);

BUFx3_ASAP7_75t_L g5597 ( 
.A(n_5408),
.Y(n_5597)
);

OR2x6_ASAP7_75t_L g5598 ( 
.A(n_5476),
.B(n_5196),
.Y(n_5598)
);

HB1xp67_ASAP7_75t_L g5599 ( 
.A(n_5473),
.Y(n_5599)
);

OAI21x1_ASAP7_75t_L g5600 ( 
.A1(n_5412),
.A2(n_5294),
.B(n_4984),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5440),
.Y(n_5601)
);

INVx3_ASAP7_75t_L g5602 ( 
.A(n_5488),
.Y(n_5602)
);

OA21x2_ASAP7_75t_L g5603 ( 
.A1(n_5537),
.A2(n_5245),
.B(n_5070),
.Y(n_5603)
);

AND2x2_ASAP7_75t_L g5604 ( 
.A(n_5520),
.B(n_5220),
.Y(n_5604)
);

INVx2_ASAP7_75t_SL g5605 ( 
.A(n_5444),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5435),
.Y(n_5606)
);

INVxp67_ASAP7_75t_L g5607 ( 
.A(n_5407),
.Y(n_5607)
);

AOI22xp33_ASAP7_75t_L g5608 ( 
.A1(n_5451),
.A2(n_5361),
.B1(n_5320),
.B2(n_5363),
.Y(n_5608)
);

AND2x2_ASAP7_75t_L g5609 ( 
.A(n_5406),
.B(n_5285),
.Y(n_5609)
);

AND2x2_ASAP7_75t_L g5610 ( 
.A(n_5424),
.B(n_5280),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5447),
.Y(n_5611)
);

AO21x2_ASAP7_75t_L g5612 ( 
.A1(n_5538),
.A2(n_5257),
.B(n_5110),
.Y(n_5612)
);

AND2x2_ASAP7_75t_L g5613 ( 
.A(n_5455),
.B(n_5371),
.Y(n_5613)
);

AO21x2_ASAP7_75t_L g5614 ( 
.A1(n_5525),
.A2(n_4681),
.B(n_5251),
.Y(n_5614)
);

BUFx2_ASAP7_75t_L g5615 ( 
.A(n_5542),
.Y(n_5615)
);

INVx3_ASAP7_75t_L g5616 ( 
.A(n_5413),
.Y(n_5616)
);

OR2x2_ASAP7_75t_L g5617 ( 
.A(n_5500),
.B(n_5153),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_5437),
.Y(n_5618)
);

AND2x4_ASAP7_75t_L g5619 ( 
.A(n_5395),
.B(n_5163),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5448),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5529),
.B(n_5297),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5421),
.Y(n_5622)
);

OA21x2_ASAP7_75t_L g5623 ( 
.A1(n_5436),
.A2(n_5074),
.B(n_4773),
.Y(n_5623)
);

AO21x2_ASAP7_75t_L g5624 ( 
.A1(n_5431),
.A2(n_5231),
.B(n_5105),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_5425),
.Y(n_5625)
);

BUFx2_ASAP7_75t_L g5626 ( 
.A(n_5396),
.Y(n_5626)
);

AND2x4_ASAP7_75t_L g5627 ( 
.A(n_5430),
.B(n_5068),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5429),
.Y(n_5628)
);

INVx3_ASAP7_75t_L g5629 ( 
.A(n_5444),
.Y(n_5629)
);

INVx1_ASAP7_75t_SL g5630 ( 
.A(n_5414),
.Y(n_5630)
);

BUFx2_ASAP7_75t_L g5631 ( 
.A(n_5442),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_5386),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_5391),
.Y(n_5633)
);

BUFx2_ASAP7_75t_L g5634 ( 
.A(n_5504),
.Y(n_5634)
);

AND2x2_ASAP7_75t_L g5635 ( 
.A(n_5526),
.B(n_5371),
.Y(n_5635)
);

BUFx3_ASAP7_75t_L g5636 ( 
.A(n_5438),
.Y(n_5636)
);

AND2x4_ASAP7_75t_L g5637 ( 
.A(n_5469),
.B(n_5152),
.Y(n_5637)
);

AO21x2_ASAP7_75t_L g5638 ( 
.A1(n_5515),
.A2(n_5516),
.B(n_5460),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5439),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5454),
.Y(n_5640)
);

INVx1_ASAP7_75t_SL g5641 ( 
.A(n_5393),
.Y(n_5641)
);

CKINVDCx5p33_ASAP7_75t_R g5642 ( 
.A(n_5404),
.Y(n_5642)
);

NAND3xp33_ASAP7_75t_L g5643 ( 
.A(n_5419),
.B(n_5207),
.C(n_5364),
.Y(n_5643)
);

NAND2xp5_ASAP7_75t_L g5644 ( 
.A(n_5523),
.B(n_5314),
.Y(n_5644)
);

NOR2xp33_ASAP7_75t_L g5645 ( 
.A(n_5505),
.B(n_5132),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_L g5646 ( 
.A(n_5503),
.B(n_5506),
.Y(n_5646)
);

AND2x2_ASAP7_75t_L g5647 ( 
.A(n_5389),
.B(n_5112),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5456),
.Y(n_5648)
);

INVx1_ASAP7_75t_L g5649 ( 
.A(n_5457),
.Y(n_5649)
);

HB1xp67_ASAP7_75t_L g5650 ( 
.A(n_5501),
.Y(n_5650)
);

INVx3_ASAP7_75t_L g5651 ( 
.A(n_5514),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5394),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_5459),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_5397),
.Y(n_5654)
);

HB1xp67_ASAP7_75t_L g5655 ( 
.A(n_5502),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5461),
.Y(n_5656)
);

OR2x2_ASAP7_75t_L g5657 ( 
.A(n_5417),
.B(n_5322),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5534),
.B(n_5254),
.Y(n_5658)
);

INVxp67_ASAP7_75t_SL g5659 ( 
.A(n_5481),
.Y(n_5659)
);

AOI22xp33_ASAP7_75t_L g5660 ( 
.A1(n_5409),
.A2(n_5363),
.B1(n_5255),
.B2(n_5339),
.Y(n_5660)
);

HB1xp67_ASAP7_75t_L g5661 ( 
.A(n_5452),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5462),
.Y(n_5662)
);

BUFx2_ASAP7_75t_L g5663 ( 
.A(n_5513),
.Y(n_5663)
);

INVx3_ASAP7_75t_L g5664 ( 
.A(n_5449),
.Y(n_5664)
);

AOI21x1_ASAP7_75t_L g5665 ( 
.A1(n_5475),
.A2(n_5107),
.B(n_5310),
.Y(n_5665)
);

BUFx2_ASAP7_75t_L g5666 ( 
.A(n_5490),
.Y(n_5666)
);

INVx2_ASAP7_75t_L g5667 ( 
.A(n_5483),
.Y(n_5667)
);

INVx2_ASAP7_75t_L g5668 ( 
.A(n_5485),
.Y(n_5668)
);

NOR3xp33_ASAP7_75t_L g5669 ( 
.A(n_5495),
.B(n_5164),
.C(n_5091),
.Y(n_5669)
);

AND2x4_ASAP7_75t_L g5670 ( 
.A(n_5469),
.B(n_5472),
.Y(n_5670)
);

OR2x6_ASAP7_75t_L g5671 ( 
.A(n_5398),
.B(n_5196),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5464),
.Y(n_5672)
);

HB1xp67_ASAP7_75t_L g5673 ( 
.A(n_5463),
.Y(n_5673)
);

CKINVDCx5p33_ASAP7_75t_R g5674 ( 
.A(n_5422),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5466),
.Y(n_5675)
);

AND2x2_ASAP7_75t_L g5676 ( 
.A(n_5559),
.B(n_5527),
.Y(n_5676)
);

HB1xp67_ASAP7_75t_L g5677 ( 
.A(n_5561),
.Y(n_5677)
);

AND2x2_ASAP7_75t_L g5678 ( 
.A(n_5562),
.B(n_5541),
.Y(n_5678)
);

NAND2xp5_ASAP7_75t_L g5679 ( 
.A(n_5644),
.B(n_5477),
.Y(n_5679)
);

AND2x2_ASAP7_75t_L g5680 ( 
.A(n_5670),
.B(n_5532),
.Y(n_5680)
);

INVx1_ASAP7_75t_SL g5681 ( 
.A(n_5642),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5615),
.Y(n_5682)
);

HB1xp67_ASAP7_75t_L g5683 ( 
.A(n_5650),
.Y(n_5683)
);

AOI22xp33_ASAP7_75t_L g5684 ( 
.A1(n_5669),
.A2(n_5521),
.B1(n_5474),
.B2(n_5398),
.Y(n_5684)
);

OR2x2_ASAP7_75t_L g5685 ( 
.A(n_5661),
.B(n_5450),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5615),
.Y(n_5686)
);

NOR2x1_ASAP7_75t_SL g5687 ( 
.A(n_5575),
.B(n_5085),
.Y(n_5687)
);

AND2x2_ASAP7_75t_L g5688 ( 
.A(n_5670),
.B(n_5627),
.Y(n_5688)
);

AND2x2_ASAP7_75t_L g5689 ( 
.A(n_5627),
.B(n_5574),
.Y(n_5689)
);

NAND2xp5_ASAP7_75t_L g5690 ( 
.A(n_5564),
.B(n_5539),
.Y(n_5690)
);

INVx2_ASAP7_75t_L g5691 ( 
.A(n_5655),
.Y(n_5691)
);

AND2x4_ASAP7_75t_L g5692 ( 
.A(n_5577),
.B(n_5492),
.Y(n_5692)
);

AND2x4_ASAP7_75t_L g5693 ( 
.A(n_5577),
.B(n_5522),
.Y(n_5693)
);

AND2x2_ASAP7_75t_L g5694 ( 
.A(n_5589),
.B(n_5524),
.Y(n_5694)
);

OAI221xp5_ASAP7_75t_L g5695 ( 
.A1(n_5660),
.A2(n_5518),
.B1(n_5528),
.B2(n_5405),
.C(n_5465),
.Y(n_5695)
);

INVx2_ASAP7_75t_SL g5696 ( 
.A(n_5560),
.Y(n_5696)
);

INVx2_ASAP7_75t_L g5697 ( 
.A(n_5673),
.Y(n_5697)
);

NOR2xp33_ASAP7_75t_L g5698 ( 
.A(n_5560),
.B(n_5122),
.Y(n_5698)
);

OA21x2_ASAP7_75t_L g5699 ( 
.A1(n_5621),
.A2(n_5494),
.B(n_5446),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_L g5700 ( 
.A(n_5570),
.B(n_5468),
.Y(n_5700)
);

INVx8_ASAP7_75t_L g5701 ( 
.A(n_5558),
.Y(n_5701)
);

BUFx3_ASAP7_75t_L g5702 ( 
.A(n_5543),
.Y(n_5702)
);

AND2x2_ASAP7_75t_L g5703 ( 
.A(n_5647),
.B(n_5533),
.Y(n_5703)
);

INVx2_ASAP7_75t_L g5704 ( 
.A(n_5602),
.Y(n_5704)
);

INVx2_ASAP7_75t_L g5705 ( 
.A(n_5602),
.Y(n_5705)
);

AND2x2_ASAP7_75t_L g5706 ( 
.A(n_5613),
.B(n_5634),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_SL g5707 ( 
.A(n_5643),
.B(n_5122),
.Y(n_5707)
);

AND2x2_ASAP7_75t_L g5708 ( 
.A(n_5634),
.B(n_5387),
.Y(n_5708)
);

AOI22xp5_ASAP7_75t_L g5709 ( 
.A1(n_5612),
.A2(n_5591),
.B1(n_5608),
.B2(n_5580),
.Y(n_5709)
);

NAND2xp5_ASAP7_75t_L g5710 ( 
.A(n_5563),
.B(n_5480),
.Y(n_5710)
);

NAND2xp5_ASAP7_75t_L g5711 ( 
.A(n_5646),
.B(n_5487),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5587),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5588),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5619),
.B(n_5486),
.Y(n_5714)
);

OR2x2_ASAP7_75t_L g5715 ( 
.A(n_5544),
.B(n_5489),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_5567),
.Y(n_5716)
);

AND2x2_ASAP7_75t_L g5717 ( 
.A(n_5619),
.B(n_5491),
.Y(n_5717)
);

AND2x2_ASAP7_75t_L g5718 ( 
.A(n_5626),
.B(n_5496),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_5632),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5586),
.Y(n_5720)
);

HB1xp67_ASAP7_75t_L g5721 ( 
.A(n_5599),
.Y(n_5721)
);

INVx2_ASAP7_75t_L g5722 ( 
.A(n_5633),
.Y(n_5722)
);

OAI31xp33_ASAP7_75t_SL g5723 ( 
.A1(n_5578),
.A2(n_5177),
.A3(n_5499),
.B(n_5094),
.Y(n_5723)
);

NAND2x1p5_ASAP7_75t_L g5724 ( 
.A(n_5560),
.B(n_5167),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5546),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5547),
.Y(n_5726)
);

INVx1_ASAP7_75t_L g5727 ( 
.A(n_5579),
.Y(n_5727)
);

AO21x2_ASAP7_75t_L g5728 ( 
.A1(n_5553),
.A2(n_5432),
.B(n_5467),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_L g5729 ( 
.A(n_5566),
.B(n_5497),
.Y(n_5729)
);

AND2x2_ASAP7_75t_L g5730 ( 
.A(n_5626),
.B(n_5498),
.Y(n_5730)
);

AND2x2_ASAP7_75t_L g5731 ( 
.A(n_5635),
.B(n_5540),
.Y(n_5731)
);

AND2x2_ASAP7_75t_L g5732 ( 
.A(n_5573),
.B(n_5484),
.Y(n_5732)
);

HB1xp67_ASAP7_75t_L g5733 ( 
.A(n_5631),
.Y(n_5733)
);

AOI21xp5_ASAP7_75t_L g5734 ( 
.A1(n_5671),
.A2(n_5198),
.B(n_5474),
.Y(n_5734)
);

HB1xp67_ASAP7_75t_L g5735 ( 
.A(n_5631),
.Y(n_5735)
);

AND2x4_ASAP7_75t_SL g5736 ( 
.A(n_5575),
.B(n_5123),
.Y(n_5736)
);

BUFx6f_ASAP7_75t_L g5737 ( 
.A(n_5569),
.Y(n_5737)
);

INVx2_ASAP7_75t_L g5738 ( 
.A(n_5652),
.Y(n_5738)
);

HB1xp67_ASAP7_75t_L g5739 ( 
.A(n_5555),
.Y(n_5739)
);

AND2x2_ASAP7_75t_L g5740 ( 
.A(n_5576),
.B(n_5484),
.Y(n_5740)
);

INVx2_ASAP7_75t_SL g5741 ( 
.A(n_5597),
.Y(n_5741)
);

INVx1_ASAP7_75t_L g5742 ( 
.A(n_5596),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5667),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5668),
.Y(n_5744)
);

AND2x2_ASAP7_75t_L g5745 ( 
.A(n_5666),
.B(n_5445),
.Y(n_5745)
);

AND2x2_ASAP7_75t_L g5746 ( 
.A(n_5666),
.B(n_5445),
.Y(n_5746)
);

AOI221x1_ASAP7_75t_L g5747 ( 
.A1(n_5590),
.A2(n_5270),
.B1(n_5248),
.B2(n_5146),
.C(n_4893),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5622),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5654),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_5625),
.Y(n_5750)
);

BUFx3_ASAP7_75t_L g5751 ( 
.A(n_5636),
.Y(n_5751)
);

NAND2xp5_ASAP7_75t_L g5752 ( 
.A(n_5595),
.B(n_5418),
.Y(n_5752)
);

OR2x2_ASAP7_75t_L g5753 ( 
.A(n_5628),
.B(n_5471),
.Y(n_5753)
);

NAND2xp5_ASAP7_75t_L g5754 ( 
.A(n_5639),
.B(n_5493),
.Y(n_5754)
);

BUFx2_ASAP7_75t_L g5755 ( 
.A(n_5598),
.Y(n_5755)
);

HB1xp67_ASAP7_75t_L g5756 ( 
.A(n_5641),
.Y(n_5756)
);

AOI22xp33_ASAP7_75t_L g5757 ( 
.A1(n_5614),
.A2(n_5521),
.B1(n_5339),
.B2(n_5362),
.Y(n_5757)
);

AND2x2_ASAP7_75t_L g5758 ( 
.A(n_5637),
.B(n_5256),
.Y(n_5758)
);

OR2x2_ASAP7_75t_L g5759 ( 
.A(n_5549),
.B(n_5471),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5548),
.Y(n_5760)
);

NAND2xp5_ASAP7_75t_L g5761 ( 
.A(n_5592),
.B(n_5531),
.Y(n_5761)
);

NOR2xp33_ASAP7_75t_L g5762 ( 
.A(n_5568),
.B(n_5217),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_5657),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_5550),
.Y(n_5764)
);

HB1xp67_ASAP7_75t_L g5765 ( 
.A(n_5607),
.Y(n_5765)
);

HB1xp67_ASAP7_75t_L g5766 ( 
.A(n_5659),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5551),
.Y(n_5767)
);

AOI22xp33_ASAP7_75t_L g5768 ( 
.A1(n_5603),
.A2(n_5284),
.B1(n_5223),
.B2(n_5367),
.Y(n_5768)
);

AND2x2_ASAP7_75t_L g5769 ( 
.A(n_5637),
.B(n_5190),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5552),
.Y(n_5770)
);

HB1xp67_ASAP7_75t_L g5771 ( 
.A(n_5630),
.Y(n_5771)
);

NAND2xp5_ASAP7_75t_L g5772 ( 
.A(n_5593),
.B(n_5531),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5554),
.Y(n_5773)
);

INVx3_ASAP7_75t_L g5774 ( 
.A(n_5598),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5557),
.Y(n_5775)
);

AND2x2_ASAP7_75t_L g5776 ( 
.A(n_5663),
.B(n_5651),
.Y(n_5776)
);

HB1xp67_ASAP7_75t_L g5777 ( 
.A(n_5663),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5571),
.Y(n_5778)
);

INVxp67_ASAP7_75t_L g5779 ( 
.A(n_5584),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5581),
.Y(n_5780)
);

INVx3_ASAP7_75t_L g5781 ( 
.A(n_5671),
.Y(n_5781)
);

AOI22xp33_ASAP7_75t_L g5782 ( 
.A1(n_5603),
.A2(n_5313),
.B1(n_5247),
.B2(n_5347),
.Y(n_5782)
);

HB1xp67_ASAP7_75t_L g5783 ( 
.A(n_5545),
.Y(n_5783)
);

HB1xp67_ASAP7_75t_L g5784 ( 
.A(n_5583),
.Y(n_5784)
);

AND2x2_ASAP7_75t_L g5785 ( 
.A(n_5572),
.B(n_5205),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5640),
.Y(n_5786)
);

AND2x2_ASAP7_75t_L g5787 ( 
.A(n_5664),
.B(n_5205),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_5648),
.Y(n_5788)
);

OR2x2_ASAP7_75t_L g5789 ( 
.A(n_5594),
.B(n_5471),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5649),
.Y(n_5790)
);

INVx2_ASAP7_75t_L g5791 ( 
.A(n_5653),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5656),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5662),
.Y(n_5793)
);

AND2x4_ASAP7_75t_L g5794 ( 
.A(n_5565),
.B(n_5287),
.Y(n_5794)
);

BUFx2_ASAP7_75t_L g5795 ( 
.A(n_5751),
.Y(n_5795)
);

AND2x2_ASAP7_75t_L g5796 ( 
.A(n_5755),
.B(n_5604),
.Y(n_5796)
);

BUFx3_ASAP7_75t_L g5797 ( 
.A(n_5701),
.Y(n_5797)
);

OR2x2_ASAP7_75t_L g5798 ( 
.A(n_5683),
.B(n_5601),
.Y(n_5798)
);

INVx2_ASAP7_75t_SL g5799 ( 
.A(n_5736),
.Y(n_5799)
);

HB1xp67_ASAP7_75t_L g5800 ( 
.A(n_5777),
.Y(n_5800)
);

OR2x2_ASAP7_75t_L g5801 ( 
.A(n_5690),
.B(n_5606),
.Y(n_5801)
);

OR2x2_ASAP7_75t_L g5802 ( 
.A(n_5766),
.B(n_5611),
.Y(n_5802)
);

OR2x6_ASAP7_75t_L g5803 ( 
.A(n_5701),
.B(n_5228),
.Y(n_5803)
);

HB1xp67_ASAP7_75t_L g5804 ( 
.A(n_5677),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5774),
.B(n_5616),
.Y(n_5805)
);

INVx2_ASAP7_75t_L g5806 ( 
.A(n_5691),
.Y(n_5806)
);

AND2x2_ASAP7_75t_L g5807 ( 
.A(n_5774),
.B(n_5616),
.Y(n_5807)
);

INVx4_ASAP7_75t_L g5808 ( 
.A(n_5737),
.Y(n_5808)
);

AND2x2_ASAP7_75t_L g5809 ( 
.A(n_5706),
.B(n_5658),
.Y(n_5809)
);

AO221x2_ASAP7_75t_L g5810 ( 
.A1(n_5687),
.A2(n_5126),
.B1(n_5137),
.B2(n_5179),
.C(n_5181),
.Y(n_5810)
);

AO21x2_ASAP7_75t_L g5811 ( 
.A1(n_5709),
.A2(n_5624),
.B(n_5638),
.Y(n_5811)
);

BUFx2_ASAP7_75t_L g5812 ( 
.A(n_5733),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5784),
.Y(n_5813)
);

BUFx2_ASAP7_75t_L g5814 ( 
.A(n_5735),
.Y(n_5814)
);

AND2x4_ASAP7_75t_L g5815 ( 
.A(n_5687),
.B(n_5565),
.Y(n_5815)
);

OR2x2_ASAP7_75t_L g5816 ( 
.A(n_5697),
.B(n_5618),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5685),
.Y(n_5817)
);

AND2x2_ASAP7_75t_L g5818 ( 
.A(n_5680),
.B(n_5605),
.Y(n_5818)
);

AND2x2_ASAP7_75t_L g5819 ( 
.A(n_5689),
.B(n_5781),
.Y(n_5819)
);

NOR2x1_ASAP7_75t_L g5820 ( 
.A(n_5737),
.B(n_5585),
.Y(n_5820)
);

AND2x2_ASAP7_75t_L g5821 ( 
.A(n_5781),
.B(n_5609),
.Y(n_5821)
);

OR2x2_ASAP7_75t_L g5822 ( 
.A(n_5721),
.B(n_5620),
.Y(n_5822)
);

AND2x2_ASAP7_75t_L g5823 ( 
.A(n_5688),
.B(n_5610),
.Y(n_5823)
);

INVx2_ASAP7_75t_SL g5824 ( 
.A(n_5724),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5776),
.B(n_5629),
.Y(n_5825)
);

AND2x2_ASAP7_75t_L g5826 ( 
.A(n_5756),
.B(n_5629),
.Y(n_5826)
);

NAND2xp5_ASAP7_75t_SL g5827 ( 
.A(n_5723),
.B(n_5737),
.Y(n_5827)
);

AND2x2_ASAP7_75t_L g5828 ( 
.A(n_5771),
.B(n_5714),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5760),
.Y(n_5829)
);

AND2x2_ASAP7_75t_L g5830 ( 
.A(n_5717),
.B(n_5582),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_5760),
.Y(n_5831)
);

OR2x2_ASAP7_75t_L g5832 ( 
.A(n_5679),
.B(n_5682),
.Y(n_5832)
);

BUFx2_ASAP7_75t_L g5833 ( 
.A(n_5783),
.Y(n_5833)
);

BUFx2_ASAP7_75t_L g5834 ( 
.A(n_5741),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5767),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5767),
.Y(n_5836)
);

AND2x2_ASAP7_75t_L g5837 ( 
.A(n_5708),
.B(n_5582),
.Y(n_5837)
);

INVx2_ASAP7_75t_L g5838 ( 
.A(n_5727),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5770),
.Y(n_5839)
);

AND2x4_ASAP7_75t_L g5840 ( 
.A(n_5692),
.B(n_5600),
.Y(n_5840)
);

INVx3_ASAP7_75t_L g5841 ( 
.A(n_5702),
.Y(n_5841)
);

AND2x4_ASAP7_75t_L g5842 ( 
.A(n_5692),
.B(n_5617),
.Y(n_5842)
);

NAND2xp5_ASAP7_75t_L g5843 ( 
.A(n_5718),
.B(n_5672),
.Y(n_5843)
);

INVx5_ASAP7_75t_L g5844 ( 
.A(n_5794),
.Y(n_5844)
);

BUFx2_ASAP7_75t_L g5845 ( 
.A(n_5794),
.Y(n_5845)
);

NAND2xp5_ASAP7_75t_L g5846 ( 
.A(n_5730),
.B(n_5675),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5770),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5792),
.Y(n_5848)
);

NAND2xp5_ASAP7_75t_L g5849 ( 
.A(n_5712),
.B(n_5623),
.Y(n_5849)
);

BUFx3_ASAP7_75t_L g5850 ( 
.A(n_5698),
.Y(n_5850)
);

OR2x2_ASAP7_75t_L g5851 ( 
.A(n_5686),
.B(n_5556),
.Y(n_5851)
);

AND2x2_ASAP7_75t_L g5852 ( 
.A(n_5731),
.B(n_5645),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5792),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5793),
.Y(n_5854)
);

AND2x2_ASAP7_75t_L g5855 ( 
.A(n_5693),
.B(n_5623),
.Y(n_5855)
);

INVx2_ASAP7_75t_SL g5856 ( 
.A(n_5758),
.Y(n_5856)
);

INVx2_ASAP7_75t_L g5857 ( 
.A(n_5727),
.Y(n_5857)
);

INVx3_ASAP7_75t_L g5858 ( 
.A(n_5681),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5793),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5748),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5693),
.B(n_5674),
.Y(n_5861)
);

AND2x4_ASAP7_75t_L g5862 ( 
.A(n_5779),
.B(n_5240),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5742),
.Y(n_5863)
);

AND2x2_ASAP7_75t_L g5864 ( 
.A(n_5765),
.B(n_5665),
.Y(n_5864)
);

NOR2xp33_ASAP7_75t_SL g5865 ( 
.A(n_5762),
.B(n_5218),
.Y(n_5865)
);

AND2x2_ASAP7_75t_L g5866 ( 
.A(n_5763),
.B(n_5665),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5748),
.Y(n_5867)
);

OR2x2_ASAP7_75t_L g5868 ( 
.A(n_5711),
.B(n_5531),
.Y(n_5868)
);

OR2x2_ASAP7_75t_L g5869 ( 
.A(n_5759),
.B(n_5511),
.Y(n_5869)
);

NOR2xp33_ASAP7_75t_L g5870 ( 
.A(n_5707),
.B(n_5125),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5700),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5710),
.Y(n_5872)
);

OR2x2_ASAP7_75t_L g5873 ( 
.A(n_5761),
.B(n_5772),
.Y(n_5873)
);

AND2x2_ASAP7_75t_L g5874 ( 
.A(n_5732),
.B(n_5334),
.Y(n_5874)
);

INVx2_ASAP7_75t_L g5875 ( 
.A(n_5742),
.Y(n_5875)
);

AND2x2_ASAP7_75t_L g5876 ( 
.A(n_5740),
.B(n_5787),
.Y(n_5876)
);

BUFx3_ASAP7_75t_L g5877 ( 
.A(n_5769),
.Y(n_5877)
);

OR2x2_ASAP7_75t_L g5878 ( 
.A(n_5729),
.B(n_4722),
.Y(n_5878)
);

AND2x2_ASAP7_75t_L g5879 ( 
.A(n_5694),
.B(n_5227),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5764),
.Y(n_5880)
);

AND2x4_ASAP7_75t_L g5881 ( 
.A(n_5745),
.B(n_5246),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_L g5882 ( 
.A(n_5713),
.B(n_5209),
.Y(n_5882)
);

NOR2xp67_ASAP7_75t_L g5883 ( 
.A(n_5734),
.B(n_5099),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5788),
.Y(n_5884)
);

AND2x4_ASAP7_75t_L g5885 ( 
.A(n_5795),
.B(n_5785),
.Y(n_5885)
);

INVx2_ASAP7_75t_L g5886 ( 
.A(n_5795),
.Y(n_5886)
);

NAND2xp5_ASAP7_75t_L g5887 ( 
.A(n_5804),
.B(n_5782),
.Y(n_5887)
);

AND2x4_ASAP7_75t_L g5888 ( 
.A(n_5799),
.B(n_5746),
.Y(n_5888)
);

AND2x2_ASAP7_75t_L g5889 ( 
.A(n_5845),
.B(n_5757),
.Y(n_5889)
);

AND2x2_ASAP7_75t_L g5890 ( 
.A(n_5845),
.B(n_5684),
.Y(n_5890)
);

AND2x2_ASAP7_75t_L g5891 ( 
.A(n_5834),
.B(n_5696),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5860),
.Y(n_5892)
);

NOR2xp33_ASAP7_75t_L g5893 ( 
.A(n_5797),
.B(n_5695),
.Y(n_5893)
);

AND2x4_ASAP7_75t_L g5894 ( 
.A(n_5834),
.B(n_5752),
.Y(n_5894)
);

OR2x2_ASAP7_75t_L g5895 ( 
.A(n_5878),
.B(n_5754),
.Y(n_5895)
);

NAND2xp5_ASAP7_75t_L g5896 ( 
.A(n_5813),
.B(n_5768),
.Y(n_5896)
);

AND2x4_ASAP7_75t_L g5897 ( 
.A(n_5815),
.B(n_5747),
.Y(n_5897)
);

INVx3_ASAP7_75t_L g5898 ( 
.A(n_5810),
.Y(n_5898)
);

INVx2_ASAP7_75t_L g5899 ( 
.A(n_5833),
.Y(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_5871),
.B(n_5720),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5833),
.Y(n_5901)
);

NAND2xp5_ASAP7_75t_L g5902 ( 
.A(n_5872),
.B(n_5725),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5867),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_L g5904 ( 
.A(n_5817),
.B(n_5726),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5844),
.B(n_5704),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5844),
.B(n_5705),
.Y(n_5906)
);

AND2x2_ASAP7_75t_L g5907 ( 
.A(n_5844),
.B(n_5703),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5819),
.B(n_5678),
.Y(n_5908)
);

NAND2xp5_ASAP7_75t_L g5909 ( 
.A(n_5864),
.B(n_5773),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5829),
.Y(n_5910)
);

INVx1_ASAP7_75t_L g5911 ( 
.A(n_5831),
.Y(n_5911)
);

NAND2xp5_ASAP7_75t_L g5912 ( 
.A(n_5801),
.B(n_5775),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5835),
.Y(n_5913)
);

BUFx2_ASAP7_75t_L g5914 ( 
.A(n_5815),
.Y(n_5914)
);

OR2x2_ASAP7_75t_L g5915 ( 
.A(n_5873),
.B(n_5715),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5836),
.Y(n_5916)
);

NAND2x1_ASAP7_75t_L g5917 ( 
.A(n_5803),
.B(n_5699),
.Y(n_5917)
);

AND2x2_ASAP7_75t_L g5918 ( 
.A(n_5805),
.B(n_5699),
.Y(n_5918)
);

HB1xp67_ASAP7_75t_L g5919 ( 
.A(n_5800),
.Y(n_5919)
);

AND2x2_ASAP7_75t_L g5920 ( 
.A(n_5807),
.B(n_5676),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5812),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5812),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5839),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5847),
.Y(n_5924)
);

INVx2_ASAP7_75t_L g5925 ( 
.A(n_5814),
.Y(n_5925)
);

AND2x4_ASAP7_75t_L g5926 ( 
.A(n_5808),
.B(n_5778),
.Y(n_5926)
);

NAND2xp5_ASAP7_75t_L g5927 ( 
.A(n_5868),
.B(n_5780),
.Y(n_5927)
);

AND2x2_ASAP7_75t_L g5928 ( 
.A(n_5796),
.B(n_5739),
.Y(n_5928)
);

BUFx3_ASAP7_75t_L g5929 ( 
.A(n_5810),
.Y(n_5929)
);

OR2x2_ASAP7_75t_L g5930 ( 
.A(n_5814),
.B(n_5789),
.Y(n_5930)
);

AND2x2_ASAP7_75t_L g5931 ( 
.A(n_5881),
.B(n_5750),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_5881),
.B(n_5791),
.Y(n_5932)
);

NAND2x1p5_ASAP7_75t_L g5933 ( 
.A(n_5841),
.B(n_5246),
.Y(n_5933)
);

INVx2_ASAP7_75t_L g5934 ( 
.A(n_5802),
.Y(n_5934)
);

OR2x2_ASAP7_75t_L g5935 ( 
.A(n_5798),
.B(n_5743),
.Y(n_5935)
);

AND2x2_ASAP7_75t_L g5936 ( 
.A(n_5821),
.B(n_5824),
.Y(n_5936)
);

BUFx3_ASAP7_75t_L g5937 ( 
.A(n_5803),
.Y(n_5937)
);

OR2x2_ASAP7_75t_L g5938 ( 
.A(n_5822),
.B(n_5743),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5816),
.Y(n_5939)
);

NAND2xp5_ASAP7_75t_L g5940 ( 
.A(n_5843),
.B(n_5786),
.Y(n_5940)
);

AND2x2_ASAP7_75t_L g5941 ( 
.A(n_5850),
.B(n_5728),
.Y(n_5941)
);

OR2x2_ASAP7_75t_L g5942 ( 
.A(n_5832),
.B(n_5744),
.Y(n_5942)
);

AND2x2_ASAP7_75t_L g5943 ( 
.A(n_5861),
.B(n_5790),
.Y(n_5943)
);

INVx2_ASAP7_75t_L g5944 ( 
.A(n_5806),
.Y(n_5944)
);

OAI21xp33_ASAP7_75t_L g5945 ( 
.A1(n_5827),
.A2(n_5820),
.B(n_5866),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5837),
.B(n_5716),
.Y(n_5946)
);

BUFx2_ASAP7_75t_SL g5947 ( 
.A(n_5883),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_5838),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5846),
.B(n_5744),
.Y(n_5949)
);

AND2x2_ASAP7_75t_L g5950 ( 
.A(n_5830),
.B(n_5719),
.Y(n_5950)
);

BUFx2_ASAP7_75t_L g5951 ( 
.A(n_5877),
.Y(n_5951)
);

AND2x4_ASAP7_75t_L g5952 ( 
.A(n_5856),
.B(n_5852),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_5826),
.B(n_5722),
.Y(n_5953)
);

NAND2xp5_ASAP7_75t_L g5954 ( 
.A(n_5848),
.B(n_5738),
.Y(n_5954)
);

AND2x2_ASAP7_75t_L g5955 ( 
.A(n_5825),
.B(n_5749),
.Y(n_5955)
);

AND2x2_ASAP7_75t_L g5956 ( 
.A(n_5828),
.B(n_5753),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5857),
.Y(n_5957)
);

AND2x2_ASAP7_75t_L g5958 ( 
.A(n_5842),
.B(n_5176),
.Y(n_5958)
);

AND2x2_ASAP7_75t_L g5959 ( 
.A(n_5842),
.B(n_5809),
.Y(n_5959)
);

AND2x2_ASAP7_75t_L g5960 ( 
.A(n_5818),
.B(n_5166),
.Y(n_5960)
);

INVx2_ASAP7_75t_L g5961 ( 
.A(n_5863),
.Y(n_5961)
);

INVx2_ASAP7_75t_L g5962 ( 
.A(n_5875),
.Y(n_5962)
);

AND2x2_ASAP7_75t_L g5963 ( 
.A(n_5876),
.B(n_5166),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5853),
.Y(n_5964)
);

HB1xp67_ASAP7_75t_L g5965 ( 
.A(n_5880),
.Y(n_5965)
);

BUFx2_ASAP7_75t_SL g5966 ( 
.A(n_5858),
.Y(n_5966)
);

AND2x2_ASAP7_75t_L g5967 ( 
.A(n_5823),
.B(n_5248),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5854),
.Y(n_5968)
);

NAND2xp5_ASAP7_75t_L g5969 ( 
.A(n_5859),
.B(n_5536),
.Y(n_5969)
);

INVx2_ASAP7_75t_L g5970 ( 
.A(n_5884),
.Y(n_5970)
);

INVx2_ASAP7_75t_L g5971 ( 
.A(n_5869),
.Y(n_5971)
);

AND2x2_ASAP7_75t_L g5972 ( 
.A(n_5855),
.B(n_5132),
.Y(n_5972)
);

AND2x2_ASAP7_75t_L g5973 ( 
.A(n_5879),
.B(n_5232),
.Y(n_5973)
);

AND2x2_ASAP7_75t_L g5974 ( 
.A(n_5874),
.B(n_5261),
.Y(n_5974)
);

AND2x2_ASAP7_75t_L g5975 ( 
.A(n_5840),
.B(n_5261),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5849),
.Y(n_5976)
);

NAND2x1p5_ASAP7_75t_L g5977 ( 
.A(n_5862),
.B(n_5117),
.Y(n_5977)
);

HB1xp67_ASAP7_75t_L g5978 ( 
.A(n_5811),
.Y(n_5978)
);

INVx3_ASAP7_75t_L g5979 ( 
.A(n_5840),
.Y(n_5979)
);

NAND2xp5_ASAP7_75t_L g5980 ( 
.A(n_5882),
.B(n_5151),
.Y(n_5980)
);

AND2x2_ASAP7_75t_L g5981 ( 
.A(n_5851),
.B(n_5253),
.Y(n_5981)
);

OR2x2_ASAP7_75t_L g5982 ( 
.A(n_5870),
.B(n_4991),
.Y(n_5982)
);

AND2x2_ASAP7_75t_L g5983 ( 
.A(n_5865),
.B(n_5253),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5860),
.Y(n_5984)
);

BUFx2_ASAP7_75t_L g5985 ( 
.A(n_5815),
.Y(n_5985)
);

AND2x2_ASAP7_75t_L g5986 ( 
.A(n_5845),
.B(n_5326),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5860),
.Y(n_5987)
);

AND2x2_ASAP7_75t_L g5988 ( 
.A(n_5914),
.B(n_5341),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5919),
.Y(n_5989)
);

INVx2_ASAP7_75t_L g5990 ( 
.A(n_5886),
.Y(n_5990)
);

AND2x2_ASAP7_75t_L g5991 ( 
.A(n_5985),
.B(n_5079),
.Y(n_5991)
);

NAND2xp5_ASAP7_75t_L g5992 ( 
.A(n_5969),
.B(n_5157),
.Y(n_5992)
);

OR2x2_ASAP7_75t_L g5993 ( 
.A(n_5895),
.B(n_4594),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5899),
.Y(n_5994)
);

NAND2x1p5_ASAP7_75t_L g5995 ( 
.A(n_5898),
.B(n_5120),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5901),
.Y(n_5996)
);

INVx2_ASAP7_75t_SL g5997 ( 
.A(n_5937),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5900),
.Y(n_5998)
);

OR2x2_ASAP7_75t_L g5999 ( 
.A(n_5976),
.B(n_4594),
.Y(n_5999)
);

OR2x2_ASAP7_75t_L g6000 ( 
.A(n_5976),
.B(n_4991),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5902),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5980),
.B(n_5185),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5912),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5890),
.B(n_5302),
.Y(n_6004)
);

NOR4xp75_ASAP7_75t_L g6005 ( 
.A(n_5898),
.B(n_5311),
.C(n_5346),
.D(n_5317),
.Y(n_6005)
);

INVx2_ASAP7_75t_L g6006 ( 
.A(n_5951),
.Y(n_6006)
);

INVxp67_ASAP7_75t_SL g6007 ( 
.A(n_5893),
.Y(n_6007)
);

BUFx2_ASAP7_75t_L g6008 ( 
.A(n_5929),
.Y(n_6008)
);

AND2x4_ASAP7_75t_L g6009 ( 
.A(n_5952),
.B(n_5885),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5921),
.Y(n_6010)
);

NAND2xp5_ASAP7_75t_L g6011 ( 
.A(n_5922),
.B(n_5230),
.Y(n_6011)
);

INVx1_ASAP7_75t_L g6012 ( 
.A(n_5925),
.Y(n_6012)
);

OR2x2_ASAP7_75t_L g6013 ( 
.A(n_5909),
.B(n_4904),
.Y(n_6013)
);

AND2x2_ASAP7_75t_L g6014 ( 
.A(n_5966),
.B(n_5133),
.Y(n_6014)
);

NAND2xp5_ASAP7_75t_L g6015 ( 
.A(n_5889),
.B(n_5221),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5904),
.Y(n_6016)
);

OR2x2_ASAP7_75t_L g6017 ( 
.A(n_5934),
.B(n_4904),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5965),
.Y(n_6018)
);

AND2x2_ASAP7_75t_L g6019 ( 
.A(n_5888),
.B(n_5086),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5927),
.Y(n_6020)
);

INVxp67_ASAP7_75t_L g6021 ( 
.A(n_5887),
.Y(n_6021)
);

NOR2xp33_ASAP7_75t_L g6022 ( 
.A(n_5947),
.B(n_5159),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5940),
.Y(n_6023)
);

HB1xp67_ASAP7_75t_L g6024 ( 
.A(n_5930),
.Y(n_6024)
);

NAND2xp5_ASAP7_75t_L g6025 ( 
.A(n_5888),
.B(n_5149),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5949),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5891),
.B(n_5936),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5892),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5952),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5928),
.Y(n_6030)
);

INVxp67_ASAP7_75t_L g6031 ( 
.A(n_5986),
.Y(n_6031)
);

NAND2xp5_ASAP7_75t_L g6032 ( 
.A(n_5982),
.B(n_5129),
.Y(n_6032)
);

O2A1O1Ixp5_ASAP7_75t_L g6033 ( 
.A1(n_5917),
.A2(n_5288),
.B(n_5348),
.C(n_5349),
.Y(n_6033)
);

INVx2_ASAP7_75t_L g6034 ( 
.A(n_5942),
.Y(n_6034)
);

INVxp67_ASAP7_75t_L g6035 ( 
.A(n_5896),
.Y(n_6035)
);

OR2x2_ASAP7_75t_L g6036 ( 
.A(n_5915),
.B(n_4945),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5892),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_5903),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_5903),
.Y(n_6039)
);

OR2x2_ASAP7_75t_L g6040 ( 
.A(n_5939),
.B(n_4945),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5975),
.B(n_5184),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5959),
.B(n_5268),
.Y(n_6042)
);

OR2x2_ASAP7_75t_L g6043 ( 
.A(n_5935),
.B(n_4962),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5910),
.Y(n_6044)
);

NOR2xp33_ASAP7_75t_L g6045 ( 
.A(n_5885),
.B(n_5160),
.Y(n_6045)
);

NOR2xp33_ASAP7_75t_L g6046 ( 
.A(n_5977),
.B(n_5144),
.Y(n_6046)
);

NAND2xp5_ASAP7_75t_L g6047 ( 
.A(n_5894),
.B(n_5308),
.Y(n_6047)
);

INVx1_ASAP7_75t_L g6048 ( 
.A(n_5910),
.Y(n_6048)
);

AND2x2_ASAP7_75t_L g6049 ( 
.A(n_5972),
.B(n_5113),
.Y(n_6049)
);

NOR2xp67_ASAP7_75t_L g6050 ( 
.A(n_5897),
.B(n_720),
.Y(n_6050)
);

AND2x2_ASAP7_75t_L g6051 ( 
.A(n_5897),
.B(n_5115),
.Y(n_6051)
);

OR2x2_ASAP7_75t_L g6052 ( 
.A(n_5938),
.B(n_5954),
.Y(n_6052)
);

NAND4xp75_ASAP7_75t_L g6053 ( 
.A(n_5941),
.B(n_5286),
.C(n_4787),
.D(n_4938),
.Y(n_6053)
);

INVx1_ASAP7_75t_L g6054 ( 
.A(n_5911),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_5944),
.Y(n_6055)
);

AND2x4_ASAP7_75t_L g6056 ( 
.A(n_5983),
.B(n_5155),
.Y(n_6056)
);

NOR2x1p5_ASAP7_75t_L g6057 ( 
.A(n_5979),
.B(n_5894),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5953),
.Y(n_6058)
);

NAND2xp5_ASAP7_75t_L g6059 ( 
.A(n_5956),
.B(n_5180),
.Y(n_6059)
);

NOR2xp33_ASAP7_75t_L g6060 ( 
.A(n_5958),
.B(n_5225),
.Y(n_6060)
);

AOI21xp5_ASAP7_75t_L g6061 ( 
.A1(n_5933),
.A2(n_5225),
.B(n_5001),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5911),
.Y(n_6062)
);

NAND2xp5_ASAP7_75t_L g6063 ( 
.A(n_5970),
.B(n_5075),
.Y(n_6063)
);

AND2x2_ASAP7_75t_L g6064 ( 
.A(n_5907),
.B(n_5095),
.Y(n_6064)
);

NAND2x1p5_ASAP7_75t_L g6065 ( 
.A(n_5974),
.B(n_5054),
.Y(n_6065)
);

INVxp67_ASAP7_75t_L g6066 ( 
.A(n_5926),
.Y(n_6066)
);

AND2x2_ASAP7_75t_L g6067 ( 
.A(n_5932),
.B(n_4907),
.Y(n_6067)
);

INVx2_ASAP7_75t_L g6068 ( 
.A(n_5948),
.Y(n_6068)
);

NAND2xp33_ASAP7_75t_SL g6069 ( 
.A(n_6008),
.B(n_5991),
.Y(n_6069)
);

OAI22xp33_ASAP7_75t_L g6070 ( 
.A1(n_6004),
.A2(n_5979),
.B1(n_5971),
.B2(n_5978),
.Y(n_6070)
);

OAI22xp5_ASAP7_75t_L g6071 ( 
.A1(n_6066),
.A2(n_5997),
.B1(n_6031),
.B2(n_6006),
.Y(n_6071)
);

INVx2_ASAP7_75t_L g6072 ( 
.A(n_6029),
.Y(n_6072)
);

NAND2xp5_ASAP7_75t_L g6073 ( 
.A(n_6007),
.B(n_5943),
.Y(n_6073)
);

AO221x2_ASAP7_75t_L g6074 ( 
.A1(n_5995),
.A2(n_5945),
.B1(n_5913),
.B2(n_5924),
.C(n_5923),
.Y(n_6074)
);

NAND2xp5_ASAP7_75t_L g6075 ( 
.A(n_6050),
.B(n_5926),
.Y(n_6075)
);

NOR2xp33_ASAP7_75t_L g6076 ( 
.A(n_6022),
.B(n_6015),
.Y(n_6076)
);

INVxp67_ASAP7_75t_L g6077 ( 
.A(n_6014),
.Y(n_6077)
);

NOR2xp33_ASAP7_75t_L g6078 ( 
.A(n_6009),
.B(n_5973),
.Y(n_6078)
);

NAND2xp5_ASAP7_75t_L g6079 ( 
.A(n_6035),
.B(n_5916),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_6024),
.Y(n_6080)
);

AND2x2_ASAP7_75t_L g6081 ( 
.A(n_6027),
.B(n_5908),
.Y(n_6081)
);

INVx4_ASAP7_75t_L g6082 ( 
.A(n_6056),
.Y(n_6082)
);

INVx3_ASAP7_75t_L g6083 ( 
.A(n_6056),
.Y(n_6083)
);

NAND2xp5_ASAP7_75t_L g6084 ( 
.A(n_5989),
.B(n_6021),
.Y(n_6084)
);

OAI221xp5_ASAP7_75t_L g6085 ( 
.A1(n_6033),
.A2(n_5918),
.B1(n_5905),
.B2(n_5906),
.C(n_5916),
.Y(n_6085)
);

INVxp67_ASAP7_75t_L g6086 ( 
.A(n_5989),
.Y(n_6086)
);

NAND2xp5_ASAP7_75t_L g6087 ( 
.A(n_5992),
.B(n_5913),
.Y(n_6087)
);

NOR2xp33_ASAP7_75t_L g6088 ( 
.A(n_6009),
.B(n_5960),
.Y(n_6088)
);

NAND2xp5_ASAP7_75t_L g6089 ( 
.A(n_6030),
.B(n_5923),
.Y(n_6089)
);

OAI221xp5_ASAP7_75t_L g6090 ( 
.A1(n_6065),
.A2(n_5924),
.B1(n_5984),
.B2(n_5968),
.C(n_5964),
.Y(n_6090)
);

AO221x2_ASAP7_75t_L g6091 ( 
.A1(n_6047),
.A2(n_5984),
.B1(n_5987),
.B2(n_5968),
.C(n_5964),
.Y(n_6091)
);

AOI22xp5_ASAP7_75t_L g6092 ( 
.A1(n_6051),
.A2(n_5987),
.B1(n_5931),
.B2(n_5963),
.Y(n_6092)
);

AO221x2_ASAP7_75t_L g6093 ( 
.A1(n_6032),
.A2(n_5957),
.B1(n_5962),
.B2(n_5961),
.C(n_5300),
.Y(n_6093)
);

AOI22xp5_ASAP7_75t_L g6094 ( 
.A1(n_6002),
.A2(n_5967),
.B1(n_5981),
.B2(n_5955),
.Y(n_6094)
);

NAND2xp5_ASAP7_75t_L g6095 ( 
.A(n_5998),
.B(n_6001),
.Y(n_6095)
);

INVx2_ASAP7_75t_L g6096 ( 
.A(n_5990),
.Y(n_6096)
);

NOR2xp67_ASAP7_75t_L g6097 ( 
.A(n_5994),
.B(n_5920),
.Y(n_6097)
);

NAND2xp5_ASAP7_75t_L g6098 ( 
.A(n_6016),
.B(n_5946),
.Y(n_6098)
);

OAI22xp33_ASAP7_75t_L g6099 ( 
.A1(n_6025),
.A2(n_5950),
.B1(n_5249),
.B2(n_5372),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_6019),
.B(n_5260),
.Y(n_6100)
);

NAND2xp5_ASAP7_75t_L g6101 ( 
.A(n_6023),
.B(n_5219),
.Y(n_6101)
);

NAND2xp33_ASAP7_75t_SL g6102 ( 
.A(n_6057),
.B(n_5988),
.Y(n_6102)
);

NAND2xp5_ASAP7_75t_L g6103 ( 
.A(n_6026),
.B(n_5211),
.Y(n_6103)
);

OAI22xp33_ASAP7_75t_L g6104 ( 
.A1(n_6052),
.A2(n_5249),
.B1(n_5370),
.B2(n_5022),
.Y(n_6104)
);

OAI221xp5_ASAP7_75t_L g6105 ( 
.A1(n_6018),
.A2(n_5278),
.B1(n_5272),
.B2(n_5212),
.C(n_5290),
.Y(n_6105)
);

NAND2xp5_ASAP7_75t_L g6106 ( 
.A(n_6020),
.B(n_5351),
.Y(n_6106)
);

NAND2xp5_ASAP7_75t_L g6107 ( 
.A(n_6003),
.B(n_5114),
.Y(n_6107)
);

NOR2xp33_ASAP7_75t_SL g6108 ( 
.A(n_6046),
.B(n_4931),
.Y(n_6108)
);

AOI22xp5_ASAP7_75t_L g6109 ( 
.A1(n_6064),
.A2(n_5332),
.B1(n_5333),
.B2(n_5375),
.Y(n_6109)
);

OAI221xp5_ASAP7_75t_L g6110 ( 
.A1(n_5996),
.A2(n_5222),
.B1(n_5303),
.B2(n_5369),
.C(n_5359),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_6067),
.B(n_5148),
.Y(n_6111)
);

NAND2xp5_ASAP7_75t_L g6112 ( 
.A(n_6010),
.B(n_4877),
.Y(n_6112)
);

NAND2xp5_ASAP7_75t_L g6113 ( 
.A(n_6012),
.B(n_6011),
.Y(n_6113)
);

NAND2xp5_ASAP7_75t_L g6114 ( 
.A(n_6063),
.B(n_4880),
.Y(n_6114)
);

NAND2xp5_ASAP7_75t_L g6115 ( 
.A(n_6034),
.B(n_4921),
.Y(n_6115)
);

INVxp67_ASAP7_75t_L g6116 ( 
.A(n_6045),
.Y(n_6116)
);

NAND2xp33_ASAP7_75t_SL g6117 ( 
.A(n_6041),
.B(n_5336),
.Y(n_6117)
);

OAI22xp33_ASAP7_75t_L g6118 ( 
.A1(n_6059),
.A2(n_6036),
.B1(n_6058),
.B2(n_6013),
.Y(n_6118)
);

AOI22xp5_ASAP7_75t_L g6119 ( 
.A1(n_6053),
.A2(n_5097),
.B1(n_5109),
.B2(n_5047),
.Y(n_6119)
);

AND2x2_ASAP7_75t_L g6120 ( 
.A(n_6049),
.B(n_4907),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_L g6121 ( 
.A(n_6055),
.B(n_4927),
.Y(n_6121)
);

NAND2xp5_ASAP7_75t_L g6122 ( 
.A(n_6068),
.B(n_4948),
.Y(n_6122)
);

AO221x2_ASAP7_75t_L g6123 ( 
.A1(n_6028),
.A2(n_5014),
.B1(n_4878),
.B2(n_4896),
.C(n_4892),
.Y(n_6123)
);

INVxp67_ASAP7_75t_L g6124 ( 
.A(n_6042),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_6043),
.B(n_4950),
.Y(n_6125)
);

NOR2xp33_ASAP7_75t_L g6126 ( 
.A(n_6060),
.B(n_6037),
.Y(n_6126)
);

NOR2xp67_ASAP7_75t_SL g6127 ( 
.A(n_6082),
.B(n_6083),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_6072),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_6080),
.Y(n_6129)
);

INVx1_ASAP7_75t_SL g6130 ( 
.A(n_6069),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_6096),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_6077),
.Y(n_6132)
);

AND2x2_ASAP7_75t_L g6133 ( 
.A(n_6076),
.B(n_5993),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_6124),
.Y(n_6134)
);

INVx2_ASAP7_75t_SL g6135 ( 
.A(n_6078),
.Y(n_6135)
);

OR2x2_ASAP7_75t_L g6136 ( 
.A(n_6084),
.B(n_6040),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_6113),
.Y(n_6137)
);

NAND2xp5_ASAP7_75t_L g6138 ( 
.A(n_6071),
.B(n_6000),
.Y(n_6138)
);

NOR2xp33_ASAP7_75t_L g6139 ( 
.A(n_6116),
.B(n_6038),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_6121),
.Y(n_6140)
);

NAND2xp5_ASAP7_75t_L g6141 ( 
.A(n_6100),
.B(n_6039),
.Y(n_6141)
);

AND2x2_ASAP7_75t_SL g6142 ( 
.A(n_6075),
.B(n_6028),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_6098),
.Y(n_6143)
);

INVx3_ASAP7_75t_L g6144 ( 
.A(n_6074),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_6122),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_6086),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_6073),
.Y(n_6147)
);

HB1xp67_ASAP7_75t_L g6148 ( 
.A(n_6095),
.Y(n_6148)
);

AND2x2_ASAP7_75t_L g6149 ( 
.A(n_6081),
.B(n_6044),
.Y(n_6149)
);

BUFx2_ASAP7_75t_L g6150 ( 
.A(n_6102),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_6107),
.Y(n_6151)
);

AND2x2_ASAP7_75t_L g6152 ( 
.A(n_6088),
.B(n_6048),
.Y(n_6152)
);

NAND2xp5_ASAP7_75t_L g6153 ( 
.A(n_6119),
.B(n_6054),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_6097),
.B(n_6062),
.Y(n_6154)
);

AND2x2_ASAP7_75t_L g6155 ( 
.A(n_6094),
.B(n_6017),
.Y(n_6155)
);

INVx1_ASAP7_75t_SL g6156 ( 
.A(n_6112),
.Y(n_6156)
);

AND2x4_ASAP7_75t_L g6157 ( 
.A(n_6126),
.B(n_6061),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_6089),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_6115),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_6114),
.Y(n_6160)
);

AND2x2_ASAP7_75t_L g6161 ( 
.A(n_6092),
.B(n_5999),
.Y(n_6161)
);

AOI21xp33_ASAP7_75t_SL g6162 ( 
.A1(n_6070),
.A2(n_722),
.B(n_723),
.Y(n_6162)
);

AOI22xp5_ASAP7_75t_L g6163 ( 
.A1(n_6117),
.A2(n_6005),
.B1(n_4614),
.B2(n_4724),
.Y(n_6163)
);

AOI22xp5_ASAP7_75t_L g6164 ( 
.A1(n_6108),
.A2(n_4965),
.B1(n_4826),
.B2(n_4814),
.Y(n_6164)
);

AOI22xp33_ASAP7_75t_L g6165 ( 
.A1(n_6093),
.A2(n_4879),
.B1(n_4745),
.B2(n_4846),
.Y(n_6165)
);

INVxp67_ASAP7_75t_L g6166 ( 
.A(n_6085),
.Y(n_6166)
);

OAI22xp5_ASAP7_75t_L g6167 ( 
.A1(n_6111),
.A2(n_4851),
.B1(n_4728),
.B2(n_4812),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_6079),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_6125),
.Y(n_6169)
);

NAND2xp5_ASAP7_75t_L g6170 ( 
.A(n_6120),
.B(n_722),
.Y(n_6170)
);

NOR2xp33_ASAP7_75t_L g6171 ( 
.A(n_6087),
.B(n_723),
.Y(n_6171)
);

NAND2xp5_ASAP7_75t_L g6172 ( 
.A(n_6118),
.B(n_723),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_6106),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_6074),
.B(n_4962),
.Y(n_6174)
);

INVxp67_ASAP7_75t_L g6175 ( 
.A(n_6101),
.Y(n_6175)
);

NAND2xp5_ASAP7_75t_L g6176 ( 
.A(n_6091),
.B(n_6103),
.Y(n_6176)
);

AOI21xp5_ASAP7_75t_SL g6177 ( 
.A1(n_6093),
.A2(n_4784),
.B(n_4783),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_6123),
.Y(n_6178)
);

NAND2x2_ASAP7_75t_L g6179 ( 
.A(n_6099),
.B(n_724),
.Y(n_6179)
);

AND2x2_ASAP7_75t_L g6180 ( 
.A(n_6091),
.B(n_4977),
.Y(n_6180)
);

OR2x2_ASAP7_75t_L g6181 ( 
.A(n_6123),
.B(n_724),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_6104),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_6090),
.Y(n_6183)
);

O2A1O1Ixp33_ASAP7_75t_L g6184 ( 
.A1(n_6105),
.A2(n_4917),
.B(n_4715),
.C(n_4712),
.Y(n_6184)
);

INVxp67_ASAP7_75t_L g6185 ( 
.A(n_6110),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_6109),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_6072),
.Y(n_6187)
);

HB1xp67_ASAP7_75t_L g6188 ( 
.A(n_6080),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_6072),
.Y(n_6189)
);

INVx2_ASAP7_75t_SL g6190 ( 
.A(n_6132),
.Y(n_6190)
);

OAI22xp5_ASAP7_75t_L g6191 ( 
.A1(n_6166),
.A2(n_4864),
.B1(n_4866),
.B2(n_4766),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_6128),
.Y(n_6192)
);

NAND2xp5_ASAP7_75t_L g6193 ( 
.A(n_6163),
.B(n_724),
.Y(n_6193)
);

OA21x2_ASAP7_75t_L g6194 ( 
.A1(n_6172),
.A2(n_4849),
.B(n_4845),
.Y(n_6194)
);

OAI21xp33_ASAP7_75t_SL g6195 ( 
.A1(n_6144),
.A2(n_4785),
.B(n_4763),
.Y(n_6195)
);

AOI22xp5_ASAP7_75t_L g6196 ( 
.A1(n_6127),
.A2(n_4705),
.B1(n_4664),
.B2(n_4725),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_6187),
.Y(n_6197)
);

INVx2_ASAP7_75t_L g6198 ( 
.A(n_6189),
.Y(n_6198)
);

AOI22xp33_ASAP7_75t_L g6199 ( 
.A1(n_6150),
.A2(n_4860),
.B1(n_4739),
.B2(n_4757),
.Y(n_6199)
);

AOI21xp5_ASAP7_75t_L g6200 ( 
.A1(n_6130),
.A2(n_4747),
.B(n_4713),
.Y(n_6200)
);

INVx2_ASAP7_75t_L g6201 ( 
.A(n_6131),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_6188),
.Y(n_6202)
);

INVx2_ASAP7_75t_L g6203 ( 
.A(n_6134),
.Y(n_6203)
);

NAND2xp5_ASAP7_75t_L g6204 ( 
.A(n_6185),
.B(n_725),
.Y(n_6204)
);

AOI22xp5_ASAP7_75t_L g6205 ( 
.A1(n_6182),
.A2(n_4618),
.B1(n_4750),
.B2(n_4706),
.Y(n_6205)
);

OAI21xp33_ASAP7_75t_L g6206 ( 
.A1(n_6135),
.A2(n_4609),
.B(n_4798),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_6186),
.B(n_725),
.Y(n_6207)
);

INVx2_ASAP7_75t_SL g6208 ( 
.A(n_6157),
.Y(n_6208)
);

AOI22xp5_ASAP7_75t_L g6209 ( 
.A1(n_6157),
.A2(n_4822),
.B1(n_4841),
.B2(n_4802),
.Y(n_6209)
);

O2A1O1Ixp5_ASAP7_75t_L g6210 ( 
.A1(n_6144),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_6210)
);

AOI22xp5_ASAP7_75t_L g6211 ( 
.A1(n_6179),
.A2(n_4887),
.B1(n_4906),
.B2(n_4856),
.Y(n_6211)
);

OAI21xp33_ASAP7_75t_L g6212 ( 
.A1(n_6183),
.A2(n_4978),
.B(n_4926),
.Y(n_6212)
);

NOR3xp33_ASAP7_75t_L g6213 ( 
.A(n_6162),
.B(n_726),
.C(n_727),
.Y(n_6213)
);

OAI31xp33_ASAP7_75t_L g6214 ( 
.A1(n_6178),
.A2(n_4876),
.A3(n_4977),
.B(n_5049),
.Y(n_6214)
);

AOI221xp5_ASAP7_75t_L g6215 ( 
.A1(n_6139),
.A2(n_730),
.B1(n_728),
.B2(n_729),
.C(n_731),
.Y(n_6215)
);

NOR2xp33_ASAP7_75t_SL g6216 ( 
.A(n_6147),
.B(n_6129),
.Y(n_6216)
);

A2O1A1Ixp33_ASAP7_75t_L g6217 ( 
.A1(n_6138),
.A2(n_5007),
.B(n_5011),
.C(n_5008),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_6181),
.Y(n_6218)
);

AOI22xp5_ASAP7_75t_L g6219 ( 
.A1(n_6133),
.A2(n_4971),
.B1(n_5028),
.B2(n_4891),
.Y(n_6219)
);

OAI22xp5_ASAP7_75t_L g6220 ( 
.A1(n_6165),
.A2(n_5028),
.B1(n_4891),
.B2(n_5049),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_L g6221 ( 
.A(n_6156),
.B(n_729),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_6149),
.Y(n_6222)
);

OR2x2_ASAP7_75t_L g6223 ( 
.A(n_6141),
.B(n_6170),
.Y(n_6223)
);

NAND2xp5_ASAP7_75t_L g6224 ( 
.A(n_6173),
.B(n_729),
.Y(n_6224)
);

NAND2xp33_ASAP7_75t_SL g6225 ( 
.A(n_6148),
.B(n_6153),
.Y(n_6225)
);

A2O1A1Ixp33_ASAP7_75t_L g6226 ( 
.A1(n_6175),
.A2(n_732),
.B(n_730),
.C(n_731),
.Y(n_6226)
);

AND2x2_ASAP7_75t_L g6227 ( 
.A(n_6152),
.B(n_731),
.Y(n_6227)
);

AOI22xp5_ASAP7_75t_L g6228 ( 
.A1(n_6143),
.A2(n_5057),
.B1(n_734),
.B2(n_732),
.Y(n_6228)
);

NAND2xp5_ASAP7_75t_L g6229 ( 
.A(n_6151),
.B(n_732),
.Y(n_6229)
);

AOI22xp5_ASAP7_75t_L g6230 ( 
.A1(n_6155),
.A2(n_5057),
.B1(n_735),
.B2(n_733),
.Y(n_6230)
);

OAI22xp5_ASAP7_75t_L g6231 ( 
.A1(n_6176),
.A2(n_735),
.B1(n_733),
.B2(n_734),
.Y(n_6231)
);

NAND2xp5_ASAP7_75t_L g6232 ( 
.A(n_6137),
.B(n_735),
.Y(n_6232)
);

OAI22xp33_ASAP7_75t_L g6233 ( 
.A1(n_6136),
.A2(n_4983),
.B1(n_738),
.B2(n_736),
.Y(n_6233)
);

NAND2xp5_ASAP7_75t_L g6234 ( 
.A(n_6171),
.B(n_736),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_6140),
.Y(n_6235)
);

INVx1_ASAP7_75t_SL g6236 ( 
.A(n_6146),
.Y(n_6236)
);

NAND2xp5_ASAP7_75t_L g6237 ( 
.A(n_6145),
.B(n_736),
.Y(n_6237)
);

INVx1_ASAP7_75t_SL g6238 ( 
.A(n_6159),
.Y(n_6238)
);

OAI22xp5_ASAP7_75t_L g6239 ( 
.A1(n_6168),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.Y(n_6239)
);

AOI311xp33_ASAP7_75t_L g6240 ( 
.A1(n_6169),
.A2(n_740),
.A3(n_737),
.B(n_739),
.C(n_741),
.Y(n_6240)
);

O2A1O1Ixp33_ASAP7_75t_L g6241 ( 
.A1(n_6158),
.A2(n_741),
.B(n_737),
.C(n_739),
.Y(n_6241)
);

NAND2xp5_ASAP7_75t_L g6242 ( 
.A(n_6160),
.B(n_742),
.Y(n_6242)
);

NAND4xp25_ASAP7_75t_L g6243 ( 
.A(n_6177),
.B(n_744),
.C(n_742),
.D(n_743),
.Y(n_6243)
);

INVx3_ASAP7_75t_L g6244 ( 
.A(n_6154),
.Y(n_6244)
);

INVx2_ASAP7_75t_SL g6245 ( 
.A(n_6142),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_6158),
.Y(n_6246)
);

AOI211xp5_ASAP7_75t_SL g6247 ( 
.A1(n_6174),
.A2(n_745),
.B(n_743),
.C(n_744),
.Y(n_6247)
);

INVx1_ASAP7_75t_L g6248 ( 
.A(n_6180),
.Y(n_6248)
);

AND2x2_ASAP7_75t_L g6249 ( 
.A(n_6161),
.B(n_743),
.Y(n_6249)
);

AND2x2_ASAP7_75t_L g6250 ( 
.A(n_6218),
.B(n_6164),
.Y(n_6250)
);

NOR2xp67_ASAP7_75t_SL g6251 ( 
.A(n_6208),
.B(n_744),
.Y(n_6251)
);

OR2x2_ASAP7_75t_L g6252 ( 
.A(n_6190),
.B(n_6207),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_6203),
.Y(n_6253)
);

NOR2xp33_ASAP7_75t_L g6254 ( 
.A(n_6243),
.B(n_6184),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_6221),
.Y(n_6255)
);

OAI21xp33_ASAP7_75t_L g6256 ( 
.A1(n_6204),
.A2(n_6167),
.B(n_745),
.Y(n_6256)
);

NAND2xp5_ASAP7_75t_L g6257 ( 
.A(n_6213),
.B(n_745),
.Y(n_6257)
);

NOR2xp33_ASAP7_75t_L g6258 ( 
.A(n_6244),
.B(n_746),
.Y(n_6258)
);

AOI21xp33_ASAP7_75t_L g6259 ( 
.A1(n_6231),
.A2(n_746),
.B(n_747),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_6247),
.B(n_6244),
.Y(n_6260)
);

NAND3xp33_ASAP7_75t_L g6261 ( 
.A(n_6210),
.B(n_746),
.C(n_747),
.Y(n_6261)
);

AOI21xp33_ASAP7_75t_SL g6262 ( 
.A1(n_6193),
.A2(n_747),
.B(n_748),
.Y(n_6262)
);

NOR2xp67_ASAP7_75t_L g6263 ( 
.A(n_6198),
.B(n_748),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_6201),
.Y(n_6264)
);

AOI221x1_ASAP7_75t_L g6265 ( 
.A1(n_6225),
.A2(n_750),
.B1(n_748),
.B2(n_749),
.C(n_751),
.Y(n_6265)
);

NOR2xp33_ASAP7_75t_L g6266 ( 
.A(n_6216),
.B(n_749),
.Y(n_6266)
);

NAND2xp5_ASAP7_75t_L g6267 ( 
.A(n_6249),
.B(n_749),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_6227),
.Y(n_6268)
);

OAI21xp5_ASAP7_75t_SL g6269 ( 
.A1(n_6236),
.A2(n_750),
.B(n_751),
.Y(n_6269)
);

OAI21xp33_ASAP7_75t_L g6270 ( 
.A1(n_6222),
.A2(n_750),
.B(n_751),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_6202),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_6192),
.Y(n_6272)
);

O2A1O1Ixp5_ASAP7_75t_L g6273 ( 
.A1(n_6197),
.A2(n_755),
.B(n_752),
.C(n_753),
.Y(n_6273)
);

INVxp67_ASAP7_75t_L g6274 ( 
.A(n_6234),
.Y(n_6274)
);

OAI221xp5_ASAP7_75t_L g6275 ( 
.A1(n_6212),
.A2(n_755),
.B1(n_752),
.B2(n_753),
.C(n_756),
.Y(n_6275)
);

AOI21xp5_ASAP7_75t_L g6276 ( 
.A1(n_6232),
.A2(n_6229),
.B(n_6224),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_6235),
.Y(n_6277)
);

AND2x4_ASAP7_75t_L g6278 ( 
.A(n_6238),
.B(n_752),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_6237),
.Y(n_6279)
);

OR2x2_ASAP7_75t_L g6280 ( 
.A(n_6242),
.B(n_753),
.Y(n_6280)
);

OAI22xp5_ASAP7_75t_L g6281 ( 
.A1(n_6245),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.Y(n_6281)
);

AOI22xp5_ASAP7_75t_L g6282 ( 
.A1(n_6248),
.A2(n_6230),
.B1(n_6239),
.B2(n_6223),
.Y(n_6282)
);

OR2x2_ASAP7_75t_L g6283 ( 
.A(n_6226),
.B(n_757),
.Y(n_6283)
);

AOI22xp33_ASAP7_75t_SL g6284 ( 
.A1(n_6246),
.A2(n_6195),
.B1(n_6194),
.B2(n_6191),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6194),
.Y(n_6285)
);

INVx1_ASAP7_75t_L g6286 ( 
.A(n_6241),
.Y(n_6286)
);

OAI32xp33_ASAP7_75t_L g6287 ( 
.A1(n_6220),
.A2(n_759),
.A3(n_757),
.B1(n_758),
.B2(n_760),
.Y(n_6287)
);

INVx2_ASAP7_75t_L g6288 ( 
.A(n_6205),
.Y(n_6288)
);

NOR2xp33_ASAP7_75t_L g6289 ( 
.A(n_6233),
.B(n_758),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_6219),
.Y(n_6290)
);

A2O1A1Ixp33_ASAP7_75t_L g6291 ( 
.A1(n_6215),
.A2(n_761),
.B(n_759),
.C(n_760),
.Y(n_6291)
);

AOI322xp5_ASAP7_75t_L g6292 ( 
.A1(n_6199),
.A2(n_4983),
.A3(n_761),
.B1(n_762),
.B2(n_763),
.C1(n_764),
.C2(n_765),
.Y(n_6292)
);

NOR3xp33_ASAP7_75t_L g6293 ( 
.A(n_6206),
.B(n_759),
.C(n_761),
.Y(n_6293)
);

AOI221xp5_ASAP7_75t_L g6294 ( 
.A1(n_6217),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.C(n_765),
.Y(n_6294)
);

HB1xp67_ASAP7_75t_L g6295 ( 
.A(n_6200),
.Y(n_6295)
);

NAND3xp33_ASAP7_75t_L g6296 ( 
.A(n_6240),
.B(n_763),
.C(n_764),
.Y(n_6296)
);

NOR2xp33_ASAP7_75t_L g6297 ( 
.A(n_6228),
.B(n_765),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_6211),
.Y(n_6298)
);

O2A1O1Ixp5_ASAP7_75t_L g6299 ( 
.A1(n_6214),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_6299)
);

OR2x2_ASAP7_75t_L g6300 ( 
.A(n_6209),
.B(n_766),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_6196),
.Y(n_6301)
);

NAND2xp5_ASAP7_75t_L g6302 ( 
.A(n_6218),
.B(n_767),
.Y(n_6302)
);

AOI22xp33_ASAP7_75t_L g6303 ( 
.A1(n_6208),
.A2(n_769),
.B1(n_767),
.B2(n_768),
.Y(n_6303)
);

OAI22xp33_ASAP7_75t_L g6304 ( 
.A1(n_6243),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_6304)
);

AOI21xp5_ASAP7_75t_L g6305 ( 
.A1(n_6204),
.A2(n_769),
.B(n_770),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6190),
.Y(n_6306)
);

AOI22xp5_ASAP7_75t_L g6307 ( 
.A1(n_6218),
.A2(n_773),
.B1(n_771),
.B2(n_772),
.Y(n_6307)
);

NAND2xp5_ASAP7_75t_L g6308 ( 
.A(n_6218),
.B(n_772),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_6190),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_6190),
.Y(n_6310)
);

AOI22xp5_ASAP7_75t_L g6311 ( 
.A1(n_6218),
.A2(n_774),
.B1(n_772),
.B2(n_773),
.Y(n_6311)
);

OA22x2_ASAP7_75t_L g6312 ( 
.A1(n_6208),
.A2(n_775),
.B1(n_773),
.B2(n_774),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_6190),
.Y(n_6313)
);

O2A1O1Ixp33_ASAP7_75t_SL g6314 ( 
.A1(n_6218),
.A2(n_776),
.B(n_774),
.C(n_775),
.Y(n_6314)
);

NAND2xp5_ASAP7_75t_L g6315 ( 
.A(n_6218),
.B(n_777),
.Y(n_6315)
);

AOI32xp33_ASAP7_75t_L g6316 ( 
.A1(n_6225),
.A2(n_779),
.A3(n_777),
.B1(n_778),
.B2(n_780),
.Y(n_6316)
);

OAI21xp33_ASAP7_75t_L g6317 ( 
.A1(n_6204),
.A2(n_778),
.B(n_779),
.Y(n_6317)
);

INVxp67_ASAP7_75t_SL g6318 ( 
.A(n_6207),
.Y(n_6318)
);

INVx2_ASAP7_75t_L g6319 ( 
.A(n_6208),
.Y(n_6319)
);

AOI22xp5_ASAP7_75t_L g6320 ( 
.A1(n_6218),
.A2(n_780),
.B1(n_778),
.B2(n_779),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_6190),
.Y(n_6321)
);

NAND2xp5_ASAP7_75t_L g6322 ( 
.A(n_6218),
.B(n_780),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_6190),
.Y(n_6323)
);

INVx1_ASAP7_75t_L g6324 ( 
.A(n_6190),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6190),
.Y(n_6325)
);

OAI22xp33_ASAP7_75t_L g6326 ( 
.A1(n_6243),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.Y(n_6326)
);

OAI22xp33_ASAP7_75t_L g6327 ( 
.A1(n_6243),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.Y(n_6327)
);

AOI22xp5_ASAP7_75t_L g6328 ( 
.A1(n_6218),
.A2(n_784),
.B1(n_781),
.B2(n_783),
.Y(n_6328)
);

OAI22xp33_ASAP7_75t_SL g6329 ( 
.A1(n_6218),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.Y(n_6329)
);

AOI322xp5_ASAP7_75t_L g6330 ( 
.A1(n_6254),
.A2(n_784),
.A3(n_785),
.B1(n_786),
.B2(n_787),
.C1(n_788),
.C2(n_789),
.Y(n_6330)
);

OAI21xp5_ASAP7_75t_L g6331 ( 
.A1(n_6299),
.A2(n_785),
.B(n_786),
.Y(n_6331)
);

AND2x2_ASAP7_75t_L g6332 ( 
.A(n_6319),
.B(n_787),
.Y(n_6332)
);

AOI221xp5_ASAP7_75t_L g6333 ( 
.A1(n_6287),
.A2(n_789),
.B1(n_787),
.B2(n_788),
.C(n_790),
.Y(n_6333)
);

OAI21xp5_ASAP7_75t_L g6334 ( 
.A1(n_6261),
.A2(n_788),
.B(n_789),
.Y(n_6334)
);

OAI211xp5_ASAP7_75t_L g6335 ( 
.A1(n_6256),
.A2(n_792),
.B(n_790),
.C(n_791),
.Y(n_6335)
);

OAI211xp5_ASAP7_75t_L g6336 ( 
.A1(n_6306),
.A2(n_793),
.B(n_791),
.C(n_792),
.Y(n_6336)
);

OAI22xp5_ASAP7_75t_L g6337 ( 
.A1(n_6309),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.Y(n_6337)
);

NAND2xp5_ASAP7_75t_L g6338 ( 
.A(n_6251),
.B(n_6278),
.Y(n_6338)
);

OAI22xp5_ASAP7_75t_L g6339 ( 
.A1(n_6310),
.A2(n_795),
.B1(n_793),
.B2(n_794),
.Y(n_6339)
);

OAI22xp5_ASAP7_75t_L g6340 ( 
.A1(n_6313),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_6340)
);

AOI22xp33_ASAP7_75t_L g6341 ( 
.A1(n_6321),
.A2(n_797),
.B1(n_795),
.B2(n_796),
.Y(n_6341)
);

OAI21xp33_ASAP7_75t_L g6342 ( 
.A1(n_6260),
.A2(n_796),
.B(n_797),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_6312),
.Y(n_6343)
);

OAI211xp5_ASAP7_75t_SL g6344 ( 
.A1(n_6323),
.A2(n_799),
.B(n_797),
.C(n_798),
.Y(n_6344)
);

NOR2x1_ASAP7_75t_L g6345 ( 
.A(n_6324),
.B(n_798),
.Y(n_6345)
);

OA21x2_ASAP7_75t_L g6346 ( 
.A1(n_6325),
.A2(n_800),
.B(n_801),
.Y(n_6346)
);

AOI31xp33_ASAP7_75t_L g6347 ( 
.A1(n_6286),
.A2(n_802),
.A3(n_800),
.B(n_801),
.Y(n_6347)
);

AOI322xp5_ASAP7_75t_L g6348 ( 
.A1(n_6250),
.A2(n_801),
.A3(n_802),
.B1(n_803),
.B2(n_804),
.C1(n_806),
.C2(n_807),
.Y(n_6348)
);

AOI322xp5_ASAP7_75t_L g6349 ( 
.A1(n_6253),
.A2(n_802),
.A3(n_803),
.B1(n_804),
.B2(n_807),
.C1(n_808),
.C2(n_809),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_6264),
.Y(n_6350)
);

OAI21xp33_ASAP7_75t_L g6351 ( 
.A1(n_6282),
.A2(n_6308),
.B(n_6302),
.Y(n_6351)
);

NAND2xp5_ASAP7_75t_SL g6352 ( 
.A(n_6329),
.B(n_803),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6278),
.Y(n_6353)
);

AOI221xp5_ASAP7_75t_L g6354 ( 
.A1(n_6277),
.A2(n_808),
.B1(n_804),
.B2(n_807),
.C(n_809),
.Y(n_6354)
);

AOI22xp33_ASAP7_75t_L g6355 ( 
.A1(n_6293),
.A2(n_811),
.B1(n_809),
.B2(n_810),
.Y(n_6355)
);

AOI222xp33_ASAP7_75t_L g6356 ( 
.A1(n_6298),
.A2(n_812),
.B1(n_814),
.B2(n_810),
.C1(n_811),
.C2(n_813),
.Y(n_6356)
);

AOI22xp5_ASAP7_75t_L g6357 ( 
.A1(n_6304),
.A2(n_812),
.B1(n_810),
.B2(n_811),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_6314),
.Y(n_6358)
);

OAI21xp5_ASAP7_75t_L g6359 ( 
.A1(n_6269),
.A2(n_812),
.B(n_813),
.Y(n_6359)
);

AOI332xp33_ASAP7_75t_L g6360 ( 
.A1(n_6271),
.A2(n_814),
.A3(n_815),
.B1(n_816),
.B2(n_817),
.B3(n_818),
.C1(n_819),
.C2(n_820),
.Y(n_6360)
);

AOI221xp5_ASAP7_75t_L g6361 ( 
.A1(n_6275),
.A2(n_6259),
.B1(n_6294),
.B2(n_6327),
.C(n_6326),
.Y(n_6361)
);

AND2x4_ASAP7_75t_L g6362 ( 
.A(n_6263),
.B(n_814),
.Y(n_6362)
);

AOI32xp33_ASAP7_75t_L g6363 ( 
.A1(n_6284),
.A2(n_817),
.A3(n_815),
.B1(n_816),
.B2(n_818),
.Y(n_6363)
);

NAND2xp5_ASAP7_75t_L g6364 ( 
.A(n_6266),
.B(n_815),
.Y(n_6364)
);

AOI21xp5_ASAP7_75t_L g6365 ( 
.A1(n_6315),
.A2(n_6322),
.B(n_6281),
.Y(n_6365)
);

OAI22xp5_ASAP7_75t_L g6366 ( 
.A1(n_6307),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.Y(n_6366)
);

NOR2x1_ASAP7_75t_L g6367 ( 
.A(n_6258),
.B(n_819),
.Y(n_6367)
);

AOI22xp5_ASAP7_75t_L g6368 ( 
.A1(n_6289),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.Y(n_6368)
);

A2O1A1Ixp33_ASAP7_75t_L g6369 ( 
.A1(n_6316),
.A2(n_822),
.B(n_820),
.C(n_821),
.Y(n_6369)
);

INVx2_ASAP7_75t_L g6370 ( 
.A(n_6252),
.Y(n_6370)
);

AOI221x1_ASAP7_75t_L g6371 ( 
.A1(n_6272),
.A2(n_824),
.B1(n_822),
.B2(n_823),
.C(n_825),
.Y(n_6371)
);

O2A1O1Ixp33_ASAP7_75t_L g6372 ( 
.A1(n_6291),
.A2(n_6273),
.B(n_6262),
.C(n_6257),
.Y(n_6372)
);

AOI221xp5_ASAP7_75t_L g6373 ( 
.A1(n_6268),
.A2(n_824),
.B1(n_822),
.B2(n_823),
.C(n_825),
.Y(n_6373)
);

A2O1A1Ixp33_ASAP7_75t_L g6374 ( 
.A1(n_6305),
.A2(n_825),
.B(n_823),
.C(n_824),
.Y(n_6374)
);

AOI22xp5_ASAP7_75t_L g6375 ( 
.A1(n_6270),
.A2(n_829),
.B1(n_826),
.B2(n_828),
.Y(n_6375)
);

NOR4xp25_ASAP7_75t_L g6376 ( 
.A(n_6255),
.B(n_829),
.C(n_826),
.D(n_828),
.Y(n_6376)
);

O2A1O1Ixp5_ASAP7_75t_L g6377 ( 
.A1(n_6318),
.A2(n_830),
.B(n_828),
.C(n_829),
.Y(n_6377)
);

OAI221xp5_ASAP7_75t_L g6378 ( 
.A1(n_6317),
.A2(n_6328),
.B1(n_6320),
.B2(n_6311),
.C(n_6303),
.Y(n_6378)
);

OAI22xp5_ASAP7_75t_L g6379 ( 
.A1(n_6288),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_6379)
);

OAI211xp5_ASAP7_75t_L g6380 ( 
.A1(n_6265),
.A2(n_833),
.B(n_831),
.C(n_832),
.Y(n_6380)
);

NOR2xp33_ASAP7_75t_L g6381 ( 
.A(n_6267),
.B(n_832),
.Y(n_6381)
);

OAI221xp5_ASAP7_75t_L g6382 ( 
.A1(n_6296),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.C(n_836),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6280),
.Y(n_6383)
);

OAI21xp5_ASAP7_75t_L g6384 ( 
.A1(n_6276),
.A2(n_834),
.B(n_835),
.Y(n_6384)
);

OAI21xp33_ASAP7_75t_SL g6385 ( 
.A1(n_6290),
.A2(n_834),
.B(n_835),
.Y(n_6385)
);

AOI22xp5_ASAP7_75t_L g6386 ( 
.A1(n_6297),
.A2(n_6301),
.B1(n_6274),
.B2(n_6279),
.Y(n_6386)
);

AOI22xp5_ASAP7_75t_L g6387 ( 
.A1(n_6283),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_6387)
);

INVx2_ASAP7_75t_SL g6388 ( 
.A(n_6300),
.Y(n_6388)
);

AND2x2_ASAP7_75t_L g6389 ( 
.A(n_6295),
.B(n_837),
.Y(n_6389)
);

AOI211xp5_ASAP7_75t_SL g6390 ( 
.A1(n_6285),
.A2(n_6292),
.B(n_839),
.C(n_837),
.Y(n_6390)
);

NOR4xp25_ASAP7_75t_L g6391 ( 
.A(n_6306),
.B(n_840),
.C(n_838),
.D(n_839),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6343),
.Y(n_6392)
);

INVx2_ASAP7_75t_L g6393 ( 
.A(n_6350),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_6346),
.Y(n_6394)
);

BUFx2_ASAP7_75t_L g6395 ( 
.A(n_6346),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_6370),
.Y(n_6396)
);

INVxp67_ASAP7_75t_L g6397 ( 
.A(n_6332),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_6358),
.Y(n_6398)
);

INVx1_ASAP7_75t_SL g6399 ( 
.A(n_6338),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6345),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_6353),
.Y(n_6401)
);

NAND2xp5_ASAP7_75t_SL g6402 ( 
.A(n_6363),
.B(n_6356),
.Y(n_6402)
);

INVx1_ASAP7_75t_SL g6403 ( 
.A(n_6389),
.Y(n_6403)
);

BUFx2_ASAP7_75t_L g6404 ( 
.A(n_6331),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_6347),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6364),
.Y(n_6406)
);

NOR2xp33_ASAP7_75t_L g6407 ( 
.A(n_6382),
.B(n_838),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_6337),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_6339),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6340),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6334),
.B(n_840),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_6362),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_6362),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6379),
.Y(n_6414)
);

HB1xp67_ASAP7_75t_L g6415 ( 
.A(n_6388),
.Y(n_6415)
);

INVx2_ASAP7_75t_L g6416 ( 
.A(n_6383),
.Y(n_6416)
);

INVx1_ASAP7_75t_L g6417 ( 
.A(n_6352),
.Y(n_6417)
);

HB1xp67_ASAP7_75t_L g6418 ( 
.A(n_6359),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_6357),
.Y(n_6419)
);

INVx2_ASAP7_75t_L g6420 ( 
.A(n_6377),
.Y(n_6420)
);

INVx2_ASAP7_75t_SL g6421 ( 
.A(n_6367),
.Y(n_6421)
);

INVx2_ASAP7_75t_L g6422 ( 
.A(n_6375),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_6387),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6342),
.Y(n_6424)
);

INVx2_ASAP7_75t_L g6425 ( 
.A(n_6368),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6336),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_6381),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6371),
.Y(n_6428)
);

INVx8_ASAP7_75t_L g6429 ( 
.A(n_6386),
.Y(n_6429)
);

BUFx12f_ASAP7_75t_L g6430 ( 
.A(n_6391),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6366),
.Y(n_6431)
);

BUFx4f_ASAP7_75t_SL g6432 ( 
.A(n_6384),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_6380),
.Y(n_6433)
);

INVxp33_ASAP7_75t_SL g6434 ( 
.A(n_6341),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6335),
.Y(n_6435)
);

HB1xp67_ASAP7_75t_L g6436 ( 
.A(n_6385),
.Y(n_6436)
);

INVx2_ASAP7_75t_L g6437 ( 
.A(n_6378),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_6369),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6344),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6360),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6374),
.Y(n_6441)
);

INVx2_ASAP7_75t_SL g6442 ( 
.A(n_6348),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_6372),
.Y(n_6443)
);

INVx2_ASAP7_75t_L g6444 ( 
.A(n_6349),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6351),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6333),
.Y(n_6446)
);

BUFx12f_ASAP7_75t_L g6447 ( 
.A(n_6361),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_6394),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6394),
.Y(n_6449)
);

NOR2xp67_ASAP7_75t_L g6450 ( 
.A(n_6398),
.B(n_6365),
.Y(n_6450)
);

NOR2xp33_ASAP7_75t_L g6451 ( 
.A(n_6436),
.B(n_6355),
.Y(n_6451)
);

AOI21xp33_ASAP7_75t_SL g6452 ( 
.A1(n_6426),
.A2(n_6376),
.B(n_6390),
.Y(n_6452)
);

NOR3x1_ASAP7_75t_L g6453 ( 
.A(n_6442),
.B(n_6373),
.C(n_6354),
.Y(n_6453)
);

AND2x2_ASAP7_75t_L g6454 ( 
.A(n_6396),
.B(n_6330),
.Y(n_6454)
);

NAND4xp25_ASAP7_75t_L g6455 ( 
.A(n_6399),
.B(n_843),
.C(n_840),
.D(n_842),
.Y(n_6455)
);

NAND3xp33_ASAP7_75t_L g6456 ( 
.A(n_6392),
.B(n_842),
.C(n_843),
.Y(n_6456)
);

NOR3xp33_ASAP7_75t_L g6457 ( 
.A(n_6392),
.B(n_843),
.C(n_844),
.Y(n_6457)
);

NOR2xp67_ASAP7_75t_L g6458 ( 
.A(n_6437),
.B(n_844),
.Y(n_6458)
);

NAND4xp25_ASAP7_75t_L g6459 ( 
.A(n_6433),
.B(n_848),
.C(n_846),
.D(n_847),
.Y(n_6459)
);

NOR2x1_ASAP7_75t_L g6460 ( 
.A(n_6443),
.B(n_6393),
.Y(n_6460)
);

NAND4xp25_ASAP7_75t_L g6461 ( 
.A(n_6435),
.B(n_849),
.C(n_846),
.D(n_848),
.Y(n_6461)
);

AOI22xp33_ASAP7_75t_L g6462 ( 
.A1(n_6447),
.A2(n_850),
.B1(n_846),
.B2(n_849),
.Y(n_6462)
);

NOR3xp33_ASAP7_75t_L g6463 ( 
.A(n_6445),
.B(n_850),
.C(n_851),
.Y(n_6463)
);

NOR2x1_ASAP7_75t_L g6464 ( 
.A(n_6420),
.B(n_6428),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6415),
.Y(n_6465)
);

NOR2x1_ASAP7_75t_L g6466 ( 
.A(n_6405),
.B(n_850),
.Y(n_6466)
);

AND2x2_ASAP7_75t_L g6467 ( 
.A(n_6411),
.B(n_852),
.Y(n_6467)
);

NOR2x2_ASAP7_75t_L g6468 ( 
.A(n_6440),
.B(n_852),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_6412),
.Y(n_6469)
);

NOR2x1_ASAP7_75t_L g6470 ( 
.A(n_6401),
.B(n_853),
.Y(n_6470)
);

HB1xp67_ASAP7_75t_L g6471 ( 
.A(n_6413),
.Y(n_6471)
);

AOI22xp5_ASAP7_75t_L g6472 ( 
.A1(n_6434),
.A2(n_855),
.B1(n_853),
.B2(n_854),
.Y(n_6472)
);

HB1xp67_ASAP7_75t_L g6473 ( 
.A(n_6417),
.Y(n_6473)
);

OAI22xp33_ASAP7_75t_L g6474 ( 
.A1(n_6432),
.A2(n_856),
.B1(n_854),
.B2(n_855),
.Y(n_6474)
);

XNOR2x2_ASAP7_75t_L g6475 ( 
.A(n_6407),
.B(n_854),
.Y(n_6475)
);

OA21x2_ASAP7_75t_L g6476 ( 
.A1(n_6395),
.A2(n_856),
.B(n_857),
.Y(n_6476)
);

NAND3xp33_ASAP7_75t_L g6477 ( 
.A(n_6444),
.B(n_6424),
.C(n_6446),
.Y(n_6477)
);

AOI21xp5_ASAP7_75t_L g6478 ( 
.A1(n_6402),
.A2(n_856),
.B(n_857),
.Y(n_6478)
);

NAND3xp33_ASAP7_75t_L g6479 ( 
.A(n_6446),
.B(n_858),
.C(n_859),
.Y(n_6479)
);

NAND4xp75_ASAP7_75t_L g6480 ( 
.A(n_6439),
.B(n_860),
.C(n_858),
.D(n_859),
.Y(n_6480)
);

INVxp67_ASAP7_75t_SL g6481 ( 
.A(n_6416),
.Y(n_6481)
);

NAND2x1_ASAP7_75t_SL g6482 ( 
.A(n_6418),
.B(n_858),
.Y(n_6482)
);

OAI211xp5_ASAP7_75t_L g6483 ( 
.A1(n_6429),
.A2(n_861),
.B(n_859),
.C(n_860),
.Y(n_6483)
);

NAND3xp33_ASAP7_75t_L g6484 ( 
.A(n_6438),
.B(n_860),
.C(n_861),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6404),
.Y(n_6485)
);

OAI21xp5_ASAP7_75t_L g6486 ( 
.A1(n_6397),
.A2(n_862),
.B(n_863),
.Y(n_6486)
);

NAND4xp25_ASAP7_75t_SL g6487 ( 
.A(n_6403),
.B(n_865),
.C(n_862),
.D(n_864),
.Y(n_6487)
);

NOR2x1p5_ASAP7_75t_SL g6488 ( 
.A(n_6441),
.B(n_6422),
.Y(n_6488)
);

AND2x2_ASAP7_75t_SL g6489 ( 
.A(n_6400),
.B(n_862),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_6429),
.Y(n_6490)
);

NAND3xp33_ASAP7_75t_L g6491 ( 
.A(n_6408),
.B(n_864),
.C(n_865),
.Y(n_6491)
);

AOI211xp5_ASAP7_75t_L g6492 ( 
.A1(n_6409),
.A2(n_867),
.B(n_864),
.C(n_866),
.Y(n_6492)
);

AO22x2_ASAP7_75t_L g6493 ( 
.A1(n_6410),
.A2(n_868),
.B1(n_866),
.B2(n_867),
.Y(n_6493)
);

OAI21xp33_ASAP7_75t_SL g6494 ( 
.A1(n_6414),
.A2(n_866),
.B(n_868),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6419),
.Y(n_6495)
);

OAI22xp5_ASAP7_75t_L g6496 ( 
.A1(n_6477),
.A2(n_6431),
.B1(n_6425),
.B2(n_6423),
.Y(n_6496)
);

NAND2xp5_ASAP7_75t_L g6497 ( 
.A(n_6448),
.B(n_6421),
.Y(n_6497)
);

NAND3xp33_ASAP7_75t_SL g6498 ( 
.A(n_6492),
.B(n_6406),
.C(n_6427),
.Y(n_6498)
);

NAND4xp25_ASAP7_75t_L g6499 ( 
.A(n_6453),
.B(n_6451),
.C(n_6490),
.D(n_6462),
.Y(n_6499)
);

AND2x2_ASAP7_75t_L g6500 ( 
.A(n_6465),
.B(n_6430),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6449),
.Y(n_6501)
);

NAND4xp25_ASAP7_75t_L g6502 ( 
.A(n_6478),
.B(n_871),
.C(n_869),
.D(n_870),
.Y(n_6502)
);

NOR2x1_ASAP7_75t_L g6503 ( 
.A(n_6491),
.B(n_869),
.Y(n_6503)
);

AOI21xp5_ASAP7_75t_L g6504 ( 
.A1(n_6481),
.A2(n_6464),
.B(n_6487),
.Y(n_6504)
);

NOR2xp33_ASAP7_75t_L g6505 ( 
.A(n_6494),
.B(n_870),
.Y(n_6505)
);

NOR2x1_ASAP7_75t_L g6506 ( 
.A(n_6479),
.B(n_870),
.Y(n_6506)
);

NOR5xp2_ASAP7_75t_L g6507 ( 
.A(n_6473),
.B(n_873),
.C(n_871),
.D(n_872),
.E(n_874),
.Y(n_6507)
);

AOI21xp5_ASAP7_75t_L g6508 ( 
.A1(n_6493),
.A2(n_871),
.B(n_872),
.Y(n_6508)
);

NOR4xp25_ASAP7_75t_L g6509 ( 
.A(n_6495),
.B(n_875),
.C(n_873),
.D(n_874),
.Y(n_6509)
);

NOR2x1_ASAP7_75t_L g6510 ( 
.A(n_6456),
.B(n_873),
.Y(n_6510)
);

CKINVDCx16_ASAP7_75t_R g6511 ( 
.A(n_6472),
.Y(n_6511)
);

AOI221xp5_ASAP7_75t_L g6512 ( 
.A1(n_6452),
.A2(n_876),
.B1(n_874),
.B2(n_875),
.C(n_877),
.Y(n_6512)
);

NOR2x1_ASAP7_75t_L g6513 ( 
.A(n_6484),
.B(n_875),
.Y(n_6513)
);

NAND4xp25_ASAP7_75t_SL g6514 ( 
.A(n_6454),
.B(n_878),
.C(n_876),
.D(n_877),
.Y(n_6514)
);

NOR3xp33_ASAP7_75t_SL g6515 ( 
.A(n_6461),
.B(n_876),
.C(n_879),
.Y(n_6515)
);

NOR2x1_ASAP7_75t_L g6516 ( 
.A(n_6460),
.B(n_879),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_6493),
.Y(n_6517)
);

NOR3xp33_ASAP7_75t_L g6518 ( 
.A(n_6483),
.B(n_879),
.C(n_880),
.Y(n_6518)
);

OAI21xp5_ASAP7_75t_L g6519 ( 
.A1(n_6458),
.A2(n_880),
.B(n_881),
.Y(n_6519)
);

AND4x2_ASAP7_75t_L g6520 ( 
.A(n_6466),
.B(n_884),
.C(n_882),
.D(n_883),
.Y(n_6520)
);

NOR4xp25_ASAP7_75t_L g6521 ( 
.A(n_6469),
.B(n_884),
.C(n_882),
.D(n_883),
.Y(n_6521)
);

NAND4xp25_ASAP7_75t_L g6522 ( 
.A(n_6459),
.B(n_885),
.C(n_882),
.D(n_884),
.Y(n_6522)
);

NAND3xp33_ASAP7_75t_SL g6523 ( 
.A(n_6463),
.B(n_885),
.C(n_886),
.Y(n_6523)
);

NOR3xp33_ASAP7_75t_L g6524 ( 
.A(n_6455),
.B(n_886),
.C(n_887),
.Y(n_6524)
);

NAND2xp5_ASAP7_75t_SL g6525 ( 
.A(n_6457),
.B(n_886),
.Y(n_6525)
);

NOR3x1_ASAP7_75t_L g6526 ( 
.A(n_6480),
.B(n_887),
.C(n_888),
.Y(n_6526)
);

NOR2x1_ASAP7_75t_L g6527 ( 
.A(n_6470),
.B(n_888),
.Y(n_6527)
);

A2O1A1Ixp33_ASAP7_75t_SL g6528 ( 
.A1(n_6485),
.A2(n_890),
.B(n_888),
.C(n_889),
.Y(n_6528)
);

AOI221xp5_ASAP7_75t_L g6529 ( 
.A1(n_6474),
.A2(n_890),
.B1(n_891),
.B2(n_892),
.C(n_893),
.Y(n_6529)
);

OAI211xp5_ASAP7_75t_SL g6530 ( 
.A1(n_6486),
.A2(n_892),
.B(n_890),
.C(n_891),
.Y(n_6530)
);

OAI21xp5_ASAP7_75t_L g6531 ( 
.A1(n_6450),
.A2(n_891),
.B(n_892),
.Y(n_6531)
);

NAND4xp25_ASAP7_75t_SL g6532 ( 
.A(n_6467),
.B(n_895),
.C(n_893),
.D(n_894),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6471),
.Y(n_6533)
);

OAI211xp5_ASAP7_75t_L g6534 ( 
.A1(n_6482),
.A2(n_895),
.B(n_893),
.C(n_894),
.Y(n_6534)
);

NAND4xp25_ASAP7_75t_L g6535 ( 
.A(n_6499),
.B(n_6488),
.C(n_6475),
.D(n_6468),
.Y(n_6535)
);

NOR3xp33_ASAP7_75t_SL g6536 ( 
.A(n_6496),
.B(n_6489),
.C(n_6476),
.Y(n_6536)
);

AOI22xp33_ASAP7_75t_L g6537 ( 
.A1(n_6514),
.A2(n_6476),
.B1(n_897),
.B2(n_894),
.Y(n_6537)
);

NOR3xp33_ASAP7_75t_L g6538 ( 
.A(n_6512),
.B(n_896),
.C(n_897),
.Y(n_6538)
);

NAND4xp25_ASAP7_75t_L g6539 ( 
.A(n_6524),
.B(n_899),
.C(n_896),
.D(n_898),
.Y(n_6539)
);

NAND2xp5_ASAP7_75t_SL g6540 ( 
.A(n_6509),
.B(n_898),
.Y(n_6540)
);

OR3x1_ASAP7_75t_L g6541 ( 
.A(n_6522),
.B(n_6523),
.C(n_6532),
.Y(n_6541)
);

NOR2x1p5_ASAP7_75t_L g6542 ( 
.A(n_6533),
.B(n_899),
.Y(n_6542)
);

NOR4xp25_ASAP7_75t_L g6543 ( 
.A(n_6498),
.B(n_902),
.C(n_900),
.D(n_901),
.Y(n_6543)
);

NAND3xp33_ASAP7_75t_L g6544 ( 
.A(n_6529),
.B(n_900),
.C(n_901),
.Y(n_6544)
);

AOI221xp5_ASAP7_75t_L g6545 ( 
.A1(n_6521),
.A2(n_901),
.B1(n_902),
.B2(n_903),
.C(n_904),
.Y(n_6545)
);

NOR2x1_ASAP7_75t_L g6546 ( 
.A(n_6516),
.B(n_902),
.Y(n_6546)
);

NAND2xp5_ASAP7_75t_L g6547 ( 
.A(n_6505),
.B(n_903),
.Y(n_6547)
);

NAND4xp25_ASAP7_75t_SL g6548 ( 
.A(n_6518),
.B(n_905),
.C(n_903),
.D(n_904),
.Y(n_6548)
);

A2O1A1Ixp33_ASAP7_75t_L g6549 ( 
.A1(n_6504),
.A2(n_906),
.B(n_904),
.C(n_905),
.Y(n_6549)
);

NAND3xp33_ASAP7_75t_SL g6550 ( 
.A(n_6507),
.B(n_906),
.C(n_907),
.Y(n_6550)
);

AND3x2_ASAP7_75t_L g6551 ( 
.A(n_6531),
.B(n_906),
.C(n_907),
.Y(n_6551)
);

NOR5xp2_ASAP7_75t_L g6552 ( 
.A(n_6534),
.B(n_908),
.C(n_909),
.D(n_910),
.E(n_911),
.Y(n_6552)
);

OR5x1_ASAP7_75t_L g6553 ( 
.A(n_6502),
.B(n_908),
.C(n_909),
.D(n_910),
.E(n_911),
.Y(n_6553)
);

NAND3xp33_ASAP7_75t_SL g6554 ( 
.A(n_6497),
.B(n_908),
.C(n_909),
.Y(n_6554)
);

NAND2xp5_ASAP7_75t_L g6555 ( 
.A(n_6517),
.B(n_910),
.Y(n_6555)
);

NOR2x1_ASAP7_75t_L g6556 ( 
.A(n_6527),
.B(n_912),
.Y(n_6556)
);

AOI322xp5_ASAP7_75t_L g6557 ( 
.A1(n_6500),
.A2(n_912),
.A3(n_913),
.B1(n_914),
.B2(n_915),
.C1(n_916),
.C2(n_917),
.Y(n_6557)
);

AOI211xp5_ASAP7_75t_L g6558 ( 
.A1(n_6530),
.A2(n_914),
.B(n_912),
.C(n_913),
.Y(n_6558)
);

NAND2xp5_ASAP7_75t_L g6559 ( 
.A(n_6508),
.B(n_913),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6503),
.Y(n_6560)
);

OAI211xp5_ASAP7_75t_L g6561 ( 
.A1(n_6528),
.A2(n_916),
.B(n_914),
.C(n_915),
.Y(n_6561)
);

OAI211xp5_ASAP7_75t_L g6562 ( 
.A1(n_6515),
.A2(n_918),
.B(n_915),
.C(n_917),
.Y(n_6562)
);

NOR2x1_ASAP7_75t_L g6563 ( 
.A(n_6535),
.B(n_6501),
.Y(n_6563)
);

INVx1_ASAP7_75t_L g6564 ( 
.A(n_6555),
.Y(n_6564)
);

NOR3xp33_ASAP7_75t_L g6565 ( 
.A(n_6554),
.B(n_6525),
.C(n_6511),
.Y(n_6565)
);

AND3x4_ASAP7_75t_L g6566 ( 
.A(n_6538),
.B(n_6513),
.C(n_6510),
.Y(n_6566)
);

AOI22xp33_ASAP7_75t_L g6567 ( 
.A1(n_6548),
.A2(n_6506),
.B1(n_6519),
.B2(n_6520),
.Y(n_6567)
);

NOR2x1_ASAP7_75t_L g6568 ( 
.A(n_6550),
.B(n_6526),
.Y(n_6568)
);

AOI22xp5_ASAP7_75t_L g6569 ( 
.A1(n_6541),
.A2(n_919),
.B1(n_917),
.B2(n_918),
.Y(n_6569)
);

OAI22xp5_ASAP7_75t_L g6570 ( 
.A1(n_6537),
.A2(n_920),
.B1(n_918),
.B2(n_919),
.Y(n_6570)
);

XOR2xp5_ASAP7_75t_L g6571 ( 
.A(n_6539),
.B(n_919),
.Y(n_6571)
);

NAND2xp5_ASAP7_75t_L g6572 ( 
.A(n_6557),
.B(n_920),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6559),
.Y(n_6573)
);

INVx2_ASAP7_75t_L g6574 ( 
.A(n_6542),
.Y(n_6574)
);

AND2x4_ASAP7_75t_L g6575 ( 
.A(n_6560),
.B(n_922),
.Y(n_6575)
);

NOR2x1p5_ASAP7_75t_L g6576 ( 
.A(n_6547),
.B(n_922),
.Y(n_6576)
);

NAND3xp33_ASAP7_75t_L g6577 ( 
.A(n_6536),
.B(n_923),
.C(n_924),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_6546),
.Y(n_6578)
);

NOR2x1_ASAP7_75t_L g6579 ( 
.A(n_6540),
.B(n_923),
.Y(n_6579)
);

HB1xp67_ASAP7_75t_L g6580 ( 
.A(n_6556),
.Y(n_6580)
);

OR2x2_ASAP7_75t_L g6581 ( 
.A(n_6543),
.B(n_923),
.Y(n_6581)
);

NOR3xp33_ASAP7_75t_L g6582 ( 
.A(n_6562),
.B(n_924),
.C(n_925),
.Y(n_6582)
);

INVx2_ASAP7_75t_L g6583 ( 
.A(n_6551),
.Y(n_6583)
);

AOI32xp33_ASAP7_75t_L g6584 ( 
.A1(n_6558),
.A2(n_925),
.A3(n_926),
.B1(n_927),
.B2(n_928),
.Y(n_6584)
);

AND2x2_ASAP7_75t_L g6585 ( 
.A(n_6549),
.B(n_925),
.Y(n_6585)
);

AND2x2_ASAP7_75t_L g6586 ( 
.A(n_6545),
.B(n_926),
.Y(n_6586)
);

AND3x2_ASAP7_75t_L g6587 ( 
.A(n_6552),
.B(n_926),
.C(n_927),
.Y(n_6587)
);

AND2x4_ASAP7_75t_L g6588 ( 
.A(n_6583),
.B(n_6544),
.Y(n_6588)
);

AND2x4_ASAP7_75t_L g6589 ( 
.A(n_6563),
.B(n_6553),
.Y(n_6589)
);

AND4x1_ASAP7_75t_L g6590 ( 
.A(n_6568),
.B(n_6577),
.C(n_6565),
.D(n_6579),
.Y(n_6590)
);

OR2x2_ASAP7_75t_L g6591 ( 
.A(n_6581),
.B(n_6561),
.Y(n_6591)
);

OR2x2_ASAP7_75t_L g6592 ( 
.A(n_6572),
.B(n_927),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6575),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6575),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6571),
.Y(n_6595)
);

NAND2xp5_ASAP7_75t_SL g6596 ( 
.A(n_6569),
.B(n_928),
.Y(n_6596)
);

NOR3xp33_ASAP7_75t_L g6597 ( 
.A(n_6570),
.B(n_928),
.C(n_929),
.Y(n_6597)
);

INVx2_ASAP7_75t_L g6598 ( 
.A(n_6587),
.Y(n_6598)
);

OR2x2_ASAP7_75t_L g6599 ( 
.A(n_6586),
.B(n_929),
.Y(n_6599)
);

AND2x4_ASAP7_75t_L g6600 ( 
.A(n_6574),
.B(n_929),
.Y(n_6600)
);

AND3x4_ASAP7_75t_L g6601 ( 
.A(n_6582),
.B(n_930),
.C(n_931),
.Y(n_6601)
);

INVx1_ASAP7_75t_L g6602 ( 
.A(n_6585),
.Y(n_6602)
);

BUFx2_ASAP7_75t_L g6603 ( 
.A(n_6564),
.Y(n_6603)
);

NAND3x1_ASAP7_75t_L g6604 ( 
.A(n_6573),
.B(n_930),
.C(n_931),
.Y(n_6604)
);

NOR3xp33_ASAP7_75t_L g6605 ( 
.A(n_6578),
.B(n_930),
.C(n_931),
.Y(n_6605)
);

NOR3xp33_ASAP7_75t_SL g6606 ( 
.A(n_6566),
.B(n_932),
.C(n_933),
.Y(n_6606)
);

NOR3xp33_ASAP7_75t_SL g6607 ( 
.A(n_6584),
.B(n_932),
.C(n_933),
.Y(n_6607)
);

NAND4xp25_ASAP7_75t_L g6608 ( 
.A(n_6567),
.B(n_936),
.C(n_933),
.D(n_934),
.Y(n_6608)
);

AND4x1_ASAP7_75t_L g6609 ( 
.A(n_6606),
.B(n_6576),
.C(n_6580),
.D(n_937),
.Y(n_6609)
);

INVxp67_ASAP7_75t_SL g6610 ( 
.A(n_6604),
.Y(n_6610)
);

AOI22xp5_ASAP7_75t_L g6611 ( 
.A1(n_6601),
.A2(n_937),
.B1(n_934),
.B2(n_936),
.Y(n_6611)
);

AOI21xp5_ASAP7_75t_L g6612 ( 
.A1(n_6596),
.A2(n_936),
.B(n_937),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_6591),
.Y(n_6613)
);

OAI22xp5_ASAP7_75t_L g6614 ( 
.A1(n_6592),
.A2(n_940),
.B1(n_938),
.B2(n_939),
.Y(n_6614)
);

NAND4xp75_ASAP7_75t_L g6615 ( 
.A(n_6595),
.B(n_940),
.C(n_938),
.D(n_939),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6600),
.B(n_941),
.Y(n_6616)
);

AOI31xp33_ASAP7_75t_L g6617 ( 
.A1(n_6593),
.A2(n_943),
.A3(n_941),
.B(n_942),
.Y(n_6617)
);

NAND2xp5_ASAP7_75t_L g6618 ( 
.A(n_6605),
.B(n_941),
.Y(n_6618)
);

AO211x2_ASAP7_75t_L g6619 ( 
.A1(n_6608),
.A2(n_6597),
.B(n_6594),
.C(n_6602),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6599),
.Y(n_6620)
);

AOI22xp5_ASAP7_75t_L g6621 ( 
.A1(n_6613),
.A2(n_6588),
.B1(n_6598),
.B2(n_6589),
.Y(n_6621)
);

OAI22xp5_ASAP7_75t_L g6622 ( 
.A1(n_6616),
.A2(n_6618),
.B1(n_6611),
.B2(n_6610),
.Y(n_6622)
);

AOI22xp5_ASAP7_75t_L g6623 ( 
.A1(n_6620),
.A2(n_6614),
.B1(n_6619),
.B2(n_6603),
.Y(n_6623)
);

INVxp67_ASAP7_75t_SL g6624 ( 
.A(n_6612),
.Y(n_6624)
);

INVx2_ASAP7_75t_L g6625 ( 
.A(n_6615),
.Y(n_6625)
);

AOI22xp33_ASAP7_75t_SL g6626 ( 
.A1(n_6609),
.A2(n_6590),
.B1(n_6607),
.B2(n_944),
.Y(n_6626)
);

HB1xp67_ASAP7_75t_L g6627 ( 
.A(n_6617),
.Y(n_6627)
);

AOI22xp5_ASAP7_75t_L g6628 ( 
.A1(n_6613),
.A2(n_944),
.B1(n_942),
.B2(n_943),
.Y(n_6628)
);

AOI22xp5_ASAP7_75t_L g6629 ( 
.A1(n_6613),
.A2(n_946),
.B1(n_942),
.B2(n_945),
.Y(n_6629)
);

OAI22x1_ASAP7_75t_L g6630 ( 
.A1(n_6611),
.A2(n_947),
.B1(n_945),
.B2(n_946),
.Y(n_6630)
);

OAI22x1_ASAP7_75t_L g6631 ( 
.A1(n_6611),
.A2(n_949),
.B1(n_947),
.B2(n_948),
.Y(n_6631)
);

CKINVDCx5p33_ASAP7_75t_R g6632 ( 
.A(n_6621),
.Y(n_6632)
);

OAI22xp5_ASAP7_75t_L g6633 ( 
.A1(n_6623),
.A2(n_949),
.B1(n_947),
.B2(n_948),
.Y(n_6633)
);

AOI22xp5_ASAP7_75t_L g6634 ( 
.A1(n_6624),
.A2(n_951),
.B1(n_948),
.B2(n_950),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6628),
.Y(n_6635)
);

AND2x2_ASAP7_75t_L g6636 ( 
.A(n_6626),
.B(n_950),
.Y(n_6636)
);

AOI22xp5_ASAP7_75t_L g6637 ( 
.A1(n_6622),
.A2(n_952),
.B1(n_950),
.B2(n_951),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_6629),
.B(n_952),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6637),
.Y(n_6639)
);

AOI22xp5_ASAP7_75t_L g6640 ( 
.A1(n_6632),
.A2(n_6627),
.B1(n_6625),
.B2(n_6630),
.Y(n_6640)
);

HB1xp67_ASAP7_75t_L g6641 ( 
.A(n_6633),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6634),
.Y(n_6642)
);

OAI222xp33_ASAP7_75t_L g6643 ( 
.A1(n_6640),
.A2(n_6638),
.B1(n_6635),
.B2(n_6636),
.C1(n_6631),
.C2(n_957),
.Y(n_6643)
);

NAND2xp5_ASAP7_75t_L g6644 ( 
.A(n_6641),
.B(n_6639),
.Y(n_6644)
);

OAI22xp5_ASAP7_75t_L g6645 ( 
.A1(n_6642),
.A2(n_953),
.B1(n_954),
.B2(n_955),
.Y(n_6645)
);

NAND2xp5_ASAP7_75t_L g6646 ( 
.A(n_6644),
.B(n_953),
.Y(n_6646)
);

AOI21xp5_ASAP7_75t_L g6647 ( 
.A1(n_6643),
.A2(n_953),
.B(n_954),
.Y(n_6647)
);

AO22x2_ASAP7_75t_L g6648 ( 
.A1(n_6647),
.A2(n_6645),
.B1(n_1083),
.B2(n_1081),
.Y(n_6648)
);

AOI21xp5_ASAP7_75t_L g6649 ( 
.A1(n_6648),
.A2(n_6646),
.B(n_954),
.Y(n_6649)
);

AOI22xp33_ASAP7_75t_L g6650 ( 
.A1(n_6649),
.A2(n_955),
.B1(n_956),
.B2(n_957),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_6650),
.Y(n_6651)
);

AOI211xp5_ASAP7_75t_L g6652 ( 
.A1(n_6651),
.A2(n_956),
.B(n_957),
.C(n_958),
.Y(n_6652)
);


endmodule