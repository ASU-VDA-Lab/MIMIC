module fake_jpeg_24705_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_31),
.Y(n_64)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_63),
.B1(n_38),
.B2(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_64),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_73),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_69),
.B(n_47),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_36),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_44),
.C(n_40),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_37),
.B1(n_45),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_72),
.A2(n_27),
.B1(n_19),
.B2(n_35),
.Y(n_125)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_83),
.B1(n_34),
.B2(n_48),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_23),
.B1(n_20),
.B2(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_43),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_95),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_37),
.B1(n_45),
.B2(n_39),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_91),
.B1(n_61),
.B2(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_39),
.B1(n_34),
.B2(n_20),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_97),
.B1(n_30),
.B2(n_44),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_43),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_115),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_109),
.B1(n_125),
.B2(n_19),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_53),
.B1(n_62),
.B2(n_47),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_53),
.C(n_32),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_74),
.B(n_28),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_42),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_42),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_46),
.B1(n_28),
.B2(n_27),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_31),
.B1(n_25),
.B2(n_41),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_88),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_SL g151 ( 
.A(n_126),
.Y(n_151)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_136),
.Y(n_160)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_134),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_147),
.C(n_77),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_76),
.B1(n_97),
.B2(n_94),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_150),
.Y(n_180)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_144),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_35),
.B1(n_77),
.B2(n_85),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_70),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_71),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_91),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_72),
.B1(n_40),
.B2(n_44),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_127),
.B1(n_113),
.B2(n_21),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_101),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_89),
.B1(n_118),
.B2(n_110),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_181),
.B1(n_179),
.B2(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_137),
.B1(n_25),
.B2(n_21),
.Y(n_211)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_164),
.B(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_129),
.B(n_17),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_17),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_110),
.B1(n_92),
.B2(n_105),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_107),
.B1(n_82),
.B2(n_79),
.Y(n_213)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_174),
.B(n_179),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_44),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_182),
.C(n_184),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_111),
.B(n_101),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_148),
.B(n_140),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_111),
.B1(n_126),
.B2(n_113),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_40),
.C(n_124),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_40),
.C(n_17),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_107),
.C(n_66),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_17),
.C(n_32),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_148),
.B1(n_142),
.B2(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_190),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_191),
.A2(n_198),
.B(n_211),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_199),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_209),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_168),
.B1(n_188),
.B2(n_183),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_128),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_32),
.B(n_17),
.C(n_21),
.D(n_22),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_208),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_144),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_0),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_168),
.B1(n_165),
.B2(n_184),
.Y(n_212)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_33),
.B(n_22),
.C(n_3),
.D(n_4),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_175),
.C(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_216),
.B(n_217),
.Y(n_226)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_218),
.B(n_8),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_171),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_243),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_212),
.B1(n_214),
.B2(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_33),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_33),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_22),
.C(n_2),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_242),
.C(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_11),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_195),
.B1(n_203),
.B2(n_194),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_3),
.C(n_4),
.Y(n_242)
);

NOR4xp25_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_190),
.A2(n_5),
.B(n_7),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_201),
.B(n_200),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_9),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_242),
.C(n_233),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_257),
.B(n_239),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_227),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_235),
.C(n_234),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_198),
.B(n_208),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_223),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_197),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_9),
.C(n_10),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_240),
.C(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_16),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_10),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_239),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_270),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_225),
.C(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

OA21x2_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_230),
.B(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_266),
.B1(n_264),
.B2(n_236),
.Y(n_291)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_283),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_229),
.C(n_222),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_249),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_300),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_286),
.A2(n_254),
.B1(n_266),
.B2(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_295),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_258),
.B1(n_262),
.B2(n_271),
.Y(n_303)
);

BUFx12_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_274),
.C(n_226),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_238),
.B1(n_268),
.B2(n_260),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_279),
.B1(n_280),
.B2(n_275),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_303),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_311),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_313),
.C(n_294),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_13),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_301),
.CI(n_297),
.CON(n_309),
.SN(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_13),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_14),
.C(n_15),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_321),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_309),
.B(n_295),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_303),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_295),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_307),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_310),
.B(n_313),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_328),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_318),
.C2(n_325),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_309),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_315),
.B(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_314),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_332),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_327),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

AOI31xp67_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_330),
.A3(n_327),
.B(n_15),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);


endmodule