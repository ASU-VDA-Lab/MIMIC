module fake_jpeg_23554_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_149;
wire n_35;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_61),
.B1(n_24),
.B2(n_32),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_66),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_19),
.C(n_34),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_49),
.C(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_36),
.Y(n_100)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_28),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_74),
.Y(n_106)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_44),
.B1(n_33),
.B2(n_39),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_75),
.A2(n_104),
.B1(n_63),
.B2(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_78),
.B1(n_83),
.B2(n_103),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_33),
.B1(n_44),
.B2(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_87),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_32),
.B1(n_24),
.B2(n_17),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_93),
.B1(n_48),
.B2(n_41),
.Y(n_107)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_94),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_42),
.B1(n_39),
.B2(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_102),
.Y(n_126)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_41),
.B(n_36),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_42),
.B1(n_32),
.B2(n_24),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_46),
.A2(n_36),
.B(n_26),
.C(n_29),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_130),
.B1(n_48),
.B2(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_121),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_1),
.Y(n_113)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_122),
.Y(n_138)
);

OAI22x1_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_26),
.B1(n_42),
.B2(n_62),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_96),
.B1(n_43),
.B2(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_129),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_68),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_64),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_50),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_71),
.B1(n_94),
.B2(n_89),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_92),
.A2(n_50),
.B1(n_41),
.B2(n_48),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_72),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_55),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_132),
.B(n_31),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_102),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_104),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_119),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_136),
.B(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_147),
.B1(n_158),
.B2(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_162),
.B(n_158),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_129),
.B1(n_109),
.B2(n_123),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_165),
.B(n_111),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_99),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_80),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_101),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_160),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_35),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_63),
.B1(n_43),
.B2(n_76),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_28),
.B(n_27),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_31),
.B(n_19),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_43),
.B1(n_88),
.B2(n_87),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_27),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

AO22x2_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_43),
.B1(n_25),
.B2(n_20),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_150),
.B1(n_118),
.B2(n_22),
.Y(n_213)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_172),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_112),
.C(n_110),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_179),
.C(n_188),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_113),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_190),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_161),
.C(n_135),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_106),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_184),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_165),
.B1(n_145),
.B2(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_111),
.B(n_125),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_116),
.C(n_119),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_22),
.Y(n_216)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_113),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_122),
.C(n_131),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_22),
.C(n_20),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_147),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_136),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_203),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

AOI221xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_159),
.B1(n_165),
.B2(n_143),
.C(n_140),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_209),
.A3(n_212),
.B1(n_35),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_18),
.B1(n_25),
.B2(n_35),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_150),
.B1(n_165),
.B2(n_31),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_213),
.B1(n_214),
.B2(n_169),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_183),
.B1(n_185),
.B2(n_184),
.C(n_194),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_165),
.C(n_17),
.Y(n_210)
);

OAI322xp33_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_180),
.A3(n_192),
.B1(n_189),
.B2(n_178),
.C1(n_171),
.C2(n_166),
.Y(n_221)
);

AOI221xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_20),
.B1(n_18),
.B2(n_35),
.C(n_25),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_17),
.B1(n_19),
.B2(n_34),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_118),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_195),
.C(n_177),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_11),
.C(n_3),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_225),
.C(n_228),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_188),
.B(n_172),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_239),
.B(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_215),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_176),
.C(n_169),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_231),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_197),
.C(n_207),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_168),
.B1(n_2),
.B2(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_219),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_20),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_237),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_2),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_216),
.B(n_205),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_25),
.C(n_35),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_200),
.A2(n_196),
.B1(n_199),
.B2(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_35),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_218),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_232),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_202),
.B1(n_2),
.B2(n_7),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_257),
.B1(n_227),
.B2(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_16),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_234),
.B(n_223),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_264),
.B(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_249),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_233),
.B(n_231),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_226),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_249),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_225),
.C(n_222),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.C(n_2),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_242),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_244),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_273),
.B(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_250),
.B1(n_255),
.B2(n_247),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_265),
.B(n_254),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_277),
.B(n_278),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_276),
.B(n_261),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_245),
.B(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_252),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_281),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_246),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_264),
.B(n_268),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_285),
.B(n_289),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_9),
.C(n_10),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_8),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_289),
.A2(n_269),
.B(n_9),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_291),
.B(n_292),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_10),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_293),
.B(n_13),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_11),
.C(n_13),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_11),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_297),
.B1(n_14),
.B2(n_15),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_294),
.C(n_15),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_301),
.B(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_14),
.Y(n_303)
);


endmodule