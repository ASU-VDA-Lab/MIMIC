module fake_jpeg_4849_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_72),
.B1(n_49),
.B2(n_52),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_48),
.B1(n_61),
.B2(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_59),
.CON(n_70),
.SN(n_70)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_46),
.B1(n_45),
.B2(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_0),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_58),
.B1(n_54),
.B2(n_48),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_61),
.B1(n_65),
.B2(n_64),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_77),
.B1(n_53),
.B2(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_57),
.B1(n_47),
.B2(n_50),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_46),
.B(n_60),
.C(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_73),
.B1(n_78),
.B2(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_75),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_90),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_95),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_75),
.B1(n_5),
.B2(n_7),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_97),
.B(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_94),
.C(n_93),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.C(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_89),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_16),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_18),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_19),
.B(n_21),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_24),
.A3(n_27),
.B1(n_30),
.B2(n_31),
.C1(n_32),
.C2(n_34),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_36),
.B(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_39),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_41),
.Y(n_111)
);


endmodule