module fake_jpeg_17112_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_50),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_54),
.B1(n_51),
.B2(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_53),
.B1(n_56),
.B2(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_53),
.B1(n_56),
.B2(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_55),
.B1(n_47),
.B2(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_63),
.B(n_1),
.C(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_108),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_4),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_104),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_6),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_19),
.Y(n_115)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_120),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_91),
.C(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_119),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_123),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_96),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_119),
.C(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_141),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_93),
.B(n_110),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_140),
.C(n_139),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_147),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_144),
.C(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_27),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_30),
.B(n_33),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_34),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_127),
.B(n_36),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_156),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_35),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_37),
.CI(n_38),
.CON(n_159),
.SN(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_127),
.Y(n_160)
);


endmodule