module fake_jpeg_1110_n_681 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_681);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_681;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g176 ( 
.A(n_60),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_61),
.A2(n_56),
.B1(n_53),
.B2(n_50),
.Y(n_177)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_10),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_64),
.B(n_76),
.Y(n_146)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_67),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_46),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_77),
.B(n_79),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_78),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_19),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_80),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_117),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_92),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_34),
.B(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_93),
.B(n_96),
.Y(n_210)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_18),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_98),
.B(n_55),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_108),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_18),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_17),
.Y(n_161)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

CKINVDCx6p67_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_22),
.B(n_17),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g207 ( 
.A(n_121),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_124),
.B(n_127),
.Y(n_200)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_56),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_26),
.B1(n_32),
.B2(n_22),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_139),
.A2(n_224),
.B1(n_108),
.B2(n_88),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_67),
.A2(n_52),
.B1(n_32),
.B2(n_45),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_143),
.A2(n_147),
.B1(n_149),
.B2(n_153),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_63),
.A2(n_26),
.B1(n_32),
.B2(n_45),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_26),
.B1(n_45),
.B2(n_49),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_49),
.B1(n_55),
.B2(n_50),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_161),
.B(n_203),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_165),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_49),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_171),
.B(n_172),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_55),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_177),
.A2(n_226),
.B1(n_99),
.B2(n_97),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_178),
.B(n_187),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_68),
.A2(n_50),
.B1(n_42),
.B2(n_56),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_180),
.A2(n_194),
.B1(n_195),
.B2(n_206),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_24),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_24),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_189),
.B(n_193),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_24),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_122),
.A2(n_42),
.B1(n_53),
.B2(n_57),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_42),
.B1(n_53),
.B2(n_57),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_60),
.B(n_40),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_198),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_40),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_73),
.B(n_40),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_204),
.B(n_214),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_70),
.A2(n_58),
.B1(n_57),
.B2(n_51),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_94),
.A2(n_39),
.B1(n_58),
.B2(n_51),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_211),
.B1(n_125),
.B2(n_126),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_78),
.A2(n_39),
.B1(n_58),
.B2(n_51),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_130),
.A2(n_39),
.B(n_29),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_213),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_65),
.B(n_29),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_104),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_215),
.B(n_216),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_124),
.B(n_59),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_131),
.A2(n_59),
.B1(n_23),
.B2(n_21),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_85),
.A2(n_59),
.B(n_23),
.C(n_21),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_225),
.B(n_1),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_72),
.A2(n_115),
.B1(n_111),
.B2(n_80),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_228),
.Y(n_326)
);

NAND2xp67_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_198),
.Y(n_229)
);

NAND2xp67_ASAP7_75t_L g339 ( 
.A(n_229),
.B(n_241),
.Y(n_339)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_230),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_231),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_23),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_232),
.B(n_243),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_233),
.A2(n_240),
.B1(n_154),
.B2(n_159),
.Y(n_366)
);

INVx4_ASAP7_75t_SL g234 ( 
.A(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_234),
.Y(n_356)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_235),
.Y(n_334)
);

OA22x2_ASAP7_75t_L g357 ( 
.A1(n_237),
.A2(n_222),
.B1(n_202),
.B2(n_218),
.Y(n_357)
);

AO22x1_ASAP7_75t_SL g238 ( 
.A1(n_135),
.A2(n_83),
.B1(n_81),
.B2(n_86),
.Y(n_238)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_238),
.Y(n_341)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_0),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_90),
.B1(n_100),
.B2(n_103),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_242),
.A2(n_292),
.B1(n_154),
.B2(n_218),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_140),
.B(n_0),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_176),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_146),
.B(n_0),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_261),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_247),
.B(n_279),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_174),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_248),
.B(n_249),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_174),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_251),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_132),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_253),
.B(n_255),
.Y(n_331)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_150),
.Y(n_254)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_158),
.Y(n_259)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_260),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_1),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_262),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_176),
.A2(n_82),
.B1(n_74),
.B2(n_69),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_263),
.A2(n_264),
.B1(n_276),
.B2(n_300),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_148),
.A2(n_66),
.B1(n_48),
.B2(n_12),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_173),
.Y(n_265)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_167),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_1),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_287),
.Y(n_310)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_213),
.A2(n_48),
.B1(n_17),
.B2(n_16),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_270),
.A2(n_305),
.B1(n_170),
.B2(n_164),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_273),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_160),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_212),
.B(n_1),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_283),
.B(n_182),
.Y(n_322)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_169),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_155),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_281),
.B(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_184),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_282),
.B(n_285),
.Y(n_350)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_168),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_143),
.B(n_1),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_155),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_134),
.B(n_48),
.C(n_16),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_271),
.C(n_246),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_157),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_291),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_137),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_294),
.Y(n_365)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_197),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_163),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_296),
.Y(n_361)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_209),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_162),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_298),
.Y(n_362)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_163),
.Y(n_298)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_133),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_205),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_301),
.B(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_306),
.B1(n_220),
.B2(n_144),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_183),
.A2(n_185),
.B1(n_170),
.B2(n_142),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_133),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_149),
.B(n_2),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_2),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_309),
.B(n_325),
.Y(n_410)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_229),
.A2(n_200),
.B(n_208),
.C(n_211),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_315),
.A2(n_241),
.B(n_278),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_256),
.A2(n_144),
.B1(n_160),
.B2(n_182),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_320),
.A2(n_323),
.B1(n_337),
.B2(n_357),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_321),
.B(n_332),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_322),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_257),
.A2(n_188),
.B1(n_192),
.B2(n_166),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_221),
.C(n_201),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_261),
.B(n_183),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_344),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_232),
.B(n_304),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_202),
.C(n_222),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_245),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_260),
.A2(n_192),
.B1(n_166),
.B2(n_220),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_268),
.B(n_185),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_233),
.A2(n_145),
.B1(n_152),
.B2(n_142),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_345),
.A2(n_351),
.B1(n_358),
.B2(n_366),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_349),
.A2(n_228),
.B1(n_276),
.B2(n_300),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_242),
.A2(n_145),
.B1(n_152),
.B2(n_164),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_290),
.B(n_162),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_359),
.B(n_306),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_283),
.B(n_2),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_364),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_283),
.B(n_3),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_277),
.A2(n_138),
.B1(n_4),
.B2(n_5),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_287),
.B1(n_234),
.B2(n_307),
.Y(n_388)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_354),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_375),
.Y(n_449)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_378),
.Y(n_429)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_383),
.Y(n_459)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_386),
.Y(n_431)
);

AOI211xp5_ASAP7_75t_L g387 ( 
.A1(n_310),
.A2(n_339),
.B(n_321),
.C(n_364),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_387),
.B(n_404),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_388),
.A2(n_394),
.B1(n_397),
.B2(n_408),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_341),
.A2(n_299),
.B1(n_252),
.B2(n_236),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_389),
.A2(n_393),
.B1(n_399),
.B2(n_417),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_395),
.Y(n_451)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_310),
.B(n_275),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_405),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_341),
.A2(n_238),
.B1(n_266),
.B2(n_243),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_396),
.A2(n_415),
.B(n_312),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_358),
.A2(n_238),
.B1(n_292),
.B2(n_276),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_311),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_398),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_366),
.A2(n_297),
.B1(n_279),
.B2(n_285),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_362),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_401),
.Y(n_450)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_336),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_402),
.Y(n_442)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_403),
.B(n_406),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_350),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_308),
.B(n_289),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_365),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_365),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_407),
.B(n_409),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_347),
.A2(n_250),
.B1(n_235),
.B2(n_262),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

AOI22x1_ASAP7_75t_L g411 ( 
.A1(n_322),
.A2(n_315),
.B1(n_368),
.B2(n_339),
.Y(n_411)
);

AO22x1_ASAP7_75t_SL g447 ( 
.A1(n_411),
.A2(n_357),
.B1(n_351),
.B2(n_345),
.Y(n_447)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_414),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_347),
.A2(n_267),
.B1(n_254),
.B2(n_273),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_413),
.A2(n_353),
.B1(n_355),
.B2(n_356),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_327),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_327),
.A2(n_230),
.B1(n_251),
.B2(n_286),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_317),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_353),
.A2(n_296),
.B1(n_294),
.B2(n_239),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_SL g418 ( 
.A(n_308),
.B(n_302),
.C(n_301),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_418),
.B(n_363),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_333),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_420),
.B(n_423),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_404),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_424),
.C(n_438),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_333),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_309),
.C(n_335),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_425),
.B(n_453),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_372),
.A2(n_346),
.B(n_331),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_435),
.A2(n_439),
.B(n_457),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_381),
.B(n_325),
.Y(n_438)
);

XNOR2x1_ASAP7_75t_L g441 ( 
.A(n_372),
.B(n_344),
.Y(n_441)
);

XOR2x1_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_396),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_392),
.B(n_328),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_444),
.C(n_377),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_359),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_452),
.Y(n_468)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_448),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_380),
.B(n_350),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_398),
.B(n_361),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_386),
.B(n_356),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_373),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_411),
.A2(n_327),
.B(n_319),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_458),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_428),
.A2(n_389),
.B1(n_371),
.B2(n_397),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_463),
.A2(n_478),
.B1(n_482),
.B2(n_495),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_401),
.C(n_406),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_435),
.Y(n_505)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_433),
.Y(n_465)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_456),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_466),
.B(n_496),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_467),
.B(n_471),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_371),
.B1(n_407),
.B2(n_411),
.Y(n_469)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_469),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_391),
.C(n_382),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_472),
.C(n_489),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_382),
.C(n_387),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_376),
.Y(n_473)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_473),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_440),
.Y(n_474)
);

INVx13_ASAP7_75t_L g534 ( 
.A(n_474),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_475),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_428),
.A2(n_388),
.B1(n_385),
.B2(n_403),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_477),
.A2(n_431),
.B1(n_447),
.B2(n_444),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_457),
.A2(n_393),
.B1(n_399),
.B2(n_416),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_479),
.B(n_481),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_432),
.A2(n_412),
.B1(n_374),
.B2(n_414),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_483),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_438),
.B(n_370),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_486),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_426),
.B(n_375),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_485),
.B(n_488),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_418),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_446),
.A2(n_413),
.B1(n_408),
.B2(n_379),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_490),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_426),
.B(n_409),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_227),
.C(n_280),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_384),
.Y(n_490)
);

OAI32xp33_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_318),
.A3(n_348),
.B1(n_367),
.B2(n_330),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_434),
.B(n_449),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_400),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_442),
.Y(n_501)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_427),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_493),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_439),
.A2(n_357),
.B(n_317),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_494),
.A2(n_480),
.B(n_478),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_431),
.A2(n_357),
.B1(n_355),
.B2(n_378),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_443),
.B(n_369),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_427),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_497),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_500),
.A2(n_505),
.B1(n_509),
.B2(n_512),
.Y(n_564)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_501),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_451),
.Y(n_506)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_506),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_434),
.Y(n_507)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_459),
.Y(n_510)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_477),
.A2(n_463),
.B1(n_462),
.B2(n_468),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_468),
.A2(n_447),
.B1(n_442),
.B2(n_441),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_513),
.A2(n_531),
.B1(n_519),
.B2(n_502),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_480),
.A2(n_430),
.B(n_422),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_462),
.A2(n_448),
.B1(n_430),
.B2(n_422),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_515),
.A2(n_522),
.B1(n_532),
.B2(n_497),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_484),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_461),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_527),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_518),
.A2(n_402),
.B(n_314),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_454),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_520),
.B(n_521),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_460),
.B(n_318),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_465),
.A2(n_436),
.B1(n_437),
.B2(n_429),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_476),
.B(n_338),
.Y(n_524)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_524),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_475),
.B(n_419),
.Y(n_525)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_525),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_481),
.B(n_436),
.C(n_419),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_489),
.C(n_471),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_492),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_483),
.A2(n_437),
.B1(n_429),
.B2(n_378),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_535),
.B(n_562),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_536),
.A2(n_538),
.B1(n_541),
.B2(n_498),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_537),
.B(n_560),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_495),
.B1(n_482),
.B2(n_479),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_519),
.A2(n_491),
.B1(n_494),
.B2(n_486),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_543),
.B(n_565),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_545),
.A2(n_554),
.B1(n_567),
.B2(n_530),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_507),
.B(n_490),
.Y(n_548)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_520),
.C(n_504),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_552),
.C(n_557),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_504),
.B(n_470),
.C(n_472),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_525),
.Y(n_553)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_553),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_512),
.A2(n_493),
.B1(n_352),
.B2(n_313),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_508),
.B(n_338),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_556),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_526),
.B(n_334),
.C(n_369),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_558),
.A2(n_563),
.B(n_533),
.Y(n_586)
);

FAx1_ASAP7_75t_SL g559 ( 
.A(n_513),
.B(n_336),
.CI(n_402),
.CON(n_559),
.SN(n_559)
);

FAx1_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_258),
.CI(n_303),
.CON(n_587),
.SN(n_587)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_499),
.B(n_367),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_501),
.Y(n_561)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_561),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_516),
.B(n_348),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_518),
.A2(n_334),
.B(n_383),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_534),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_511),
.B(n_499),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_511),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_509),
.A2(n_352),
.B1(n_313),
.B2(n_383),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g568 ( 
.A1(n_537),
.A2(n_529),
.B(n_500),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g611 ( 
.A(n_568),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_582),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_542),
.A2(n_514),
.B(n_528),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_574),
.A2(n_576),
.B1(n_563),
.B2(n_540),
.Y(n_603)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_575),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_542),
.A2(n_528),
.B(n_503),
.Y(n_576)
);

OAI22x1_ASAP7_75t_L g579 ( 
.A1(n_541),
.A2(n_515),
.B1(n_531),
.B2(n_498),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_579),
.A2(n_580),
.B1(n_585),
.B2(n_591),
.Y(n_600)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_581),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_522),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_549),
.B(n_532),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_583),
.B(n_590),
.Y(n_606)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_548),
.Y(n_584)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_584),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_538),
.A2(n_533),
.B1(n_530),
.B2(n_534),
.Y(n_585)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_586),
.Y(n_605)
);

AOI211xp5_ASAP7_75t_L g612 ( 
.A1(n_587),
.A2(n_567),
.B(n_545),
.C(n_554),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_549),
.B(n_330),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_536),
.A2(n_291),
.B1(n_272),
.B2(n_244),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_535),
.B(n_269),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_593),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_265),
.Y(n_593)
);

INVx11_ASAP7_75t_L g595 ( 
.A(n_587),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g620 ( 
.A1(n_595),
.A2(n_603),
.B1(n_609),
.B2(n_610),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_571),
.B(n_552),
.C(n_557),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_597),
.B(n_599),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_571),
.B(n_560),
.C(n_546),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_561),
.Y(n_602)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_602),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_593),
.B(n_564),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_583),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_562),
.C(n_558),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_569),
.C(n_590),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_578),
.A2(n_550),
.B1(n_555),
.B2(n_559),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_587),
.A2(n_555),
.B1(n_559),
.B2(n_543),
.Y(n_610)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_612),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_580),
.A2(n_544),
.B1(n_547),
.B2(n_231),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_613),
.A2(n_575),
.B1(n_577),
.B2(n_572),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_570),
.B(n_259),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_3),
.Y(n_632)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_576),
.Y(n_615)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_615),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_616),
.A2(n_626),
.B1(n_629),
.B2(n_630),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_619),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_602),
.B(n_585),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_621),
.B(n_622),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_582),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_623),
.B(n_634),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_597),
.B(n_588),
.C(n_573),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_631),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_SL g626 ( 
.A1(n_605),
.A2(n_579),
.B(n_574),
.C(n_586),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_605),
.A2(n_569),
.B(n_591),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_627),
.A2(n_607),
.B(n_608),
.Y(n_646)
);

OAI321xp33_ASAP7_75t_L g629 ( 
.A1(n_596),
.A2(n_592),
.A3(n_16),
.B1(n_14),
.B2(n_13),
.C(n_3),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_600),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_615),
.B(n_3),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_632),
.B(n_633),
.Y(n_642)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_609),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_612),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_618),
.B(n_598),
.C(n_604),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_639),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_628),
.A2(n_611),
.B1(n_598),
.B2(n_610),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_638),
.Y(n_656)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_617),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_620),
.A2(n_624),
.B(n_633),
.Y(n_640)
);

AOI21xp33_ASAP7_75t_L g653 ( 
.A1(n_640),
.A2(n_621),
.B(n_624),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_616),
.A2(n_613),
.B1(n_600),
.B2(n_594),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_643),
.B(n_647),
.Y(n_658)
);

XNOR2x1_ASAP7_75t_SL g644 ( 
.A(n_627),
.B(n_604),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_644),
.A2(n_637),
.B(n_638),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_646),
.A2(n_606),
.B(n_626),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_622),
.B(n_601),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_625),
.B(n_606),
.C(n_601),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_649),
.B(n_595),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_651),
.Y(n_663)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_646),
.B(n_619),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_653),
.A2(n_639),
.B(n_648),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_654),
.B(n_655),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_623),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_636),
.B(n_630),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_657),
.B(n_659),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_641),
.B(n_631),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_660),
.Y(n_662)
);

AOI21x1_ASAP7_75t_L g669 ( 
.A1(n_665),
.A2(n_656),
.B(n_649),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_652),
.B(n_645),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_SL g670 ( 
.A1(n_666),
.A2(n_656),
.B(n_635),
.C(n_644),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_658),
.A2(n_635),
.B(n_642),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_667),
.B(n_668),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_651),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_669),
.A2(n_662),
.B(n_661),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_670),
.B(n_663),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_664),
.B(n_643),
.C(n_6),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_673),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_666),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_674),
.A2(n_675),
.B(n_4),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_671),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_677),
.A2(n_678),
.B(n_6),
.C(n_7),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_6),
.Y(n_680)
);

FAx1_ASAP7_75t_SL g681 ( 
.A(n_680),
.B(n_7),
.CI(n_678),
.CON(n_681),
.SN(n_681)
);


endmodule