module real_jpeg_6904_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_128),
.B1(n_129),
.B2(n_134),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_1),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_128),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_1),
.A2(n_128),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_3),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_3),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_3),
.A2(n_143),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_4),
.A2(n_50),
.B1(n_177),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_4),
.A2(n_50),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_4),
.A2(n_50),
.B1(n_280),
.B2(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_5),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_5),
.A2(n_63),
.B1(n_161),
.B2(n_271),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_5),
.A2(n_63),
.B1(n_92),
.B2(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_6),
.A2(n_190),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_6),
.B(n_167),
.C(n_251),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_6),
.A2(n_157),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_6),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_6),
.A2(n_85),
.B1(n_300),
.B2(n_303),
.Y(n_307)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_8),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_9),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_9),
.A2(n_93),
.B1(n_218),
.B2(n_221),
.Y(n_217)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_12),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_13),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_14),
.Y(n_119)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_14),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_15),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_243),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_241),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_171),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_19),
.B(n_171),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.C(n_146),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_20),
.A2(n_21),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_67),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_22),
.B(n_68),
.C(n_105),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_48),
.B2(n_57),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_23),
.A2(n_25),
.B1(n_57),
.B2(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_24),
.A2(n_49),
.B1(n_268),
.B2(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_25),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_28),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_28),
.Y(n_220)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_29),
.Y(n_136)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_29),
.Y(n_162)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_29),
.Y(n_222)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_30),
.Y(n_155)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_32),
.Y(n_160)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_33),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_40),
.Y(n_185)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_40),
.Y(n_211)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_46),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_52),
.Y(n_321)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_56),
.Y(n_176)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_64),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_97),
.B2(n_105),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_79),
.B(n_84),
.Y(n_69)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_72),
.Y(n_302)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_78),
.Y(n_290)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_80),
.B(n_157),
.Y(n_309)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_85),
.A2(n_164),
.B(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_85),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_85),
.A2(n_274),
.B(n_281),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_85),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_85),
.A2(n_289),
.B1(n_300),
.B2(n_303),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_90),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_95),
.B(n_309),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_99),
.A2(n_224),
.B1(n_227),
.B2(n_236),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_100),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_106),
.A2(n_146),
.B1(n_147),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_106),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_126),
.B(n_137),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_107),
.A2(n_140),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_108),
.A2(n_216),
.B1(n_254),
.B2(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_108),
.A2(n_216),
.B1(n_258),
.B2(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_108),
.A2(n_127),
.B1(n_216),
.B2(n_270),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_109)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_110),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_116),
.Y(n_263)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_117),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_118)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_123),
.Y(n_276)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_123),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_125),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_136),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_139),
.B(n_157),
.Y(n_298)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_163),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_148),
.B(n_163),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.A3(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g319 ( 
.A1(n_156),
.A2(n_157),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_164),
.Y(n_282)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_205),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_204),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_194),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_177),
.A3(n_180),
.B1(n_184),
.B2(n_189),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx6_ASAP7_75t_SL g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_197),
.Y(n_284)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_205),
.Y(n_331)
);

FAx1_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_214),
.CI(n_223),
.CON(n_205),
.SN(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_234),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_324),
.B(n_330),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_313),
.B(n_323),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_285),
.B(n_312),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_264),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_264),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_253),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_272),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_272),
.C(n_273),
.Y(n_314)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_269),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_296),
.B(n_311),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_295),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_295),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_306),
.B(n_310),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_315),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_318),
.C(n_322),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_322),
.Y(n_317)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule