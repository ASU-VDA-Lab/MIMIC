module real_jpeg_19114_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_286;
wire n_288;
wire n_292;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx13_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_151),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_151),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_3),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_116),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_116),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_116),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_4),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_4),
.B(n_24),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_12),
.B(n_49),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_81),
.B1(n_83),
.B2(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_27),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_4),
.A2(n_27),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_48),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_53),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_25),
.B1(n_27),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_8),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_145),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_145),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_145),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_32),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_11),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_12),
.A2(n_43),
.B(n_46),
.C(n_47),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_12),
.B(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_35),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_14),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_14),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_107)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_95),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_19),
.B(n_95),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_19),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_68),
.CI(n_77),
.CON(n_19),
.SN(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_33),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_23),
.A2(n_91),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_23),
.A2(n_91),
.B1(n_115),
.B2(n_162),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_24),
.B(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_24),
.A2(n_36),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_25),
.A2(n_37),
.B1(n_148),
.B2(n_155),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_25),
.A2(n_43),
.A3(n_62),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_26),
.B(n_27),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_30),
.B(n_149),
.CON(n_148),
.SN(n_148)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_51),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_42),
.A2(n_47),
.B1(n_87),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_42),
.A2(n_51),
.B(n_88),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_42),
.A2(n_47),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_42),
.A2(n_47),
.B1(n_205),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_42),
.A2(n_47),
.B1(n_225),
.B2(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_42),
.A2(n_72),
.B(n_241),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_44),
.A2(n_50),
.B(n_149),
.C(n_201),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_44),
.B(n_58),
.Y(n_235)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_47),
.A2(n_74),
.B(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_47),
.B(n_149),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_48),
.B(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_66),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_56),
.B(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_56),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_56),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_56),
.A2(n_66),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_57),
.A2(n_61),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_57),
.A2(n_61),
.B1(n_182),
.B2(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_70),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_61),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_67),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_90),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_79),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_80),
.A2(n_86),
.B1(n_89),
.B2(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B(n_84),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_81),
.A2(n_83),
.B1(n_134),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_81),
.A2(n_110),
.B1(n_194),
.B2(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_81),
.A2(n_108),
.B(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_82),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_82),
.A2(n_85),
.B(n_136),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_107),
.Y(n_136)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_83),
.B(n_149),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_86),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_94),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_115),
.B(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_101),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_96),
.B(n_100),
.Y(n_301)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_101),
.A2(n_102),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.C(n_118),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_103),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_104),
.B(n_111),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

OAI21x1_ASAP7_75t_SL g177 ( 
.A1(n_105),
.A2(n_157),
.B(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_297),
.B(n_302),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_285),
.B(n_296),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_185),
.B(n_264),
.C(n_284),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_169),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_128),
.B(n_169),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_152),
.B2(n_168),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_139),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_131),
.B(n_139),
.C(n_168),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_132),
.B(n_138),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_147),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_153),
.B(n_159),
.C(n_164),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_167),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_180),
.B(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_263),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_258),
.B(n_262),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_246),
.B(n_257),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_228),
.B(n_245),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_217),
.B(n_227),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_206),
.B(n_216),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_202),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_211),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_231),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_237),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_255),
.C(n_256),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_282),
.B2(n_283),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_272),
.C(n_283),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_281),
.Y(n_272)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_293),
.C(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);


endmodule