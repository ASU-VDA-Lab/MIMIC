module fake_aes_4759_n_542 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_542);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_542;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_70), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_59), .Y(n_79) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_62), .B(n_58), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_33), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_69), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_64), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_9), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_38), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_60), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_28), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_32), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_54), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_16), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_66), .Y(n_92) );
OR2x2_ASAP7_75t_L g93 ( .A(n_16), .B(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_30), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_48), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_37), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_1), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_24), .Y(n_100) );
BUFx10_ASAP7_75t_L g101 ( .A(n_31), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_14), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_9), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_46), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_71), .Y(n_106) );
BUFx5_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_3), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_1), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_44), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_107), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_110), .B(n_0), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_96), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_97), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_102), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_97), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_110), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_78), .B(n_2), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_96), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_84), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_85), .B(n_4), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_102), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_103), .B(n_5), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_103), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_108), .B(n_6), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_107), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_115), .B(n_98), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_122), .B(n_128), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_131), .B(n_83), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_131), .B(n_101), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_122), .B(n_128), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_133), .B(n_100), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_115), .B(n_93), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_133), .B(n_106), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_115), .A2(n_95), .B1(n_91), .B2(n_90), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_130), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_129), .B(n_101), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
AO21x1_ASAP7_75t_L g151 ( .A1(n_121), .A2(n_79), .B(n_105), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_120), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_120), .B(n_109), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_117), .B(n_112), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_132), .B(n_111), .Y(n_156) );
AO22x2_ASAP7_75t_L g157 ( .A1(n_124), .A2(n_113), .B1(n_92), .B2(n_107), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_125), .B(n_101), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_132), .B(n_107), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_132), .B(n_117), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_119), .B(n_107), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_143), .B(n_125), .Y(n_163) );
INVxp67_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_141), .B(n_127), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_147), .B(n_141), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_157), .A2(n_118), .B1(n_113), .B2(n_126), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_141), .B(n_158), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_158), .B(n_134), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
AOI221xp5_ASAP7_75t_L g173 ( .A1(n_157), .A2(n_119), .B1(n_99), .B2(n_92), .C(n_130), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_151), .A2(n_136), .B1(n_135), .B2(n_123), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_151), .A2(n_136), .B1(n_135), .B2(n_104), .Y(n_175) );
AND3x1_ASAP7_75t_L g176 ( .A(n_149), .B(n_80), .C(n_81), .Y(n_176) );
NOR2xp33_ASAP7_75t_SL g177 ( .A(n_138), .B(n_104), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_138), .A2(n_89), .B1(n_81), .B2(n_123), .Y(n_179) );
NAND2xp33_ASAP7_75t_L g180 ( .A(n_138), .B(n_89), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_139), .B(n_88), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_140), .B(n_123), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_149), .B(n_123), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_138), .A2(n_123), .B1(n_116), .B2(n_10), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_149), .B(n_7), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_139), .B(n_116), .Y(n_188) );
NOR2x2_ASAP7_75t_L g189 ( .A(n_157), .B(n_8), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_142), .B(n_116), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_138), .A2(n_116), .B1(n_10), .B2(n_11), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_144), .B(n_8), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_144), .B(n_43), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_169), .A2(n_144), .B1(n_164), .B2(n_184), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_168), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_167), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_167), .A2(n_157), .B1(n_144), .B2(n_153), .Y(n_199) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_174), .A2(n_159), .B(n_156), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_171), .B(n_138), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_165), .B(n_138), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_187), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_189), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_177), .B(n_153), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_163), .B(n_138), .Y(n_209) );
NAND3xp33_ASAP7_75t_SL g210 ( .A(n_173), .B(n_162), .C(n_145), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_185), .A2(n_137), .B(n_146), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_181), .B(n_153), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_166), .A2(n_162), .B(n_156), .C(n_154), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_191), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_168), .B(n_153), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_178), .B(n_152), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_191), .A2(n_183), .B(n_178), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_175), .A2(n_157), .B1(n_148), .B2(n_146), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_195), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_188), .A2(n_148), .B(n_137), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_193), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_180), .A2(n_159), .B(n_155), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_170), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_179), .B(n_176), .Y(n_226) );
NOR3xp33_ASAP7_75t_SL g227 ( .A(n_182), .B(n_11), .C(n_12), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_176), .A2(n_160), .B1(n_155), .B2(n_15), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_223), .A2(n_186), .B(n_194), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_218), .A2(n_177), .B(n_192), .C(n_155), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_209), .A2(n_194), .B(n_172), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
CKINVDCx6p67_ASAP7_75t_R g233 ( .A(n_204), .Y(n_233) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_227), .B(n_179), .C(n_160), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_210), .A2(n_155), .B(n_160), .C(n_170), .Y(n_235) );
INVxp67_ASAP7_75t_L g236 ( .A(n_208), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_208), .B(n_13), .Y(n_238) );
INVx3_ASAP7_75t_SL g239 ( .A(n_198), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_206), .B(n_13), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_215), .B(n_14), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_225), .B(n_194), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_225), .B(n_17), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_196), .A2(n_172), .B1(n_170), .B2(n_17), .Y(n_245) );
AO31x2_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_172), .A3(n_20), .B(n_21), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_206), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_207), .A2(n_19), .B(n_22), .C(n_23), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_212), .B(n_25), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_202), .B(n_26), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_221), .B(n_27), .Y(n_252) );
AO32x2_ASAP7_75t_L g253 ( .A1(n_199), .A2(n_29), .A3(n_34), .B1(n_35), .B2(n_36), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_205), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_247), .B(n_198), .Y(n_257) );
INVx4_ASAP7_75t_SL g258 ( .A(n_254), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_231), .A2(n_217), .B(n_213), .Y(n_259) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_228), .B(n_211), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_229), .A2(n_220), .B(n_224), .Y(n_262) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_244), .A2(n_201), .B(n_219), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_214), .B(n_203), .C(n_219), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_237), .B(n_226), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_255), .A2(n_219), .B(n_200), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_255), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_243), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_250), .A2(n_219), .B(n_200), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_233), .B(n_226), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_226), .B1(n_214), .B2(n_203), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_219), .B(n_200), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_235), .A2(n_200), .B(n_214), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_242), .A2(n_205), .B(n_42), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_234), .A2(n_205), .B(n_45), .Y(n_277) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_275), .A2(n_245), .B(n_249), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_268), .B(n_238), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_265), .A2(n_240), .B1(n_248), .B2(n_239), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_267), .B(n_253), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_267), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_266), .A2(n_241), .B(n_252), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_268), .B(n_253), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_269), .B(n_251), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_257), .A2(n_239), .B1(n_249), .B2(n_251), .C(n_205), .Y(n_289) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_264), .A2(n_246), .B(n_253), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_256), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_269), .B(n_254), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_262), .Y(n_296) );
INVxp33_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_272), .B(n_253), .Y(n_298) );
AOI21xp5_ASAP7_75t_SL g299 ( .A1(n_272), .A2(n_254), .B(n_253), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_287), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_285), .B(n_260), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_263), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_285), .B(n_260), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_292), .Y(n_305) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_297), .A2(n_283), .B1(n_279), .B2(n_288), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_293), .B(n_263), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_291), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_299), .B(n_273), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_291), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_295), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_285), .B(n_298), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_298), .B(n_260), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_260), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_281), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_281), .B(n_263), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_322), .B(n_281), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_290), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_322), .B(n_290), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_305), .Y(n_333) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_309), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_303), .B(n_294), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_318), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_325), .B(n_290), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_325), .B(n_290), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_306), .B(n_279), .Y(n_340) );
INVx6_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_302), .B(n_280), .C(n_289), .D(n_279), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_325), .B(n_284), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_323), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_303), .B(n_294), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_326), .B(n_284), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_326), .B(n_284), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_306), .B(n_297), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_310), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_302), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_307), .B(n_288), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_307), .B(n_233), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_303), .B(n_284), .Y(n_357) );
NOR4xp25_ASAP7_75t_SL g358 ( .A(n_310), .B(n_289), .C(n_246), .D(n_280), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_326), .B(n_284), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_301), .B(n_278), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_328), .B(n_258), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_312), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_301), .B(n_278), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_301), .B(n_278), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_309), .B(n_261), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_308), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_304), .B(n_278), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_304), .B(n_246), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_304), .B(n_246), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_246), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_329), .B(n_270), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_313), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_366), .B(n_329), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_366), .B(n_328), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_330), .B(n_328), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_344), .B(n_316), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_330), .B(n_313), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_331), .B(n_317), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_340), .B(n_308), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_353), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_335), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_316), .B1(n_305), .B2(n_320), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_362), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_333), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_340), .B(n_321), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_355), .B(n_315), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_335), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_351), .B(n_324), .C(n_311), .D(n_320), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_331), .B(n_321), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_332), .B(n_315), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_335), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_342), .A2(n_316), .B1(n_320), .B2(n_311), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_344), .B(n_316), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_332), .B(n_315), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_372), .B(n_317), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_372), .B(n_317), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_337), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_348), .B(n_327), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_336), .B(n_324), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_343), .B(n_327), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_343), .B(n_327), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_348), .B(n_327), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_345), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_336), .B(n_319), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_346), .B(n_319), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_349), .B(n_319), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_345), .B(n_314), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_347), .B(n_314), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_314), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_342), .A2(n_316), .B1(n_300), .B2(n_276), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_359), .B(n_316), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_347), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_367), .B(n_259), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_346), .B(n_274), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_359), .B(n_274), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_367), .B(n_277), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_338), .B(n_277), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_354), .B(n_41), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_378), .B(n_373), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_380), .B(n_339), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_388), .B(n_339), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_376), .B(n_334), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_374), .B(n_338), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_377), .B(n_333), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
NAND2xp33_ASAP7_75t_SL g438 ( .A(n_389), .B(n_377), .Y(n_438) );
OR2x6_ASAP7_75t_L g439 ( .A(n_399), .B(n_341), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_401), .B(n_352), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_401), .B(n_360), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_392), .B(n_354), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_402), .B(n_360), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_382), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_406), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_384), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_402), .B(n_364), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_379), .B(n_364), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_379), .B(n_365), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_393), .B(n_334), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_384), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_394), .B(n_368), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_394), .B(n_368), .Y(n_454) );
NOR4xp25_ASAP7_75t_L g455 ( .A(n_398), .B(n_417), .C(n_420), .D(n_385), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_400), .B(n_365), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_357), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_400), .B(n_371), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_386), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_375), .B(n_371), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_386), .Y(n_461) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_383), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_413), .B(n_370), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_391), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_391), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_383), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_406), .Y(n_468) );
OAI32xp33_ASAP7_75t_L g469 ( .A1(n_411), .A2(n_357), .A3(n_350), .B1(n_370), .B2(n_369), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_399), .B(n_350), .Y(n_470) );
OAI21xp33_ASAP7_75t_L g471 ( .A1(n_455), .A2(n_418), .B(n_399), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_443), .B(n_416), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_465), .Y(n_473) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_428), .B(n_418), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_468), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_469), .A2(n_418), .B1(n_403), .B2(n_404), .C(n_419), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_456), .B(n_428), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_465), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_443), .A2(n_409), .B(n_416), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_438), .A2(n_407), .B(n_408), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_457), .B(n_463), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_442), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_427), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_430), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_446), .B(n_411), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_433), .Y(n_487) );
AOI21xp33_ASAP7_75t_L g488 ( .A1(n_442), .A2(n_425), .B(n_395), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_438), .B(n_409), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_434), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_436), .A2(n_410), .B(n_423), .C(n_415), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_439), .A2(n_341), .B1(n_412), .B2(n_358), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_436), .A2(n_414), .B(n_358), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_431), .B(n_410), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_432), .B(n_422), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_435), .B(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_439), .A2(n_341), .B1(n_412), .B2(n_350), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_470), .A2(n_421), .B(n_390), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_472), .B(n_440), .Y(n_501) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_471), .A2(n_470), .B(n_451), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g503 ( .A1(n_489), .A2(n_479), .A3(n_492), .B(n_499), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_476), .B(n_462), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_483), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_484), .Y(n_506) );
OAI21xp33_ASAP7_75t_SL g507 ( .A1(n_474), .A2(n_439), .B(n_462), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_492), .A2(n_448), .B(n_444), .C(n_441), .Y(n_508) );
AOI222xp33_ASAP7_75t_L g509 ( .A1(n_480), .A2(n_458), .B1(n_454), .B2(n_453), .C1(n_449), .C2(n_450), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_475), .A2(n_429), .B1(n_437), .B2(n_460), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_487), .A2(n_341), .B1(n_466), .B2(n_464), .Y(n_511) );
OAI211xp5_ASAP7_75t_SL g512 ( .A1(n_488), .A2(n_461), .B(n_459), .C(n_452), .Y(n_512) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_491), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g514 ( .A1(n_499), .A2(n_341), .B1(n_361), .B2(n_467), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_493), .B(n_467), .C(n_421), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_481), .A2(n_397), .B(n_396), .Y(n_516) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_473), .Y(n_517) );
NOR4xp25_ASAP7_75t_L g518 ( .A(n_513), .B(n_478), .C(n_488), .D(n_500), .Y(n_518) );
OAI21xp33_ASAP7_75t_L g519 ( .A1(n_502), .A2(n_495), .B(n_496), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_503), .A2(n_498), .B1(n_485), .B2(n_494), .C(n_490), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_515), .A2(n_482), .B1(n_486), .B2(n_477), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_508), .A2(n_497), .B1(n_424), .B2(n_369), .C(n_396), .Y(n_522) );
AOI211xp5_ASAP7_75t_L g523 ( .A1(n_507), .A2(n_424), .B(n_361), .C(n_390), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_505), .A2(n_361), .B1(n_397), .B2(n_350), .Y(n_524) );
NOR2x1_ASAP7_75t_L g525 ( .A(n_504), .B(n_361), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g526 ( .A(n_509), .B(n_356), .C(n_50), .D(n_51), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_523), .B(n_514), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_520), .A2(n_517), .B1(n_501), .B2(n_516), .C(n_506), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_518), .A2(n_512), .B1(n_517), .B2(n_510), .C(n_511), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_526), .B(n_356), .Y(n_530) );
AOI211xp5_ASAP7_75t_L g531 ( .A1(n_521), .A2(n_254), .B(n_205), .C(n_258), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g532 ( .A1(n_529), .A2(n_525), .B(n_522), .C(n_519), .Y(n_532) );
NAND5xp2_ASAP7_75t_L g533 ( .A(n_528), .B(n_524), .C(n_53), .D(n_55), .E(n_56), .Y(n_533) );
NOR4xp25_ASAP7_75t_L g534 ( .A(n_527), .B(n_49), .C(n_57), .D(n_61), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_532), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_533), .B(n_531), .C(n_530), .Y(n_536) );
OAI22xp5_ASAP7_75t_SL g537 ( .A1(n_535), .A2(n_534), .B1(n_258), .B2(n_67), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_537), .A2(n_536), .B1(n_65), .B2(n_68), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_538), .B(n_63), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_539), .B(n_72), .C(n_73), .Y(n_540) );
AO21x1_ASAP7_75t_L g541 ( .A1(n_540), .A2(n_74), .B(n_75), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_541), .A2(n_76), .B(n_77), .Y(n_542) );
endmodule