module real_aes_9107_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g338 ( .A(n_0), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_1), .A2(n_183), .B1(n_184), .B2(n_188), .Y(n_182) );
INVx1_ASAP7_75t_L g188 ( .A(n_1), .Y(n_188) );
AOI21xp33_ASAP7_75t_L g245 ( .A1(n_2), .A2(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g203 ( .A(n_3), .Y(n_203) );
AND2x6_ASAP7_75t_L g220 ( .A(n_3), .B(n_201), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_3), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_4), .A2(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g254 ( .A(n_5), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_6), .B(n_306), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_7), .A2(n_15), .B1(n_84), .B2(n_101), .Y(n_83) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_8), .A2(n_25), .B1(n_90), .B2(n_95), .Y(n_98) );
INVx1_ASAP7_75t_L g217 ( .A(n_9), .Y(n_217) );
INVx1_ASAP7_75t_L g320 ( .A(n_10), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_11), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_12), .B(n_265), .Y(n_292) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_13), .A2(n_26), .B1(n_90), .B2(n_91), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_14), .B(n_246), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_16), .B(n_242), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_17), .A2(n_27), .B1(n_132), .B2(n_135), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_18), .A2(n_318), .B(n_319), .C(n_321), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_19), .A2(n_80), .B1(n_179), .B2(n_180), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_19), .Y(n_179) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_20), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_21), .B(n_252), .Y(n_339) );
INVx1_ASAP7_75t_L g230 ( .A(n_22), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_22), .A2(n_180), .B1(n_230), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_23), .A2(n_34), .B1(n_120), .B2(n_125), .Y(n_119) );
INVx2_ASAP7_75t_L g224 ( .A(n_24), .Y(n_224) );
OAI221xp5_ASAP7_75t_L g194 ( .A1(n_26), .A2(n_39), .B1(n_47), .B2(n_195), .C(n_196), .Y(n_194) );
INVxp67_ASAP7_75t_L g197 ( .A(n_26), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_28), .A2(n_220), .B(n_231), .C(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g228 ( .A(n_29), .Y(n_228) );
OAI22xp5_ASAP7_75t_SL g184 ( .A1(n_30), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
INVx1_ASAP7_75t_L g187 ( .A(n_30), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_30), .B(n_252), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_31), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_32), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_33), .B(n_246), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_35), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_36), .A2(n_222), .B1(n_225), .B2(n_231), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_37), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_38), .Y(n_335) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_39), .A2(n_55), .B1(n_90), .B2(n_91), .Y(n_89) );
INVxp67_ASAP7_75t_L g198 ( .A(n_39), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_40), .A2(n_251), .B(n_253), .C(n_256), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_41), .Y(n_295) );
INVx1_ASAP7_75t_L g248 ( .A(n_42), .Y(n_248) );
INVx1_ASAP7_75t_L g201 ( .A(n_43), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_44), .A2(n_526), .B1(n_537), .B2(n_538), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_44), .Y(n_537) );
INVx1_ASAP7_75t_L g216 ( .A(n_45), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_46), .Y(n_195) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_47), .A2(n_61), .B1(n_90), .B2(n_95), .Y(n_94) );
A2O1A1Ixp33_ASAP7_75t_SL g264 ( .A1(n_48), .A2(n_256), .B(n_265), .C(n_266), .Y(n_264) );
INVxp67_ASAP7_75t_L g267 ( .A(n_49), .Y(n_267) );
INVx1_ASAP7_75t_L g186 ( .A(n_50), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_51), .Y(n_239) );
INVx1_ASAP7_75t_L g288 ( .A(n_52), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_53), .A2(n_220), .B(n_231), .C(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_54), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_56), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_57), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g214 ( .A(n_58), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_59), .B(n_265), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_60), .A2(n_220), .B(n_231), .C(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_62), .B(n_259), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_63), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_64), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_65), .A2(n_220), .B(n_231), .C(n_303), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_66), .Y(n_310) );
INVx1_ASAP7_75t_L g263 ( .A(n_67), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_68), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_69), .B(n_278), .Y(n_304) );
INVx1_ASAP7_75t_L g90 ( .A(n_70), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_71), .B(n_244), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_72), .A2(n_182), .B1(n_189), .B2(n_190), .Y(n_181) );
INVx1_ASAP7_75t_L g189 ( .A(n_72), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_73), .A2(n_246), .B(n_262), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_74), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_75), .A2(n_76), .B1(n_109), .B2(n_113), .Y(n_108) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_191), .B1(n_204), .B2(n_516), .C(n_524), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_181), .Y(n_78) );
INVx1_ASAP7_75t_L g180 ( .A(n_80), .Y(n_180) );
INVx2_ASAP7_75t_L g538 ( .A(n_80), .Y(n_538) );
AND2x2_ASAP7_75t_SL g80 ( .A(n_81), .B(n_139), .Y(n_80) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_118), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_108), .Y(n_82) );
BUFx3_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_96), .Y(n_86) );
AND2x6_ASAP7_75t_L g105 ( .A(n_87), .B(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g123 ( .A(n_87), .B(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_L g153 ( .A(n_87), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g112 ( .A(n_88), .B(n_94), .Y(n_112) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_89), .B(n_94), .Y(n_117) );
AND2x2_ASAP7_75t_L g129 ( .A(n_89), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g161 ( .A(n_89), .B(n_98), .Y(n_161) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g95 ( .A(n_92), .Y(n_95) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
AND2x4_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g115 ( .A(n_96), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g128 ( .A(n_96), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_99), .Y(n_96) );
OR2x2_ASAP7_75t_L g107 ( .A(n_97), .B(n_100), .Y(n_107) );
AND2x2_ASAP7_75t_L g124 ( .A(n_97), .B(n_100), .Y(n_124) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g154 ( .A(n_98), .B(n_100), .Y(n_154) );
AND2x2_ASAP7_75t_L g159 ( .A(n_99), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g172 ( .A(n_99), .Y(n_172) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g138 ( .A(n_100), .Y(n_138) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx11_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g143 ( .A(n_107), .B(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_112), .B(n_124), .Y(n_148) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g137 ( .A(n_117), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_131), .Y(n_118) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g134 ( .A(n_124), .B(n_129), .Y(n_134) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx8_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx6_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_149), .C(n_168), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B1(n_145), .B2(n_146), .Y(n_140) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI221xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_155), .B1(n_156), .B2(n_162), .C(n_163), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
AND2x4_ASAP7_75t_L g166 ( .A(n_161), .B(n_167), .Y(n_166) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_161), .B(n_172), .Y(n_171) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B1(n_173), .B2(n_174), .Y(n_168) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_180), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_182), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
AND3x1_ASAP7_75t_SL g193 ( .A(n_194), .B(n_199), .C(n_202), .Y(n_193) );
INVxp67_ASAP7_75t_L g530 ( .A(n_194), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx1_ASAP7_75t_SL g532 ( .A(n_199), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_199), .A2(n_519), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g542 ( .A(n_199), .Y(n_542) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_200), .B(n_203), .Y(n_535) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_SL g541 ( .A(n_202), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND3x1_ASAP7_75t_L g205 ( .A(n_206), .B(n_441), .C(n_490), .Y(n_205) );
NOR3xp33_ASAP7_75t_SL g206 ( .A(n_207), .B(n_348), .C(n_386), .Y(n_206) );
OAI222xp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_269), .B1(n_323), .B2(n_329), .C1(n_343), .C2(n_346), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_240), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_209), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_209), .B(n_391), .Y(n_482) );
BUFx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g359 ( .A(n_210), .B(n_260), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_210), .B(n_241), .Y(n_367) );
AND2x2_ASAP7_75t_L g402 ( .A(n_210), .B(n_379), .Y(n_402) );
OR2x2_ASAP7_75t_L g426 ( .A(n_210), .B(n_241), .Y(n_426) );
OR2x2_ASAP7_75t_L g434 ( .A(n_210), .B(n_333), .Y(n_434) );
AND2x2_ASAP7_75t_L g437 ( .A(n_210), .B(n_260), .Y(n_437) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g331 ( .A(n_211), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g345 ( .A(n_211), .B(n_260), .Y(n_345) );
AND2x2_ASAP7_75t_L g395 ( .A(n_211), .B(n_333), .Y(n_395) );
AND2x2_ASAP7_75t_L g408 ( .A(n_211), .B(n_241), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_211), .B(n_494), .Y(n_515) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_238), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_212), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_212), .A2(n_334), .B(n_341), .Y(n_333) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_213), .Y(n_244) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x2_ASAP7_75t_SL g259 ( .A(n_214), .B(n_215), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_221), .B1(n_234), .B2(n_235), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_219), .A2(n_248), .B(n_249), .C(n_250), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_219), .A2(n_249), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_219), .A2(n_249), .B(n_316), .C(n_317), .Y(n_315) );
INVx4_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_220), .B(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g246 ( .A(n_220), .B(n_236), .Y(n_246) );
BUFx3_ASAP7_75t_L g518 ( .A(n_220), .Y(n_518) );
INVx2_ASAP7_75t_L g340 ( .A(n_222), .Y(n_340) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g232 ( .A(n_224), .Y(n_232) );
INVx1_ASAP7_75t_L g237 ( .A(n_224), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g225 ( .A1(n_226), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_225) );
INVx2_ASAP7_75t_L g229 ( .A(n_226), .Y(n_229) );
INVx4_ASAP7_75t_L g318 ( .A(n_226), .Y(n_318) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
AND2x2_ASAP7_75t_L g236 ( .A(n_227), .B(n_237), .Y(n_236) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_227), .Y(n_252) );
INVx3_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
INVx1_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
OAI322xp33_ASAP7_75t_L g524 ( .A1(n_228), .A2(n_525), .A3(n_527), .B1(n_531), .B2(n_533), .C1(n_536), .C2(n_539), .Y(n_524) );
INVx2_ASAP7_75t_L g523 ( .A(n_229), .Y(n_523) );
INVx5_ASAP7_75t_L g249 ( .A(n_231), .Y(n_249) );
AND2x6_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_232), .Y(n_257) );
BUFx3_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_235), .A2(n_288), .B(n_289), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_235), .A2(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g521 ( .A(n_237), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_240), .A2(n_434), .B(n_435), .C(n_438), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_240), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_240), .B(n_378), .Y(n_500) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_260), .Y(n_240) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_241), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g358 ( .A(n_241), .Y(n_358) );
AND2x2_ASAP7_75t_L g385 ( .A(n_241), .B(n_379), .Y(n_385) );
INVx1_ASAP7_75t_SL g393 ( .A(n_241), .Y(n_393) );
AND2x2_ASAP7_75t_L g416 ( .A(n_241), .B(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g494 ( .A(n_241), .Y(n_494) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_245), .B(n_258), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_243), .B(n_285), .Y(n_284) );
INVx4_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_244), .A2(n_261), .B(n_268), .Y(n_260) );
BUFx2_ASAP7_75t_L g314 ( .A(n_246), .Y(n_314) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx4_ASAP7_75t_L g306 ( .A(n_252), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_255), .B(n_267), .Y(n_266) );
INVx5_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_257), .Y(n_307) );
INVx1_ASAP7_75t_L g296 ( .A(n_259), .Y(n_296) );
INVx2_ASAP7_75t_L g300 ( .A(n_259), .Y(n_300) );
OA21x2_ASAP7_75t_L g312 ( .A1(n_259), .A2(n_313), .B(n_322), .Y(n_312) );
BUFx2_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
INVx1_ASAP7_75t_L g392 ( .A(n_260), .Y(n_392) );
INVx3_ASAP7_75t_L g417 ( .A(n_260), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_269), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_297), .Y(n_269) );
INVx1_ASAP7_75t_L g413 ( .A(n_270), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g419 ( .A1(n_270), .A2(n_358), .A3(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_270), .A2(n_424), .B1(n_427), .B2(n_432), .Y(n_423) );
INVx4_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g361 ( .A(n_271), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g439 ( .A(n_271), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g509 ( .A(n_271), .B(n_455), .Y(n_509) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_286), .Y(n_271) );
AND2x2_ASAP7_75t_L g324 ( .A(n_272), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g354 ( .A(n_272), .Y(n_354) );
INVx1_ASAP7_75t_L g373 ( .A(n_272), .Y(n_373) );
OR2x2_ASAP7_75t_L g381 ( .A(n_272), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_272), .B(n_362), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_272), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g409 ( .A(n_272), .B(n_327), .Y(n_409) );
INVx3_ASAP7_75t_L g431 ( .A(n_272), .Y(n_431) );
AND2x2_ASAP7_75t_L g456 ( .A(n_272), .B(n_328), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_272), .B(n_421), .Y(n_504) );
OR2x6_ASAP7_75t_L g272 ( .A(n_273), .B(n_284), .Y(n_272) );
AOI21xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_275), .B(n_283), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B(n_280), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_278), .A2(n_338), .B(n_339), .C(n_340), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_280), .A2(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
INVx1_ASAP7_75t_L g293 ( .A(n_283), .Y(n_293) );
INVx2_ASAP7_75t_L g328 ( .A(n_286), .Y(n_328) );
AND2x2_ASAP7_75t_L g460 ( .A(n_286), .B(n_298), .Y(n_460) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_293), .B(n_294), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_296), .B(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_296), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g502 ( .A(n_297), .Y(n_502) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_311), .Y(n_297) );
INVx1_ASAP7_75t_L g347 ( .A(n_298), .Y(n_347) );
AND2x2_ASAP7_75t_L g374 ( .A(n_298), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_298), .B(n_328), .Y(n_382) );
AND2x2_ASAP7_75t_L g440 ( .A(n_298), .B(n_363), .Y(n_440) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_299), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g362 ( .A(n_299), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_299), .B(n_328), .Y(n_428) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_309), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_307), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_311), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g375 ( .A(n_311), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_311), .B(n_328), .Y(n_421) );
AND2x2_ASAP7_75t_L g430 ( .A(n_311), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g455 ( .A(n_311), .Y(n_455) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g327 ( .A(n_312), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_318), .B(n_320), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_323), .A2(n_333), .B1(n_492), .B2(n_495), .Y(n_491) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
OAI21xp5_ASAP7_75t_SL g514 ( .A1(n_325), .A2(n_436), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_326), .B(n_431), .Y(n_448) );
INVx1_ASAP7_75t_L g473 ( .A(n_326), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_327), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g400 ( .A(n_327), .B(n_353), .Y(n_400) );
INVx2_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
INVx1_ASAP7_75t_L g406 ( .A(n_328), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g497 ( .A1(n_329), .A2(n_481), .B1(n_498), .B2(n_501), .C(n_503), .Y(n_497) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g368 ( .A(n_330), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_330), .B(n_379), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_331), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g422 ( .A(n_331), .B(n_368), .Y(n_422) );
INVx3_ASAP7_75t_SL g463 ( .A(n_331), .Y(n_463) );
AND2x2_ASAP7_75t_L g407 ( .A(n_332), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g436 ( .A(n_332), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_332), .B(n_345), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_332), .B(n_391), .Y(n_477) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g379 ( .A(n_333), .Y(n_379) );
OAI322xp33_ASAP7_75t_L g474 ( .A1(n_333), .A2(n_405), .A3(n_427), .B1(n_475), .B2(n_477), .C1(n_478), .C2(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI21xp33_ASAP7_75t_L g498 ( .A1(n_344), .A2(n_347), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_SL g424 ( .A(n_345), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g446 ( .A(n_345), .B(n_358), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_345), .B(n_385), .Y(n_461) );
INVxp67_ASAP7_75t_L g412 ( .A(n_347), .Y(n_412) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_347), .A2(n_419), .B(n_423), .C(n_433), .Y(n_418) );
OAI221xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_357), .B1(n_360), .B2(n_364), .C(n_369), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g372 ( .A(n_356), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g489 ( .A(n_356), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_357), .A2(n_506), .B1(n_511), .B2(n_512), .C(n_514), .Y(n_505) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_358), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_358), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_358), .B(n_436), .Y(n_443) );
AND2x2_ASAP7_75t_L g485 ( .A(n_358), .B(n_463), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_359), .B(n_384), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_359), .A2(n_371), .B1(n_481), .B2(n_482), .Y(n_480) );
OR2x2_ASAP7_75t_L g511 ( .A(n_359), .B(n_379), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g488 ( .A(n_362), .Y(n_488) );
AND2x2_ASAP7_75t_L g513 ( .A(n_362), .B(n_456), .Y(n_513) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g377 ( .A(n_367), .B(n_378), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_376), .B1(n_380), .B2(n_383), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g444 ( .A(n_372), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_372), .B(n_412), .Y(n_479) );
AOI322xp5_ASAP7_75t_L g403 ( .A1(n_374), .A2(n_404), .A3(n_406), .B1(n_407), .B2(n_409), .C1(n_410), .C2(n_414), .Y(n_403) );
INVxp67_ASAP7_75t_L g397 ( .A(n_375), .Y(n_397) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_377), .A2(n_382), .B1(n_399), .B2(n_401), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_378), .B(n_391), .Y(n_478) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_379), .B(n_417), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_379), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g475 ( .A(n_381), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NAND3xp33_ASAP7_75t_SL g386 ( .A(n_387), .B(n_403), .C(n_418), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_394), .B2(n_396), .C(n_398), .Y(n_387) );
AND2x2_ASAP7_75t_L g394 ( .A(n_390), .B(n_395), .Y(n_394) );
INVx3_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AND2x2_ASAP7_75t_L g404 ( .A(n_395), .B(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_397), .Y(n_476) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_402), .B(n_416), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_405), .B(n_463), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_406), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g481 ( .A(n_409), .Y(n_481) );
AND2x2_ASAP7_75t_L g496 ( .A(n_409), .B(n_473), .Y(n_496) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g490 ( .A1(n_420), .A2(n_491), .B(n_497), .C(n_505), .Y(n_490) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g459 ( .A(n_430), .B(n_460), .Y(n_459) );
NAND2x1_ASAP7_75t_SL g501 ( .A(n_431), .B(n_502), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_434), .Y(n_471) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g466 ( .A(n_440), .Y(n_466) );
AND2x2_ASAP7_75t_L g470 ( .A(n_440), .B(n_456), .Y(n_470) );
NOR5xp2_ASAP7_75t_L g441 ( .A(n_442), .B(n_457), .C(n_474), .D(n_480), .E(n_483), .Y(n_441) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_445), .B2(n_447), .C(n_449), .Y(n_442) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_446), .B(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g472 ( .A(n_456), .B(n_473), .Y(n_472) );
OAI221xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_461), .B1(n_462), .B2(n_464), .C(n_467), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g510 ( .A(n_470), .Y(n_510) );
AOI211xp5_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_486), .B(n_488), .C(n_489), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
CKINVDCx14_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
endmodule