module fake_ibex_369_n_1765 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_340, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1765);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1765;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_504;
wire n_1752;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1599;
wire n_1400;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_1455;
wire n_484;
wire n_1642;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1740;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_1744;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1755;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_341),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_342),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_296),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_148),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_97),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_319),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_193),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_202),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_80),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_0),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_150),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_346),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_299),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_117),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_47),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_146),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_232),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_236),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_133),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_45),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_256),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_110),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_52),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_180),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_287),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_190),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_265),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_297),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_253),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_165),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_282),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_8),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_246),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_63),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_262),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_260),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_138),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_55),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_32),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_144),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_111),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_276),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_38),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_63),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_82),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_69),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_178),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_251),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_35),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_4),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_137),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_340),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_54),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_122),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_66),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_288),
.Y(n_408)
);

BUFx12f_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_126),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_266),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_277),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_120),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_305),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_343),
.Y(n_415)
);

BUFx10_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_61),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_344),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_145),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_113),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_302),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_189),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_300),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_18),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_283),
.Y(n_425)
);

BUFx8_ASAP7_75t_SL g426 ( 
.A(n_261),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_285),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_314),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_68),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_57),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_87),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_224),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_87),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_125),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_244),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_159),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_307),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_321),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_248),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_183),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_80),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_255),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_243),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_194),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_128),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_281),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_269),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_184),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_8),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_263),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_208),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_286),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_3),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_268),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_112),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_51),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_279),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_149),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_324),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_270),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_75),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_301),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_152),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_161),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_136),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_195),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_271),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_304),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_325),
.Y(n_469)
);

INVxp33_ASAP7_75t_R g470 ( 
.A(n_201),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_293),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_188),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_337),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_220),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_249),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_294),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_257),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_218),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_105),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_290),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_13),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_105),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_309),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_348),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_311),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_316),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_9),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_280),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_345),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_64),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_223),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_242),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_143),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_181),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_313),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_328),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_315),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_54),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_68),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_221),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_103),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_259),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_252),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_185),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_3),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_318),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_216),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_92),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_187),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_240),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_39),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_151),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_231),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_0),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_121),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_23),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_349),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_13),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_326),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_52),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_308),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_237),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_85),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_196),
.Y(n_524)
);

BUFx5_ASAP7_75t_L g525 ( 
.A(n_65),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_267),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_203),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_40),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_39),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_62),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_176),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_339),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_320),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_306),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_92),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_219),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_327),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_99),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_114),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_55),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_274),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_12),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_291),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_254),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_51),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_264),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_317),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_278),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_70),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_167),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_61),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_250),
.Y(n_552)
);

BUFx8_ASAP7_75t_SL g553 ( 
.A(n_79),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_273),
.Y(n_554)
);

CKINVDCx14_ASAP7_75t_R g555 ( 
.A(n_78),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_258),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_11),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_292),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_275),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_206),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_147),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_50),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_303),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_334),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_94),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_310),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_49),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_245),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_169),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_107),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_57),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_59),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_338),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_60),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_64),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_32),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_347),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_157),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_289),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_168),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_24),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_4),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_199),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_312),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_59),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_142),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_31),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_272),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_333),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_298),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_62),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_335),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_247),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_329),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_284),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_72),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_7),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_139),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_295),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_336),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_2),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_28),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_173),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_426),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_369),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_371),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_L g607 ( 
.A(n_490),
.B(n_1),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_354),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_444),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_445),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_380),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_476),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_555),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_555),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_477),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_484),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_536),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_525),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_372),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_427),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_581),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_527),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_384),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_525),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_378),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_499),
.B(n_572),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_499),
.B(n_1),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_390),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_466),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_354),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_500),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_407),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_502),
.Y(n_634)
);

INVxp33_ASAP7_75t_SL g635 ( 
.A(n_359),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_435),
.B(n_2),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_409),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_382),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_382),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_549),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_409),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_562),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_553),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_414),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_585),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_585),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_582),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_414),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_581),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_370),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_438),
.B(n_5),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_581),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_525),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_375),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_525),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_525),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_373),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_375),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_360),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_397),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_400),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_365),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_389),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_405),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_417),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_424),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_394),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_396),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_401),
.Y(n_672)
);

INVxp33_ASAP7_75t_SL g673 ( 
.A(n_441),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_429),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_456),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_430),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_431),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_433),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_449),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_479),
.Y(n_680)
);

BUFx6f_ASAP7_75t_SL g681 ( 
.A(n_416),
.Y(n_681)
);

CKINVDCx16_ASAP7_75t_R g682 ( 
.A(n_416),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_453),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_461),
.B(n_5),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_481),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_605),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_606),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_633),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_609),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_610),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_657),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_633),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_608),
.B(n_388),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_613),
.B(n_416),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_619),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_638),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_619),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_639),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_625),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_658),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_640),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_660),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_625),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_612),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_648),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_657),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_640),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_685),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_616),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_617),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_655),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_618),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_656),
.Y(n_714)
);

AND3x2_ASAP7_75t_L g715 ( 
.A(n_622),
.B(n_470),
.C(n_432),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_665),
.B(n_388),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_604),
.B(n_350),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_645),
.B(n_454),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_652),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_659),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_661),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_666),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_642),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_664),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_646),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_647),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_670),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_682),
.B(n_454),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_611),
.B(n_520),
.Y(n_731)
);

CKINVDCx14_ASAP7_75t_R g732 ( 
.A(n_654),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_614),
.B(n_528),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_664),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_651),
.B(n_454),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_672),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_677),
.B(n_482),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_674),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_615),
.B(n_351),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_669),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_636),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_676),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_643),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_663),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_621),
.B(n_420),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_683),
.B(n_487),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_669),
.Y(n_750)
);

BUFx10_ASAP7_75t_L g751 ( 
.A(n_681),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_681),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_662),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_667),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_615),
.B(n_654),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_680),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_650),
.B(n_460),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_627),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_680),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_628),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_681),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_643),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_653),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_607),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_623),
.Y(n_766)
);

XNOR2xp5_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_498),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_668),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_624),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_675),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_637),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_629),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_673),
.B(n_402),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_641),
.B(n_402),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_620),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_626),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_630),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_632),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_634),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_644),
.B(n_352),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_649),
.B(n_567),
.C(n_557),
.Y(n_781)
);

OA21x2_ASAP7_75t_L g782 ( 
.A1(n_648),
.A2(n_437),
.B(n_434),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_608),
.B(n_434),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_605),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_657),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_605),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_657),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_605),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_605),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_619),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_613),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_631),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_605),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_633),
.Y(n_794)
);

BUFx8_ASAP7_75t_L g795 ( 
.A(n_681),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_645),
.B(n_353),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_619),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_605),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_654),
.A2(n_501),
.B1(n_508),
.B2(n_505),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_619),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_611),
.B(n_574),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_613),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_631),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_605),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_657),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_660),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_631),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_608),
.B(n_437),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_608),
.B(n_443),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_657),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_605),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_631),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_621),
.B(n_357),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_657),
.Y(n_816)
);

BUFx8_ASAP7_75t_L g817 ( 
.A(n_681),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_619),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_613),
.B(n_511),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_657),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_657),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_619),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_R g823 ( 
.A(n_604),
.B(n_514),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_608),
.B(n_443),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_605),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_631),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_613),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_605),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_605),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_633),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_731),
.A2(n_518),
.B1(n_523),
.B2(n_516),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_722),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_751),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_703),
.B(n_529),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_785),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_795),
.B(n_530),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_730),
.B(n_355),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_692),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_764),
.B(n_473),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_692),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_782),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_751),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_781),
.B(n_597),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_703),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_806),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_709),
.B(n_535),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_752),
.B(n_729),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_709),
.B(n_538),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_762),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_692),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_719),
.B(n_540),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_741),
.B(n_395),
.Y(n_852)
);

INVx8_ASAP7_75t_L g853 ( 
.A(n_752),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_762),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_785),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_782),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_721),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_731),
.B(n_733),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_733),
.A2(n_545),
.B1(n_551),
.B2(n_542),
.Y(n_859)
);

INVx6_ASAP7_75t_L g860 ( 
.A(n_795),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_688),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_802),
.B(n_552),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_743),
.B(n_356),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_805),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_805),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_812),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_719),
.B(n_602),
.Y(n_867)
);

OAI22xp33_ASAP7_75t_L g868 ( 
.A1(n_799),
.A2(n_565),
.B1(n_575),
.B2(n_571),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_791),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_801),
.A2(n_587),
.B1(n_591),
.B2(n_576),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_801),
.B(n_596),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_707),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_812),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_707),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_735),
.B(n_358),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_827),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_816),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_827),
.B(n_601),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_730),
.B(n_361),
.Y(n_879)
);

INVx5_ASAP7_75t_L g880 ( 
.A(n_707),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_787),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_721),
.Y(n_882)
);

AND3x4_ASAP7_75t_L g883 ( 
.A(n_781),
.B(n_475),
.C(n_457),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_775),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_802),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_L g886 ( 
.A(n_738),
.B(n_366),
.C(n_362),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_787),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_816),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_820),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_820),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_817),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_787),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_730),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_755),
.B(n_590),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_807),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_749),
.B(n_395),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_817),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_769),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_807),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_743),
.B(n_367),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_766),
.B(n_363),
.Y(n_901)
);

INVx4_ASAP7_75t_SL g902 ( 
.A(n_743),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_690),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_701),
.A2(n_395),
.B1(n_368),
.B2(n_386),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_807),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_753),
.B(n_364),
.Y(n_906)
);

AND2x6_ASAP7_75t_L g907 ( 
.A(n_695),
.B(n_377),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_819),
.B(n_754),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_821),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_754),
.B(n_395),
.Y(n_910)
);

AND3x1_ASAP7_75t_L g911 ( 
.A(n_776),
.B(n_403),
.C(n_393),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_799),
.B(n_410),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_821),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_773),
.B(n_374),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_697),
.Y(n_915)
);

OR2x6_ASAP7_75t_L g916 ( 
.A(n_746),
.B(n_411),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_821),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_768),
.B(n_413),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_724),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_726),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_758),
.B(n_376),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_727),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_768),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_699),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_773),
.B(n_379),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_723),
.B(n_381),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_792),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_747),
.A2(n_815),
.B1(n_736),
.B2(n_739),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_803),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_747),
.B(n_423),
.C(n_419),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_728),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_777),
.B(n_428),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_770),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_771),
.B(n_383),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_809),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_814),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_826),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_694),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_770),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_737),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_744),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_748),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_696),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_759),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_698),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_716),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_765),
.B(n_436),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_716),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_694),
.B(n_385),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_686),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_778),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_779),
.B(n_6),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_783),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_783),
.A2(n_446),
.B1(n_448),
.B2(n_442),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_774),
.B(n_387),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_700),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_810),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_704),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_718),
.B(n_391),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_790),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_761),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_797),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_796),
.B(n_392),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_772),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_810),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_774),
.B(n_450),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_811),
.B(n_398),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_800),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_779),
.B(n_399),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_725),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_811),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_824),
.B(n_452),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_715),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_808),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_734),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_818),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_742),
.B(n_6),
.Y(n_977)
);

AND2x6_ASAP7_75t_L g978 ( 
.A(n_824),
.B(n_455),
.Y(n_978)
);

AND2x6_ASAP7_75t_L g979 ( 
.A(n_706),
.B(n_471),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_712),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_822),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_720),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_715),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_714),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_687),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_717),
.B(n_404),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_689),
.B(n_472),
.Y(n_987)
);

BUFx10_ASAP7_75t_L g988 ( 
.A(n_691),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_740),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_780),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_705),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_710),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_711),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_713),
.B(n_485),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_784),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_823),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_786),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_788),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_756),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_789),
.B(n_406),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_793),
.B(n_408),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_750),
.B(n_7),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_798),
.B(n_412),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_757),
.B(n_9),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_804),
.A2(n_492),
.B1(n_493),
.B2(n_489),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_813),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_825),
.B(n_497),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_760),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_828),
.B(n_415),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_829),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_732),
.B(n_507),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_767),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_693),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_702),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_708),
.Y(n_1015)
);

AO21x2_ASAP7_75t_L g1016 ( 
.A1(n_745),
.A2(n_513),
.B(n_510),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_763),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_794),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_830),
.B(n_418),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_751),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_743),
.B(n_421),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_795),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_795),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_722),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_722),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_751),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_785),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_785),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_785),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_751),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_795),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_785),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_806),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_703),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_722),
.Y(n_1035)
);

AND2x6_ASAP7_75t_L g1036 ( 
.A(n_752),
.B(n_515),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_692),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_795),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_806),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_751),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_692),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_785),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_703),
.B(n_603),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_795),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_731),
.A2(n_580),
.B1(n_583),
.B2(n_573),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_795),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_731),
.B(n_593),
.Y(n_1047)
);

AND2x6_ASAP7_75t_L g1048 ( 
.A(n_752),
.B(n_457),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_751),
.Y(n_1049)
);

INVxp33_ASAP7_75t_SL g1050 ( 
.A(n_756),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_743),
.B(n_422),
.Y(n_1051)
);

BUFx10_ASAP7_75t_L g1052 ( 
.A(n_775),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_730),
.B(n_425),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_692),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_751),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_938),
.B(n_439),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_938),
.B(n_440),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_957),
.B(n_946),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_957),
.B(n_447),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_860),
.B(n_475),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_948),
.B(n_953),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_876),
.B(n_451),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_869),
.B(n_458),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_860),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_941),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_965),
.B(n_459),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_883),
.A2(n_541),
.B1(n_569),
.B2(n_478),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_922),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_923),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_971),
.B(n_462),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_885),
.B(n_463),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_892),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_858),
.B(n_933),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_858),
.B(n_464),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_941),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_843),
.A2(n_541),
.B1(n_569),
.B2(n_478),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_871),
.B(n_465),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_942),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_922),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_972),
.B(n_467),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_871),
.B(n_468),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_951),
.B(n_469),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_942),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_960),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_972),
.A2(n_978),
.B1(n_912),
.B2(n_966),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_960),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_972),
.B(n_474),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_867),
.B(n_10),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_912),
.A2(n_589),
.B1(n_595),
.B2(n_577),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_1055),
.B(n_833),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_978),
.B(n_480),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_SL g1092 ( 
.A(n_891),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_978),
.B(n_483),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_928),
.B(n_486),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_940),
.B(n_488),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_919),
.B(n_491),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1047),
.B(n_494),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1039),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_974),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1047),
.B(n_495),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_974),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1034),
.B(n_496),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_903),
.B(n_927),
.Y(n_1103)
);

O2A1O1Ixp5_ASAP7_75t_L g1104 ( 
.A1(n_955),
.A2(n_589),
.B(n_595),
.C(n_577),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_923),
.Y(n_1105)
);

INVx8_ASAP7_75t_L g1106 ( 
.A(n_852),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1026),
.B(n_503),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_896),
.Y(n_1108)
);

INVxp33_ASAP7_75t_L g1109 ( 
.A(n_939),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1031),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_903),
.B(n_504),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_966),
.A2(n_600),
.B1(n_509),
.B2(n_512),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_844),
.B(n_10),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_976),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_927),
.B(n_506),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_862),
.B(n_517),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_915),
.B(n_519),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_976),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_892),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_981),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_863),
.A2(n_600),
.B(n_522),
.C(n_524),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_1044),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_929),
.B(n_521),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_836),
.A2(n_918),
.B1(n_916),
.B2(n_997),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_980),
.A2(n_531),
.B1(n_533),
.B2(n_532),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_SL g1126 ( 
.A(n_1008),
.B(n_537),
.C(n_534),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_845),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_935),
.B(n_539),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_841),
.A2(n_544),
.B(n_543),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_937),
.B(n_546),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_908),
.B(n_11),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_949),
.B(n_547),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_982),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_909),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1026),
.B(n_1040),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_SL g1136 ( 
.A(n_833),
.B(n_548),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_878),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_909),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_875),
.A2(n_550),
.B1(n_556),
.B2(n_554),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_967),
.B(n_558),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_832),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_918),
.A2(n_559),
.B1(n_561),
.B2(n_560),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_875),
.A2(n_563),
.B1(n_566),
.B2(n_564),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_875),
.B(n_931),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_897),
.Y(n_1145)
);

INVxp67_ASAP7_75t_SL g1146 ( 
.A(n_1033),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1046),
.Y(n_1147)
);

OAI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_831),
.A2(n_570),
.B1(n_579),
.B2(n_578),
.C(n_568),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_832),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1011),
.A2(n_594),
.B1(n_598),
.B2(n_586),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_981),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_924),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_936),
.B(n_599),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_920),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1043),
.B(n_979),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1024),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_979),
.B(n_12),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1024),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1025),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_979),
.B(n_907),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_907),
.B(n_14),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1025),
.Y(n_1162)
);

AND3x1_ASAP7_75t_L g1163 ( 
.A(n_973),
.B(n_14),
.C(n_15),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_907),
.B(n_15),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1040),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_842),
.B(n_16),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_868),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1049),
.B(n_526),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1035),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1035),
.A2(n_584),
.B1(n_588),
.B2(n_526),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_894),
.B(n_17),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1049),
.B(n_526),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_842),
.B(n_19),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_851),
.B(n_19),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_910),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_857),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_835),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_852),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_932),
.A2(n_584),
.B1(n_526),
.B2(n_588),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1055),
.B(n_584),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_SL g1181 ( 
.A(n_997),
.B(n_584),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_839),
.B(n_20),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_834),
.B(n_846),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_864),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_932),
.A2(n_588),
.B1(n_22),
.B2(n_20),
.Y(n_1185)
);

NOR2xp67_ASAP7_75t_L g1186 ( 
.A(n_996),
.B(n_21),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_932),
.A2(n_588),
.B1(n_23),
.B2(n_21),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_865),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_866),
.Y(n_1189)
);

XOR2xp5_ASAP7_75t_L g1190 ( 
.A(n_861),
.B(n_22),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1045),
.B(n_24),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_893),
.B(n_25),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_857),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_954),
.B(n_25),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_947),
.B(n_26),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_873),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1011),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_911),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_882),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1022),
.B(n_29),
.Y(n_1200)
);

INVxp67_ASAP7_75t_SL g1201 ( 
.A(n_841),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_947),
.B(n_30),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_882),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_877),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_944),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_856),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_848),
.B(n_33),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_917),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_886),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_969),
.B(n_855),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_981),
.B(n_36),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_888),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_889),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_902),
.B(n_37),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_856),
.A2(n_109),
.B(n_108),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_890),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_849),
.B(n_37),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1036),
.B(n_38),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1036),
.B(n_900),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1036),
.B(n_40),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_900),
.B(n_41),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1027),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_916),
.B(n_41),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1028),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_950),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_902),
.B(n_996),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_884),
.B(n_42),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_854),
.B(n_1020),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_900),
.B(n_42),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_930),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_984),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_901),
.B(n_46),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_987),
.B(n_47),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_996),
.B(n_48),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1014),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1013),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_987),
.B(n_48),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1023),
.B(n_49),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1029),
.A2(n_56),
.B1(n_50),
.B2(n_53),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1032),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1038),
.B(n_53),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_859),
.B(n_56),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_R g1243 ( 
.A(n_1235),
.B(n_1015),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1061),
.B(n_847),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1145),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1133),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1072),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1109),
.B(n_1018),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1090),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1069),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1072),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1058),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1141),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1152),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1105),
.B(n_847),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1145),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1149),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1064),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1072),
.Y(n_1259)
);

INVx5_ASAP7_75t_L g1260 ( 
.A(n_1106),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1183),
.B(n_847),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1205),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1124),
.B(n_998),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1106),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_1179),
.B(n_1067),
.C(n_1085),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1122),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1106),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1065),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1165),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1103),
.B(n_983),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1165),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1098),
.B(n_1010),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1131),
.B(n_1016),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1073),
.B(n_870),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1208),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1208),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1158),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1075),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1078),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1083),
.B(n_994),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1110),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1137),
.B(n_1017),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1147),
.B(n_964),
.C(n_898),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1092),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1159),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1208),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1174),
.B(n_994),
.Y(n_1287)
);

AND3x1_ASAP7_75t_SL g1288 ( 
.A(n_1190),
.B(n_995),
.C(n_993),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1156),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1166),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1076),
.B(n_1007),
.Y(n_1291)
);

NOR3xp33_ASAP7_75t_SL g1292 ( 
.A(n_1223),
.B(n_975),
.C(n_970),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1076),
.B(n_1007),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1136),
.A2(n_1050),
.B1(n_993),
.B2(n_995),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1166),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1173),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1136),
.A2(n_992),
.B1(n_985),
.B2(n_991),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1238),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1175),
.B(n_952),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1162),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1142),
.B(n_884),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1181),
.B(n_1052),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1146),
.B(n_1030),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1084),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1201),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1154),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1228),
.B(n_1006),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1084),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1169),
.B(n_961),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1101),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1177),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1113),
.B(n_914),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1101),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1181),
.B(n_1173),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1184),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1222),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1188),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1120),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1060),
.Y(n_1319)
);

AND3x1_ASAP7_75t_SL g1320 ( 
.A(n_1148),
.B(n_990),
.C(n_989),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1228),
.B(n_999),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1108),
.B(n_925),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1238),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1207),
.B(n_1155),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1060),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1238),
.B(n_1013),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1225),
.B(n_1042),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1060),
.B(n_1021),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1189),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1217),
.Y(n_1330)
);

AND3x2_ASAP7_75t_SL g1331 ( 
.A(n_1163),
.B(n_1052),
.C(n_988),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1224),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1196),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1200),
.A2(n_1012),
.B1(n_983),
.B2(n_1002),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1240),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1120),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_R g1337 ( 
.A(n_1126),
.B(n_988),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1077),
.B(n_1019),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1204),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1233),
.A2(n_1063),
.B1(n_1062),
.B2(n_1102),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1176),
.Y(n_1341)
);

AND2x6_ASAP7_75t_SL g1342 ( 
.A(n_1227),
.B(n_1003),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1151),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1151),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1150),
.B(n_986),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1217),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1086),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1178),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1127),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1212),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_R g1351 ( 
.A(n_1236),
.B(n_1011),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1099),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1089),
.B(n_1005),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1114),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1193),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1210),
.B(n_1051),
.Y(n_1356)
);

AND2x4_ASAP7_75t_SL g1357 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1199),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1089),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1135),
.B(n_934),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1088),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1056),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1242),
.A2(n_1004),
.B1(n_977),
.B2(n_1048),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1203),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1125),
.B(n_837),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1057),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1059),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1097),
.B(n_1000),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1213),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1216),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1068),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1094),
.B(n_1191),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1186),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1079),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1119),
.Y(n_1375)
);

AND2x2_ASAP7_75t_SL g1376 ( 
.A(n_1163),
.B(n_1001),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1144),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1198),
.B(n_879),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1081),
.B(n_906),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1161),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1164),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1195),
.B(n_853),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1160),
.B(n_874),
.Y(n_1383)
);

NAND2xp33_ASAP7_75t_SL g1384 ( 
.A(n_1219),
.B(n_1053),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1237),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1194),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1134),
.Y(n_1387)
);

AO22x2_ASAP7_75t_L g1388 ( 
.A1(n_1263),
.A2(n_1206),
.B1(n_1234),
.B2(n_1157),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1202),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1314),
.A2(n_1215),
.B(n_1104),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1291),
.B(n_1112),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1258),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1293),
.B(n_1082),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1253),
.A2(n_1226),
.B(n_1138),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1260),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1273),
.A2(n_1230),
.A3(n_1232),
.B(n_1182),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1257),
.A2(n_1192),
.B(n_1180),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1277),
.A2(n_1172),
.B(n_1168),
.Y(n_1398)
);

AOI211x1_ASAP7_75t_L g1399 ( 
.A1(n_1274),
.A2(n_1171),
.B(n_1214),
.C(n_1211),
.Y(n_1399)
);

INVx3_ASAP7_75t_SL g1400 ( 
.A(n_1266),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1298),
.B(n_1198),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1359),
.B(n_1125),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1305),
.A2(n_1231),
.B1(n_1239),
.B2(n_1187),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1287),
.B(n_1066),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1285),
.A2(n_1170),
.B(n_840),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1386),
.A2(n_1229),
.A3(n_1221),
.B(n_1220),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1319),
.B(n_1325),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1372),
.B(n_1070),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1246),
.B(n_1071),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1302),
.A2(n_1170),
.B(n_850),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1338),
.B(n_1074),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1260),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1262),
.Y(n_1413)
);

BUFx8_ASAP7_75t_L g1414 ( 
.A(n_1245),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1268),
.B(n_1100),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1250),
.B(n_1361),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1260),
.B(n_1241),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1346),
.A2(n_1231),
.B1(n_1239),
.B2(n_1185),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_874),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1365),
.A2(n_1115),
.B(n_1111),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1289),
.A2(n_872),
.B(n_838),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1319),
.B(n_1129),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1290),
.B(n_921),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1300),
.A2(n_887),
.B(n_881),
.Y(n_1424)
);

O2A1O1Ixp5_ASAP7_75t_L g1425 ( 
.A1(n_1270),
.A2(n_1218),
.B(n_1121),
.C(n_1107),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1341),
.A2(n_913),
.B(n_895),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1330),
.A2(n_1197),
.B1(n_1209),
.B2(n_1139),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1324),
.A2(n_1167),
.B(n_1123),
.C(n_1128),
.Y(n_1428)
);

NOR2x1_ASAP7_75t_L g1429 ( 
.A(n_1256),
.B(n_1080),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1384),
.A2(n_1140),
.B(n_1132),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1264),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1244),
.A2(n_1130),
.B(n_1117),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1264),
.B(n_874),
.Y(n_1433)
);

AOI21xp33_ASAP7_75t_L g1434 ( 
.A1(n_1340),
.A2(n_1116),
.B(n_1091),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1355),
.A2(n_1041),
.B(n_1037),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1278),
.B(n_963),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1279),
.B(n_1252),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1267),
.Y(n_1438)
);

AOI31xp67_ASAP7_75t_L g1439 ( 
.A1(n_1345),
.A2(n_1054),
.A3(n_945),
.B(n_956),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1280),
.B(n_959),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1358),
.A2(n_905),
.B(n_899),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1267),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1254),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1261),
.A2(n_1153),
.B(n_1095),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1265),
.A2(n_904),
.B(n_943),
.Y(n_1445)
);

AO31x2_ASAP7_75t_L g1446 ( 
.A1(n_1364),
.A2(n_958),
.A3(n_968),
.B(n_962),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1296),
.A2(n_1143),
.B1(n_1087),
.B2(n_1093),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1373),
.A2(n_1096),
.B(n_926),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1282),
.A2(n_1048),
.B1(n_853),
.B2(n_880),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1376),
.A2(n_880),
.B(n_1048),
.C(n_65),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1311),
.A2(n_880),
.B(n_116),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1379),
.B(n_58),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1309),
.A2(n_1312),
.B(n_1378),
.Y(n_1453)
);

AOI211x1_ASAP7_75t_L g1454 ( 
.A1(n_1301),
.A2(n_66),
.B(n_58),
.C(n_60),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1325),
.B(n_67),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1249),
.B(n_67),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1306),
.Y(n_1457)
);

AO31x2_ASAP7_75t_L g1458 ( 
.A1(n_1316),
.A2(n_1335),
.A3(n_1332),
.B(n_1315),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1299),
.A2(n_118),
.B(n_115),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1366),
.B(n_69),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1317),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1363),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1329),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1380),
.A2(n_123),
.B(n_119),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1333),
.A2(n_127),
.B(n_124),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1271),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1349),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1356),
.A2(n_130),
.B(n_129),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1362),
.B(n_71),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1362),
.B(n_73),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1284),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1339),
.A2(n_132),
.B(n_131),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1367),
.B(n_73),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1368),
.B(n_74),
.Y(n_1474)
);

CKINVDCx8_ASAP7_75t_R g1475 ( 
.A(n_1326),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1350),
.A2(n_1370),
.B(n_1255),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1431),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1475),
.A2(n_1326),
.B1(n_1323),
.B2(n_1250),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1402),
.B(n_1295),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1413),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1458),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_SL g1482 ( 
.A1(n_1450),
.A2(n_1385),
.B(n_1272),
.C(n_1331),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1405),
.A2(n_1369),
.B(n_1347),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1411),
.A2(n_1334),
.B1(n_1288),
.B2(n_1248),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1412),
.B(n_1433),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1416),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1401),
.B(n_1295),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1443),
.Y(n_1488)
);

NAND2x1p5_ASAP7_75t_L g1489 ( 
.A(n_1412),
.B(n_1271),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1451),
.A2(n_1410),
.B(n_1397),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1414),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1432),
.A2(n_1259),
.B(n_1251),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1457),
.Y(n_1493)
);

INVx3_ASAP7_75t_SL g1494 ( 
.A(n_1392),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1458),
.B(n_1336),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1437),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1458),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1446),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1465),
.A2(n_1322),
.B(n_1269),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1446),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1463),
.B(n_1318),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1434),
.A2(n_1294),
.B1(n_1428),
.B2(n_1408),
.C(n_1404),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1420),
.A2(n_1297),
.B(n_1356),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1456),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1454),
.A2(n_1328),
.B1(n_1377),
.B2(n_1327),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_1433),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1476),
.A2(n_1382),
.B(n_1354),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1390),
.A2(n_1352),
.B(n_1328),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1440),
.A2(n_1307),
.B(n_1348),
.C(n_1321),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1456),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1472),
.A2(n_1259),
.B(n_1251),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1421),
.A2(n_1259),
.B(n_1251),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1418),
.A2(n_1381),
.B1(n_1348),
.B2(n_1307),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1424),
.A2(n_1247),
.B(n_1375),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1444),
.A2(n_1383),
.B(n_1360),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1469),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1403),
.A2(n_1360),
.B1(n_1327),
.B2(n_1321),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1419),
.Y(n_1519)
);

NAND2x1_ASAP7_75t_L g1520 ( 
.A(n_1399),
.B(n_1247),
.Y(n_1520)
);

AO21x2_ASAP7_75t_L g1521 ( 
.A1(n_1453),
.A2(n_1383),
.B(n_1337),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1394),
.A2(n_1375),
.B(n_1343),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1518),
.A2(n_1427),
.B1(n_1462),
.B2(n_1393),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1519),
.B(n_1395),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1480),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1492),
.A2(n_1388),
.B(n_1430),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1479),
.B(n_1486),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1484),
.A2(n_1449),
.B1(n_1470),
.B2(n_1467),
.Y(n_1529)
);

NAND2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1494),
.B(n_1351),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1490),
.A2(n_1448),
.B(n_1435),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1506),
.A2(n_1388),
.B1(n_1417),
.B2(n_1414),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1495),
.B(n_1406),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1507),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1507),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1520),
.A2(n_1422),
.B(n_1455),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_SL g1537 ( 
.A(n_1491),
.B(n_1243),
.C(n_1283),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1490),
.A2(n_1426),
.B(n_1398),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1491),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1495),
.B(n_1406),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1495),
.B(n_1446),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1508),
.A2(n_1389),
.B(n_1464),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1503),
.A2(n_1452),
.B1(n_1474),
.B2(n_1436),
.C(n_1423),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1481),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1508),
.A2(n_1459),
.B(n_1468),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1481),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1518),
.A2(n_1391),
.B1(n_1473),
.B2(n_1460),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1507),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1406),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1497),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1514),
.A2(n_1447),
.B1(n_1429),
.B2(n_1409),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1514),
.A2(n_1415),
.B1(n_1445),
.B2(n_1407),
.Y(n_1552)
);

BUFx8_ASAP7_75t_L g1553 ( 
.A(n_1477),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1525),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1529),
.A2(n_1510),
.B1(n_1478),
.B2(n_1517),
.C(n_1511),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1528),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1546),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1553),
.A2(n_1506),
.B1(n_1521),
.B2(n_1505),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1551),
.A2(n_1506),
.B1(n_1494),
.B2(n_1496),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1527),
.A2(n_1482),
.B(n_1516),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1533),
.B(n_1493),
.Y(n_1561)
);

INVx6_ASAP7_75t_L g1562 ( 
.A(n_1553),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1553),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1541),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1532),
.A2(n_1487),
.B(n_1504),
.C(n_1519),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1533),
.B(n_1540),
.Y(n_1566)
);

CKINVDCx16_ASAP7_75t_R g1567 ( 
.A(n_1539),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1502),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1543),
.A2(n_1547),
.B1(n_1523),
.B2(n_1530),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1530),
.A2(n_1487),
.B1(n_1521),
.B2(n_1500),
.Y(n_1570)
);

OAI211xp5_ASAP7_75t_L g1571 ( 
.A1(n_1537),
.A2(n_1482),
.B(n_1292),
.C(n_1519),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1552),
.A2(n_1516),
.B1(n_1502),
.B2(n_1498),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1534),
.A2(n_1485),
.B1(n_1489),
.B2(n_1516),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1485),
.Y(n_1574)
);

AOI33xp33_ASAP7_75t_L g1575 ( 
.A1(n_1541),
.A2(n_1466),
.A3(n_1342),
.B1(n_1357),
.B2(n_1498),
.B3(n_1501),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1541),
.Y(n_1576)
);

AOI222xp33_ASAP7_75t_L g1577 ( 
.A1(n_1539),
.A2(n_1501),
.B1(n_1471),
.B2(n_1442),
.C1(n_1438),
.C2(n_1281),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1535),
.B(n_1396),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1542),
.A2(n_1531),
.B(n_1538),
.Y(n_1579)
);

OAI21xp33_ASAP7_75t_L g1580 ( 
.A1(n_1549),
.A2(n_1489),
.B(n_1442),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1564),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1554),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1562),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1561),
.B(n_1549),
.Y(n_1584)
);

INVx3_ASAP7_75t_SL g1585 ( 
.A(n_1562),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1556),
.B(n_1544),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1587)
);

INVx5_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

INVx4_ASAP7_75t_R g1589 ( 
.A(n_1563),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1569),
.A2(n_1524),
.B1(n_1548),
.B2(n_1535),
.C(n_1545),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1566),
.B(n_1544),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1557),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1576),
.B(n_1564),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1578),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1564),
.B(n_1546),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1576),
.B(n_1546),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1573),
.B(n_1550),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1574),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1572),
.B(n_1550),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1579),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1589),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1583),
.A2(n_1559),
.B1(n_1558),
.B2(n_1570),
.Y(n_1603)
);

OAI211xp5_ASAP7_75t_L g1604 ( 
.A1(n_1590),
.A2(n_1565),
.B(n_1577),
.C(n_1571),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_R g1605 ( 
.A(n_1588),
.B(n_1567),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1581),
.B(n_1565),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1594),
.B(n_1555),
.C(n_1575),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1583),
.A2(n_1570),
.B1(n_1572),
.B2(n_1560),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1599),
.B(n_1580),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1591),
.B(n_1509),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1582),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1586),
.B(n_1575),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1597),
.A2(n_1548),
.B1(n_1425),
.B2(n_1438),
.C(n_1343),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1584),
.A2(n_1344),
.B1(n_1343),
.B2(n_1318),
.C(n_1303),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1610),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1612),
.B(n_1586),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1605),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1609),
.B(n_1591),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1611),
.B(n_1607),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1606),
.B(n_1587),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1606),
.B(n_1592),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1608),
.B(n_1600),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1581),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1603),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1604),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1613),
.B(n_1600),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1614),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1581),
.Y(n_1628)
);

AND2x4_ASAP7_75t_SL g1629 ( 
.A(n_1602),
.B(n_1596),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1611),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1612),
.B(n_1600),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1610),
.B(n_1593),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1632),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_1619),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1616),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1630),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1634),
.B(n_1625),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1636),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1638),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1633),
.B(n_1617),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1642),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1641),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1644),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1643),
.B(n_1625),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1643),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1644),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1645),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1648),
.B(n_1639),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1646),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1646),
.B(n_1639),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1647),
.B(n_1640),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1645),
.Y(n_1654)
);

XNOR2xp5_ASAP7_75t_L g1655 ( 
.A(n_1645),
.B(n_1627),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1650),
.B(n_1635),
.Y(n_1656)
);

NAND4xp25_ASAP7_75t_L g1657 ( 
.A(n_1649),
.B(n_1627),
.C(n_1622),
.D(n_1626),
.Y(n_1657)
);

NAND5xp2_ASAP7_75t_L g1658 ( 
.A(n_1652),
.B(n_1400),
.C(n_1623),
.D(n_1585),
.E(n_1621),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1649),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1655),
.B(n_1588),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1654),
.A2(n_1615),
.B1(n_1631),
.B2(n_1633),
.C(n_1628),
.Y(n_1661)
);

NAND4xp25_ASAP7_75t_L g1662 ( 
.A(n_1653),
.B(n_1628),
.C(n_1585),
.D(n_1620),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1615),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1649),
.B(n_1628),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1655),
.A2(n_1629),
.B(n_1588),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1655),
.A2(n_1629),
.B(n_1588),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1650),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1659),
.A2(n_1588),
.B1(n_1601),
.B2(n_1637),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1667),
.A2(n_1637),
.B1(n_1601),
.B2(n_1303),
.C(n_1595),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1664),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1670)
);

AOI222xp33_ASAP7_75t_L g1671 ( 
.A1(n_1663),
.A2(n_1596),
.B1(n_1320),
.B2(n_1336),
.C1(n_1318),
.C2(n_1344),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1660),
.A2(n_1374),
.B(n_1371),
.C(n_78),
.Y(n_1672)
);

AOI322xp5_ASAP7_75t_L g1673 ( 
.A1(n_1656),
.A2(n_1336),
.A3(n_1344),
.B1(n_79),
.B2(n_81),
.C1(n_82),
.C2(n_83),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1657),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1662),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1658),
.B(n_76),
.C(n_77),
.Y(n_1676)
);

OAI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1665),
.A2(n_1536),
.B(n_1276),
.C(n_1286),
.Y(n_1677)
);

NOR4xp75_ASAP7_75t_SL g1678 ( 
.A(n_1666),
.B(n_1661),
.C(n_83),
.D(n_77),
.Y(n_1678)
);

AOI222xp33_ASAP7_75t_L g1679 ( 
.A1(n_1667),
.A2(n_1304),
.B1(n_1308),
.B2(n_1310),
.C1(n_1313),
.C2(n_1387),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_SL g1680 ( 
.A(n_1659),
.B(n_81),
.C(n_84),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1659),
.A2(n_1276),
.B(n_1275),
.Y(n_1681)
);

XOR2x2_ASAP7_75t_L g1682 ( 
.A(n_1667),
.B(n_84),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_SL g1683 ( 
.A(n_1659),
.B(n_85),
.C(n_86),
.Y(n_1683)
);

AOI322xp5_ASAP7_75t_L g1684 ( 
.A1(n_1674),
.A2(n_86),
.A3(n_88),
.B1(n_89),
.B2(n_90),
.C1(n_91),
.C2(n_93),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_R g1685 ( 
.A(n_1680),
.B(n_88),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1675),
.A2(n_1668),
.B1(n_1676),
.B2(n_1669),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1683),
.Y(n_1687)
);

NOR5xp2_ASAP7_75t_L g1688 ( 
.A(n_1670),
.B(n_1678),
.C(n_1672),
.D(n_1677),
.E(n_1682),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1673),
.B(n_89),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1679),
.Y(n_1690)
);

OAI322xp33_ASAP7_75t_L g1691 ( 
.A1(n_1681),
.A2(n_1275),
.A3(n_1286),
.B1(n_93),
.B2(n_94),
.C1(n_95),
.C2(n_96),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1671),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1675),
.A2(n_1579),
.B1(n_1509),
.B2(n_1308),
.Y(n_1693)
);

OAI322xp33_ASAP7_75t_L g1694 ( 
.A1(n_1675),
.A2(n_90),
.A3(n_91),
.B1(n_95),
.B2(n_96),
.C1(n_97),
.C2(n_98),
.Y(n_1694)
);

CKINVDCx20_ASAP7_75t_R g1695 ( 
.A(n_1676),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_SL g1696 ( 
.A1(n_1675),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_1696)
);

AOI222xp33_ASAP7_75t_L g1697 ( 
.A1(n_1674),
.A2(n_1304),
.B1(n_1308),
.B2(n_1310),
.C1(n_1313),
.C2(n_104),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1675),
.Y(n_1698)
);

OA22x2_ASAP7_75t_L g1699 ( 
.A1(n_1675),
.A2(n_1531),
.B1(n_102),
.B2(n_100),
.Y(n_1699)
);

NOR2xp67_ASAP7_75t_L g1700 ( 
.A(n_1698),
.B(n_101),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1687),
.B(n_1304),
.Y(n_1701)
);

NAND4xp75_ASAP7_75t_L g1702 ( 
.A(n_1689),
.B(n_101),
.C(n_102),
.D(n_103),
.Y(n_1702)
);

NOR3xp33_ASAP7_75t_L g1703 ( 
.A(n_1694),
.B(n_104),
.C(n_106),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1695),
.B(n_106),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1699),
.Y(n_1705)
);

NOR2xp67_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_134),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1685),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1684),
.B(n_1579),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1696),
.A2(n_1445),
.B(n_1313),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1697),
.B(n_1396),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1690),
.A2(n_1310),
.B1(n_1499),
.B2(n_1483),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1692),
.B(n_1441),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1688),
.B(n_1693),
.C(n_1691),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1698),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_L g1715 ( 
.A(n_1694),
.B(n_135),
.C(n_140),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1698),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1698),
.Y(n_1717)
);

NOR4xp25_ASAP7_75t_L g1718 ( 
.A(n_1714),
.B(n_141),
.C(n_153),
.D(n_154),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1704),
.B(n_1375),
.Y(n_1719)
);

NOR4xp25_ASAP7_75t_L g1720 ( 
.A(n_1717),
.B(n_155),
.C(n_156),
.D(n_158),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1700),
.Y(n_1721)
);

NAND4xp25_ASAP7_75t_L g1722 ( 
.A(n_1703),
.B(n_160),
.C(n_162),
.D(n_163),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1705),
.A2(n_1499),
.B1(n_1483),
.B2(n_1538),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1713),
.A2(n_1396),
.B1(n_1439),
.B2(n_170),
.C(n_171),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1707),
.Y(n_1726)
);

NAND4xp75_ASAP7_75t_L g1727 ( 
.A(n_1706),
.B(n_164),
.C(n_166),
.D(n_172),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1702),
.B(n_174),
.Y(n_1728)
);

OAI211xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1715),
.A2(n_175),
.B(n_177),
.C(n_179),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1701),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1708),
.A2(n_1512),
.B1(n_1515),
.B2(n_1522),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1723),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1726),
.A2(n_1710),
.B1(n_1712),
.B2(n_1711),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1721),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1730),
.B(n_1712),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1728),
.B(n_1709),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1722),
.B(n_182),
.C(n_186),
.D(n_191),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1729),
.A2(n_1512),
.B(n_1515),
.C(n_1513),
.Y(n_1739)
);

NAND4xp25_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_192),
.C(n_197),
.D(n_198),
.Y(n_1740)
);

NOR3xp33_ASAP7_75t_SL g1741 ( 
.A(n_1727),
.B(n_200),
.C(n_204),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1732),
.A2(n_1720),
.B(n_1718),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1735),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1736),
.B(n_1731),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_SL g1745 ( 
.A(n_1734),
.B(n_1724),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1738),
.A2(n_1513),
.B1(n_1522),
.B2(n_209),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1733),
.B(n_205),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1741),
.B(n_207),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1739),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1743),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1748),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1742),
.A2(n_1737),
.B(n_1740),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1744),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1750),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1753),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1751),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1754),
.A2(n_1752),
.B(n_1747),
.Y(n_1757)
);

NAND2x1_ASAP7_75t_SL g1758 ( 
.A(n_1755),
.B(n_1745),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1758),
.Y(n_1759)
);

OAI321xp33_ASAP7_75t_L g1760 ( 
.A1(n_1757),
.A2(n_1749),
.A3(n_1756),
.B1(n_1746),
.B2(n_217),
.C(n_222),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1759),
.A2(n_1756),
.B1(n_1760),
.B2(n_215),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1759),
.A2(n_213),
.B1(n_214),
.B2(n_225),
.Y(n_1762)
);

AOI322xp5_ASAP7_75t_L g1763 ( 
.A1(n_1759),
.A2(n_226),
.A3(n_227),
.B1(n_228),
.B2(n_229),
.C1(n_230),
.C2(n_233),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1761),
.A2(n_234),
.B1(n_235),
.B2(n_238),
.C(n_239),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1762),
.B(n_1763),
.C(n_241),
.Y(n_1765)
);


endmodule