module fake_jpeg_10355_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_15),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_7),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_28),
.B1(n_16),
.B2(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_62),
.B1(n_28),
.B2(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_56),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_24),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_38),
.CON(n_65),
.SN(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_67),
.B(n_83),
.C(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_80),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_40),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_72),
.Y(n_118)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_87),
.Y(n_98)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_86),
.B1(n_20),
.B2(n_23),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_41),
.B(n_33),
.C(n_17),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_36),
.A3(n_39),
.B1(n_33),
.B2(n_18),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_89),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_33),
.B1(n_19),
.B2(n_23),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_36),
.C(n_35),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_30),
.B1(n_27),
.B2(n_32),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_100),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_84),
.B1(n_85),
.B2(n_66),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_89),
.B1(n_71),
.B2(n_70),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_55),
.B1(n_44),
.B2(n_21),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_97),
.A2(n_117),
.B1(n_120),
.B2(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_51),
.B1(n_44),
.B2(n_21),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_71),
.B1(n_89),
.B2(n_80),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_27),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_114),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_115),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_73),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_74),
.A2(n_20),
.B1(n_25),
.B2(n_17),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_69),
.C(n_77),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_101),
.C(n_29),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_123),
.A2(n_145),
.B(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_124),
.B(n_126),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_125),
.B(n_9),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_107),
.B1(n_103),
.B2(n_102),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_119),
.B1(n_22),
.B2(n_29),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_77),
.B(n_82),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_139),
.B(n_140),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_82),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_141),
.B(n_29),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_142),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_149),
.B1(n_150),
.B2(n_113),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_13),
.B(n_12),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_121),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_93),
.B(n_22),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_88),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_27),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_88),
.B1(n_76),
.B2(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_1),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_160),
.Y(n_188)
);

OAI211xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_30),
.B(n_22),
.C(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_181),
.Y(n_189)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_22),
.B1(n_95),
.B2(n_100),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_149),
.B1(n_150),
.B2(n_130),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_99),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_169),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_123),
.B1(n_131),
.B2(n_130),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

XOR2x2_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_101),
.Y(n_161)
);

OA21x2_ASAP7_75t_SL g201 ( 
.A1(n_161),
.A2(n_184),
.B(n_126),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_22),
.B(n_29),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_172),
.B1(n_136),
.B2(n_129),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_108),
.B1(n_115),
.B2(n_101),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_1),
.C(n_2),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_183),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_10),
.A3(n_13),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_14),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_137),
.B1(n_145),
.B2(n_144),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_198),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_190),
.A2(n_196),
.B(n_197),
.C(n_2),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_176),
.B1(n_156),
.B2(n_183),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_125),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_200),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_155),
.B(n_135),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_167),
.B(n_154),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_211),
.B(n_163),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_127),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_158),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_167),
.CI(n_169),
.CON(n_213),
.SN(n_213)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_230),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_157),
.C(n_210),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_175),
.B(n_179),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_229),
.B(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_174),
.C(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_166),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_182),
.B(n_166),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_219),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_223),
.Y(n_251)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_232),
.B1(n_196),
.B2(n_225),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_231),
.C(n_235),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_156),
.B(n_155),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_188),
.A2(n_206),
.B(n_189),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_138),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_10),
.B(n_12),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_11),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_242),
.B(n_243),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_185),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_218),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_227),
.B1(n_205),
.B2(n_198),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_232),
.B1(n_231),
.B2(n_213),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_187),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_224),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_255),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_251),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_247),
.B1(n_246),
.B2(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_244),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_250),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_232),
.B1(n_222),
.B2(n_193),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_269),
.B1(n_252),
.B2(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_211),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_202),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_232),
.B1(n_193),
.B2(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_245),
.B1(n_251),
.B2(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_266),
.B1(n_269),
.B2(n_249),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_277),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_250),
.B(n_240),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_274),
.B(n_258),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_226),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_195),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_195),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_292),
.B(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_264),
.C(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_288),
.C(n_262),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_263),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_12),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_280),
.C(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_4),
.B1(n_6),
.B2(n_11),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_259),
.B(n_260),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_186),
.B(n_212),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_297),
.C(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_216),
.C(n_228),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_4),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_302),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_13),
.C(n_11),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_2),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_306),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_293),
.B(n_288),
.Y(n_308)
);

OAI31xp33_ASAP7_75t_SL g311 ( 
.A1(n_308),
.A2(n_303),
.A3(n_287),
.B(n_291),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_310),
.B(n_309),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_304),
.C(n_3),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_3),
.B(n_304),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_3),
.Y(n_315)
);


endmodule