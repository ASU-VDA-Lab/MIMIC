module fake_jpeg_11793_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_57),
.B(n_62),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_58),
.B(n_85),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_64),
.B(n_67),
.Y(n_160)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_68),
.B(n_71),
.Y(n_162)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_72),
.Y(n_153)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_86),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_84),
.B(n_88),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_18),
.B(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_0),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_37),
.Y(n_90)
);

NAND2xp67_ASAP7_75t_SL g158 ( 
.A(n_90),
.B(n_50),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_54),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_119),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_20),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_103),
.B(n_113),
.Y(n_181)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_20),
.B(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_107),
.B(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_25),
.B(n_15),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_25),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_109),
.B(n_3),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_48),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_34),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_114),
.B(n_116),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_48),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_121),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_45),
.B1(n_42),
.B2(n_49),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_122),
.A2(n_139),
.B(n_140),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_61),
.A2(n_42),
.B1(n_45),
.B2(n_49),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_126),
.A2(n_154),
.B1(n_177),
.B2(n_180),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_45),
.B1(n_42),
.B2(n_46),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_72),
.A2(n_22),
.B1(n_53),
.B2(n_46),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_72),
.A2(n_21),
.B1(n_53),
.B2(n_31),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_143),
.A2(n_150),
.B1(n_161),
.B2(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_148),
.B(n_155),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_69),
.A2(n_21),
.B1(n_31),
.B2(n_27),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_56),
.B1(n_27),
.B2(n_22),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_70),
.B(n_55),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_158),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_78),
.B(n_28),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_159),
.B(n_163),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_50),
.B1(n_41),
.B2(n_35),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_73),
.B(n_41),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_81),
.A2(n_56),
.B1(n_35),
.B2(n_28),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_101),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_173),
.B(n_186),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_79),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_63),
.A2(n_26),
.B1(n_1),
.B2(n_3),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_102),
.B(n_0),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_182),
.B(n_188),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_194),
.C(n_196),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_89),
.B(n_3),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_3),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_110),
.B(n_5),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_192),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_112),
.B(n_7),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_79),
.B(n_7),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_197),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_80),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_196),
.A2(n_199),
.B1(n_201),
.B2(n_177),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_80),
.B(n_9),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_75),
.A2(n_11),
.B1(n_12),
.B2(n_105),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_94),
.A2(n_11),
.B1(n_12),
.B2(n_119),
.Y(n_201)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_125),
.B(n_101),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_202),
.A2(n_213),
.B(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_205),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_124),
.B(n_11),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_206),
.B(n_216),
.Y(n_279)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_208),
.B(n_217),
.Y(n_269)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_209),
.Y(n_301)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_210),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_211),
.Y(n_299)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_212),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_153),
.A2(n_59),
.B(n_94),
.C(n_120),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_146),
.B(n_92),
.Y(n_215)
);

NAND2x1p5_ASAP7_75t_L g294 ( 
.A(n_215),
.B(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_142),
.B(n_117),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_149),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_138),
.B(n_82),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_262),
.C(n_264),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_220),
.A2(n_132),
.B1(n_213),
.B2(n_219),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_147),
.B(n_106),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_239),
.Y(n_280)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_115),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_223),
.B(n_226),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_128),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_118),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_228),
.B(n_234),
.Y(n_289)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_126),
.A2(n_121),
.B1(n_200),
.B2(n_154),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_233),
.A2(n_237),
.B1(n_261),
.B2(n_263),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_129),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_164),
.A2(n_184),
.B1(n_167),
.B2(n_131),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_152),
.B(n_145),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_187),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_241),
.B(n_246),
.Y(n_302)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_242),
.B(n_243),
.Y(n_303)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_127),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_244),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_164),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_134),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_252),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_127),
.B(n_135),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_123),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_123),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_156),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_256),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_257),
.A2(n_260),
.B1(n_266),
.B2(n_236),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_129),
.A2(n_201),
.B(n_150),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_267),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_122),
.A2(n_139),
.B(n_136),
.C(n_174),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_167),
.A2(n_131),
.B1(n_171),
.B2(n_176),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_136),
.B(n_144),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_171),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_157),
.B(n_156),
.C(n_191),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_144),
.B(n_133),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_166),
.B1(n_176),
.B2(n_157),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_274),
.B1(n_291),
.B2(n_295),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_249),
.A2(n_166),
.B1(n_179),
.B2(n_191),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_141),
.B1(n_174),
.B2(n_179),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g358 ( 
.A1(n_278),
.A2(n_288),
.B1(n_294),
.B2(n_270),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_216),
.A2(n_132),
.B1(n_221),
.B2(n_245),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_224),
.C(n_239),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_293),
.C(n_297),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_206),
.B(n_218),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_246),
.A2(n_223),
.B1(n_230),
.B2(n_268),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_202),
.B(n_203),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_230),
.A2(n_229),
.B1(n_257),
.B2(n_225),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_305),
.A2(n_309),
.B1(n_310),
.B2(n_295),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_265),
.A2(n_235),
.B1(n_259),
.B2(n_264),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_219),
.A2(n_215),
.B1(n_204),
.B2(n_263),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_202),
.B(n_215),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_317),
.C(n_319),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_215),
.A2(n_212),
.B1(n_232),
.B2(n_231),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_313),
.A2(n_298),
.B1(n_285),
.B2(n_277),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_252),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_209),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_234),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_320),
.B(n_324),
.Y(n_372)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_305),
.A2(n_247),
.B1(n_238),
.B2(n_254),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_323),
.A2(n_355),
.B1(n_299),
.B2(n_275),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_205),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_242),
.C(n_227),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_340),
.C(n_299),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_243),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_266),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_343),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_300),
.A2(n_210),
.B(n_250),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_331),
.A2(n_334),
.B(n_316),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_279),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_315),
.A2(n_260),
.B(n_207),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_293),
.B(n_214),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_336),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_272),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_318),
.A2(n_222),
.B1(n_240),
.B2(n_274),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_346),
.B1(n_349),
.B2(n_356),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_297),
.C(n_292),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_289),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_341),
.Y(n_359)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_310),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_345),
.A2(n_352),
.B(n_358),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_291),
.A2(n_311),
.B1(n_307),
.B2(n_302),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_279),
.B(n_302),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_348),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_282),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_282),
.A2(n_273),
.B1(n_317),
.B2(n_288),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_286),
.B(n_315),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_354),
.Y(n_386)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_300),
.A2(n_294),
.B(n_278),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_284),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_353),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_308),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_278),
.A2(n_294),
.B1(n_290),
.B2(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_301),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_362),
.C(n_376),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_355),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_378),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_345),
.A2(n_278),
.B1(n_271),
.B2(n_276),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_368),
.A2(n_382),
.B1(n_384),
.B2(n_323),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_371),
.A2(n_329),
.B(n_326),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_316),
.C(n_270),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_352),
.A2(n_278),
.B(n_331),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_377),
.A2(n_343),
.B(n_334),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_327),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_325),
.C(n_347),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_329),
.C(n_358),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_330),
.A2(n_349),
.B1(n_346),
.B2(n_356),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_332),
.B1(n_358),
.B2(n_333),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_354),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_328),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_386),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_393),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_359),
.B(n_338),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_391),
.B(n_403),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_386),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_394),
.A2(n_396),
.B(n_412),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_377),
.A2(n_333),
.B(n_343),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_395),
.A2(n_414),
.B(n_415),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_398),
.A2(n_413),
.B1(n_389),
.B2(n_370),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_400),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_367),
.A2(n_358),
.B1(n_325),
.B2(n_322),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_401),
.A2(n_407),
.B1(n_375),
.B2(n_376),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_411),
.C(n_366),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_359),
.B(n_351),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_387),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_408),
.Y(n_423)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_378),
.A2(n_342),
.B1(n_357),
.B2(n_344),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_361),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_361),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_410),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_383),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_381),
.C(n_362),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_321),
.B(n_371),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_384),
.B1(n_375),
.B2(n_368),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_321),
.B(n_364),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_374),
.A2(n_321),
.B(n_373),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_373),
.Y(n_416)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_417),
.A2(n_418),
.B1(n_425),
.B2(n_430),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_385),
.B1(n_364),
.B2(n_372),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_383),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_439),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_433),
.C(n_397),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_399),
.A2(n_372),
.B1(n_366),
.B2(n_363),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_390),
.B1(n_407),
.B2(n_410),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_401),
.A2(n_389),
.B1(n_370),
.B2(n_388),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_388),
.Y(n_431)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_379),
.C(n_365),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_379),
.Y(n_436)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_365),
.Y(n_437)
);

XOR2x1_ASAP7_75t_SL g444 ( 
.A(n_437),
.B(n_395),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_402),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_442),
.C(n_453),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_397),
.C(n_402),
.Y(n_442)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_396),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_446),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_416),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_394),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_457),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_394),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_434),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_452),
.A2(n_456),
.B1(n_432),
.B2(n_438),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_414),
.C(n_412),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_422),
.A2(n_423),
.B(n_404),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_454),
.B(n_455),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_414),
.C(n_412),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_429),
.A2(n_391),
.B1(n_403),
.B2(n_405),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_413),
.C(n_398),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_SL g461 ( 
.A(n_448),
.B(n_423),
.C(n_428),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_462),
.Y(n_477)
);

NAND4xp25_ASAP7_75t_SL g462 ( 
.A(n_444),
.B(n_437),
.C(n_428),
.D(n_436),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_458),
.Y(n_464)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_449),
.A2(n_420),
.B1(n_435),
.B2(n_438),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_466),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_434),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_472),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_445),
.C(n_451),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_471),
.A2(n_473),
.B1(n_459),
.B2(n_440),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_455),
.A2(n_432),
.B(n_420),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_485),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_441),
.C(n_442),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_476),
.B(n_478),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_443),
.C(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_457),
.B1(n_459),
.B2(n_453),
.Y(n_481)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_481),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_440),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_482),
.B(n_483),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_464),
.B(n_431),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_467),
.A2(n_392),
.B(n_425),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_477),
.B1(n_470),
.B2(n_484),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_488),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_474),
.A2(n_461),
.B1(n_462),
.B2(n_466),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_480),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_490),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_463),
.C(n_468),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_475),
.B(n_392),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_492),
.A2(n_478),
.B(n_469),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_486),
.A2(n_487),
.B(n_490),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_503),
.Y(n_506)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_498),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_463),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_499),
.B(n_500),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_493),
.B(n_406),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_424),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_502),
.A2(n_488),
.B1(n_495),
.B2(n_424),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_493),
.B(n_468),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_501),
.B(n_492),
.Y(n_505)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_505),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_497),
.B1(n_426),
.B2(n_398),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_502),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_510),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_511),
.A2(n_506),
.B(n_508),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_512),
.A2(n_506),
.B1(n_426),
.B2(n_413),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_514),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_515),
.B(n_513),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_447),
.Y(n_517)
);


endmodule