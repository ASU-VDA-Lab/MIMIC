module fake_jpeg_28864_n_446 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_446);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_53),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_22),
.B(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_12),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_8),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_83),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_85),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_88),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_26),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_21),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_104),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_135),
.Y(n_171)
);

BUFx4f_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_137),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g132 ( 
.A(n_70),
.Y(n_132)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_71),
.Y(n_137)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_166),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_73),
.B1(n_63),
.B2(n_79),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_174),
.B1(n_176),
.B2(n_87),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_109),
.A2(n_68),
.B(n_62),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_136),
.B1(n_108),
.B2(n_121),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_165),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_78),
.B1(n_58),
.B2(n_84),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_94),
.B1(n_124),
.B2(n_128),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_175),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_43),
.B1(n_28),
.B2(n_41),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_43),
.B1(n_28),
.B2(n_41),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_128),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_110),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_143),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_94),
.B1(n_124),
.B2(n_117),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_115),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_168),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_118),
.B(n_108),
.C(n_138),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_147),
.B(n_131),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_158),
.Y(n_206)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_205),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_213),
.Y(n_232)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_214),
.B1(n_220),
.B2(n_224),
.Y(n_236)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_172),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_118),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_223),
.Y(n_233)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_163),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_225),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_101),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_186),
.C(n_180),
.Y(n_242)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_219),
.Y(n_244)
);

INVx3_ASAP7_75t_SL g221 ( 
.A(n_200),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_187),
.B1(n_183),
.B2(n_200),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_227),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_178),
.B(n_23),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_149),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_29),
.B(n_37),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_201),
.B(n_186),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_153),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_229),
.Y(n_251)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_221),
.A2(n_180),
.B1(n_177),
.B2(n_166),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_235),
.A2(n_240),
.B(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_239),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_184),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_201),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_248),
.C(n_219),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_245),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_108),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_26),
.C(n_13),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_192),
.C(n_181),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_44),
.C(n_23),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_30),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_181),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_214),
.A2(n_177),
.B1(n_165),
.B2(n_162),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_208),
.B1(n_198),
.B2(n_197),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_263),
.Y(n_290)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_226),
.B1(n_215),
.B2(n_220),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_258),
.A2(n_254),
.B1(n_197),
.B2(n_154),
.Y(n_302)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_251),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_261),
.Y(n_292)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_225),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_264),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_211),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_273),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_266),
.B(n_216),
.Y(n_304)
);

AOI22x1_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_224),
.B1(n_215),
.B2(n_229),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_268),
.A2(n_140),
.B1(n_146),
.B2(n_139),
.Y(n_310)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_281),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_233),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_233),
.B(n_228),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_244),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_224),
.B(n_221),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_277),
.A2(n_278),
.B(n_136),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_241),
.A2(n_224),
.B(n_167),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_255),
.B1(n_254),
.B2(n_230),
.Y(n_287)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_229),
.B(n_216),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_284),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_192),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_208),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_152),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_236),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_286),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_270),
.B1(n_269),
.B2(n_271),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_289),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_242),
.Y(n_296)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_245),
.B(n_230),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_310),
.B(n_280),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_253),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_302),
.A2(n_314),
.B1(n_189),
.B2(n_175),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_267),
.C(n_285),
.Y(n_323)
);

XOR2x1_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_277),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_284),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_260),
.A2(n_173),
.B(n_145),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_275),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_189),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_279),
.A2(n_44),
.B1(n_33),
.B2(n_161),
.Y(n_314)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_316),
.A2(n_319),
.B1(n_307),
.B2(n_310),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_290),
.B(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_328),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_326),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_304),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_299),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_274),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_301),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_329),
.B(n_305),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_301),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_288),
.C(n_303),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_334),
.C(n_336),
.Y(n_342)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_259),
.B(n_257),
.Y(n_333)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_293),
.C(n_298),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_281),
.C(n_258),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_292),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_275),
.C(n_272),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_337),
.A2(n_298),
.B1(n_293),
.B2(n_313),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_283),
.C(n_257),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_308),
.C(n_313),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_350),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_332),
.A2(n_302),
.B1(n_292),
.B2(n_294),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_343),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_320),
.B(n_306),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_339),
.A2(n_334),
.B1(n_319),
.B2(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_315),
.Y(n_348)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_309),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_102),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_321),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_355),
.A2(n_359),
.B1(n_145),
.B2(n_205),
.Y(n_370)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_360),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_311),
.C(n_283),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_115),
.C(n_57),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_318),
.A2(n_324),
.B1(n_329),
.B2(n_326),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_311),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_362),
.B(n_49),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_363),
.B(n_367),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_351),
.A2(n_336),
.B(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_351),
.A2(n_282),
.B(n_262),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_SL g368 ( 
.A1(n_349),
.A2(n_282),
.B(n_262),
.C(n_207),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_370),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_207),
.B(n_205),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_358),
.Y(n_385)
);

AO221x1_ASAP7_75t_L g372 ( 
.A1(n_346),
.A2(n_33),
.B1(n_37),
.B2(n_29),
.C(n_4),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_382),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_102),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_103),
.C(n_96),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_344),
.C(n_350),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_352),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_378),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_355),
.A2(n_46),
.B1(n_41),
.B2(n_103),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_381),
.B(n_353),
.Y(n_387)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_354),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_391),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_392),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_364),
.A2(n_342),
.B(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_395),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_344),
.C(n_46),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_95),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_373),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_14),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_96),
.C(n_77),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_380),
.C(n_376),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_368),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_389),
.A2(n_383),
.B(n_379),
.Y(n_400)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_400),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_403),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_407),
.Y(n_414)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_384),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_408),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_390),
.A2(n_376),
.B(n_375),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_396),
.B(n_369),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_393),
.B(n_369),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_387),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_393),
.C(n_394),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_415),
.Y(n_424)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_14),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_368),
.C(n_50),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_420),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_399),
.A2(n_368),
.B1(n_30),
.B2(n_76),
.Y(n_418)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_74),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_17),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_413),
.A2(n_405),
.B(n_402),
.Y(n_422)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_422),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_421),
.A2(n_17),
.B(n_16),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_17),
.B(n_15),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_7),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_427),
.Y(n_433)
);

AOI322xp5_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_419),
.A3(n_414),
.B1(n_417),
.B2(n_151),
.C1(n_95),
.C2(n_48),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_429),
.A2(n_424),
.B(n_425),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_432),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_428),
.A2(n_430),
.B1(n_427),
.B2(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_56),
.C(n_151),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_422),
.A2(n_114),
.B(n_156),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_436),
.B(n_156),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_438),
.C(n_15),
.Y(n_442)
);

AOI322xp5_ASAP7_75t_L g439 ( 
.A1(n_435),
.A2(n_138),
.A3(n_64),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_14),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_433),
.B(n_3),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_441),
.B(n_442),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_440),
.C(n_15),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_0),
.B(n_1),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_0),
.B(n_1),
.Y(n_446)
);


endmodule