module fake_netlist_6_104_n_44 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_8, n_44);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_8;

output n_44;

wire n_41;
wire n_16;
wire n_34;
wire n_42;
wire n_9;
wire n_10;
wire n_21;
wire n_18;
wire n_24;
wire n_37;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_38;
wire n_39;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_30;
wire n_43;
wire n_19;
wire n_29;
wire n_31;
wire n_25;
wire n_40;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx5p33_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR3xp33_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

AND2x6_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

AND2x4_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_2),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_14),
.B1(n_15),
.B2(n_13),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_20),
.Y(n_28)
);

OAI321xp33_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_23),
.A3(n_21),
.B1(n_22),
.B2(n_18),
.C(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI31xp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_16),
.A3(n_18),
.B(n_19),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_9),
.B1(n_18),
.B2(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_29),
.B(n_31),
.Y(n_37)
);

AOI221xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_19),
.B1(n_32),
.B2(n_4),
.C(n_8),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_33),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_32),
.A3(n_34),
.B1(n_41),
.B2(n_42),
.C1(n_38),
.C2(n_40),
.Y(n_44)
);


endmodule