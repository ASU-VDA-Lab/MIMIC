module fake_ariane_1802_n_3064 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_381, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_382, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_3064);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_3064;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_416;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_3063;
wire n_813;
wire n_1985;
wire n_419;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_559;
wire n_2663;
wire n_495;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_2650;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2391;
wire n_2332;
wire n_611;
wire n_2060;
wire n_1295;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_533;
wire n_3049;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_2739;
wire n_512;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_461;
wire n_1416;
wire n_2909;
wire n_490;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2326;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_444;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2926;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_2970;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_418;
wire n_2185;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_436;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_2628;
wire n_619;
wire n_967;
wire n_437;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_2598;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_489;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_397;
wire n_2467;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_3052;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_404;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_2649;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_441;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_637;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_2841;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_481;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_502;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_3022;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_699;
wire n_727;
wire n_590;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1614;
wire n_1162;
wire n_1377;
wire n_536;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_2853;
wire n_636;
wire n_427;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_390;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_451;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1975;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_403;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_1700;
wire n_862;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_1748;
wire n_873;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_2939;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_474;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_2785;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_2574;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1281;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1856;
wire n_463;
wire n_1524;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_3050;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_643;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_473;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2477;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_3043;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_640;
wire n_644;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_497;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_2343;
wire n_1048;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_2401;
wire n_2935;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_409;
wire n_2963;
wire n_519;
wire n_384;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_820;
wire n_1749;
wire n_1653;
wire n_872;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_395;
wire n_2648;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_580;
wire n_1579;
wire n_494;
wire n_2809;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_394;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_679;
wire n_3047;
wire n_1720;
wire n_663;
wire n_2409;
wire n_2966;
wire n_443;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_385;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_399;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_2967;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_2897;
wire n_816;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3038;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1409;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_488;
wire n_3018;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_459;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1983;
wire n_1273;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_448;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_450;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_1591;
wire n_664;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_2052;
wire n_2485;
wire n_1091;
wire n_1063;
wire n_537;
wire n_991;
wire n_2275;
wire n_2183;
wire n_2205;
wire n_389;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_457;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_412;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_447;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_796;
wire n_573;
wire n_2851;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_348),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_234),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_19),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_160),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_241),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_164),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_201),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_85),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_170),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_217),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_272),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_172),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_36),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_375),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_303),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_255),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_329),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_279),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_144),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_97),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_370),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_344),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_354),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_22),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_58),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_128),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_199),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_51),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_109),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_9),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_278),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_225),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_92),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_159),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_72),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_132),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_335),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_283),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_246),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_287),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_223),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_176),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_299),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_350),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_96),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_169),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_87),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_109),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_137),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_101),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_123),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_205),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_215),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_81),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_297),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_71),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_104),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_372),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_262),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_21),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_165),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_153),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_210),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_45),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_140),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_158),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_308),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_167),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_209),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_1),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_239),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_165),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_84),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_99),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_56),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_216),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_23),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_19),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_341),
.Y(n_469)
);

INVxp33_ASAP7_75t_R g470 ( 
.A(n_369),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_61),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_274),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_26),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_374),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_232),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_130),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_380),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_288),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_328),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_356),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_174),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_182),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_214),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_124),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_224),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_330),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_77),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_291),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_212),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_342),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_218),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_363),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_220),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_270),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_382),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_231),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_146),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_181),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_265),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_143),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_347),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_195),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_13),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_268),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_136),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_359),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_134),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_92),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_148),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_332),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_113),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_77),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_230),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_16),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_243),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_104),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_99),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_346),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_181),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_57),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_306),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_317),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_38),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_176),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_67),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_142),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_365),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_106),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_111),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_86),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_33),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_343),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_13),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_349),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_52),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_63),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_47),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_129),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_160),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_364),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_142),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_59),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_70),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_132),
.Y(n_545)
);

CKINVDCx14_ASAP7_75t_R g546 ( 
.A(n_21),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_353),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_158),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_295),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_75),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_95),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_37),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_254),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_357),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_233),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_340),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_100),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_89),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_251),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_352),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_47),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_244),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_164),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_54),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_207),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_286),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_377),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_337),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_197),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_138),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_381),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_76),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_61),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_373),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_257),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_22),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_138),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_68),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_137),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_39),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_69),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_170),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_242),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_376),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_260),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_321),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_339),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_249),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_143),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_83),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_309),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_338),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_345),
.Y(n_593)
);

INVxp33_ASAP7_75t_SL g594 ( 
.A(n_15),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_316),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_93),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_161),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_54),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_64),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_128),
.Y(n_600)
);

BUFx5_ASAP7_75t_L g601 ( 
.A(n_112),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_83),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_126),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_106),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_240),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_351),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_95),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_107),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_15),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_296),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_161),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_146),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_110),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_171),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_213),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_116),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_120),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_281),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_39),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_49),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_211),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_289),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_33),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_70),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_229),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_26),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_336),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_93),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_177),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_157),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_156),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_206),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_107),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_153),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_204),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_355),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_159),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_294),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_199),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_358),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_195),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_196),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_247),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_290),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_379),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_293),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_27),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_98),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_79),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_201),
.Y(n_650)
);

BUFx8_ASAP7_75t_SL g651 ( 
.A(n_63),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_42),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_171),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_320),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_64),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_94),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_252),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_238),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_79),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_361),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_202),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_127),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_25),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_8),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_67),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_185),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_245),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_136),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_177),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_58),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_75),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_111),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_124),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_118),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_100),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_227),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_6),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_334),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_118),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_187),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_98),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_144),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_27),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_101),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_154),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_277),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_300),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_97),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_52),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_601),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

INVxp33_ASAP7_75t_L g692 ( 
.A(n_661),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_526),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_529),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_601),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_601),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_601),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_601),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_601),
.Y(n_700)
);

INVxp67_ASAP7_75t_SL g701 ( 
.A(n_529),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_601),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_601),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_546),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_388),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_424),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_388),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_533),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_398),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_395),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_398),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_395),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_400),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_400),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_540),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_402),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_533),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_402),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_411),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_411),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_420),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_420),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_540),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_629),
.Y(n_724)
);

INVxp67_ASAP7_75t_SL g725 ( 
.A(n_602),
.Y(n_725)
);

INVxp33_ASAP7_75t_L g726 ( 
.A(n_651),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_448),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_622),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_448),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_622),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_408),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_454),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_602),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_454),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_476),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_476),
.Y(n_736)
);

INVxp33_ASAP7_75t_SL g737 ( 
.A(n_629),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_452),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_489),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_489),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_408),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_493),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_452),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_472),
.Y(n_744)
);

CKINVDCx14_ASAP7_75t_R g745 ( 
.A(n_475),
.Y(n_745)
);

INVxp33_ASAP7_75t_SL g746 ( 
.A(n_668),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_424),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_384),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_424),
.Y(n_750)
);

INVxp33_ASAP7_75t_SL g751 ( 
.A(n_389),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_689),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_387),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_385),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_385),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_689),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_414),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_493),
.B(n_0),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_414),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_421),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_422),
.Y(n_761)
);

INVxp33_ASAP7_75t_SL g762 ( 
.A(n_391),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_403),
.Y(n_763)
);

INVxp33_ASAP7_75t_SL g764 ( 
.A(n_392),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_422),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_431),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_431),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_434),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_434),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_435),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_435),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_424),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_438),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_424),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_438),
.Y(n_775)
);

INVxp33_ASAP7_75t_SL g776 ( 
.A(n_396),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_439),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_505),
.B(n_0),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_439),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_450),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_445),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_445),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_446),
.Y(n_783)
);

INVxp33_ASAP7_75t_L g784 ( 
.A(n_446),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_456),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_450),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_456),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_464),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_464),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_471),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_471),
.Y(n_791)
);

CKINVDCx16_ASAP7_75t_R g792 ( 
.A(n_518),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_450),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_505),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_405),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_403),
.Y(n_796)
);

CKINVDCx14_ASAP7_75t_R g797 ( 
.A(n_403),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_553),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_516),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_450),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_450),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_516),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_528),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_485),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_485),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_397),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_528),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_549),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_549),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_554),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_401),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_554),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_410),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_583),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_499),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_410),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_583),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_407),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_553),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_584),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_660),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_584),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_678),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_586),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_412),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_686),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_453),
.Y(n_827)
);

CKINVDCx16_ASAP7_75t_R g828 ( 
.A(n_518),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_586),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_780),
.Y(n_830)
);

OAI22x1_ASAP7_75t_SL g831 ( 
.A1(n_737),
.A2(n_488),
.B1(n_513),
.B2(n_455),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_738),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_706),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_753),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_780),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_705),
.B(n_386),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_706),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_738),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_780),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_691),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_813),
.B(n_462),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_813),
.B(n_462),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_690),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_695),
.B(n_591),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_710),
.B(n_390),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_738),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_816),
.B(n_543),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_747),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_745),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_747),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_750),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_750),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_772),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_784),
.B(n_518),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_772),
.Y(n_855)
);

BUFx12f_ASAP7_75t_L g856 ( 
.A(n_708),
.Y(n_856)
);

AND2x2_ASAP7_75t_SL g857 ( 
.A(n_758),
.B(n_386),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_778),
.A2(n_592),
.B(n_591),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_797),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_691),
.A2(n_635),
.B(n_592),
.Y(n_860)
);

OA21x2_ASAP7_75t_L g861 ( 
.A1(n_690),
.A2(n_645),
.B(n_635),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_738),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_738),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_786),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_786),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_743),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_792),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_753),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_696),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_816),
.B(n_543),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_793),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_793),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_705),
.B(n_597),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_751),
.B(n_645),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_746),
.A2(n_579),
.B1(n_580),
.B2(n_550),
.Y(n_875)
);

AND2x6_ASAP7_75t_L g876 ( 
.A(n_707),
.B(n_393),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_701),
.B(n_646),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_696),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_763),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_743),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_697),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_801),
.Y(n_882)
);

BUFx8_ASAP7_75t_SL g883 ( 
.A(n_748),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_743),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_708),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_801),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_725),
.B(n_534),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_697),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_733),
.B(n_534),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_741),
.B(n_597),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_743),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_806),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_760),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_743),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_698),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_698),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_699),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_699),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_700),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_763),
.B(n_796),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_707),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_710),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_700),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_702),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_774),
.B(n_646),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_702),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_703),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_703),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_796),
.B(n_553),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_709),
.B(n_393),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_709),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_811),
.Y(n_912)
);

INVx6_ASAP7_75t_L g913 ( 
.A(n_731),
.Y(n_913)
);

OA21x2_ASAP7_75t_L g914 ( 
.A1(n_711),
.A2(n_657),
.B(n_428),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_SL g915 ( 
.A1(n_818),
.A2(n_596),
.B1(n_616),
.B2(n_582),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_741),
.B(n_717),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_717),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_800),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_693),
.B(n_534),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_711),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_713),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_731),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_728),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_713),
.B(n_671),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_714),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_714),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_716),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_728),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_716),
.B(n_671),
.Y(n_929)
);

BUFx12f_ASAP7_75t_L g930 ( 
.A(n_730),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_718),
.Y(n_931)
);

CKINVDCx6p67_ASAP7_75t_R g932 ( 
.A(n_704),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_798),
.B(n_657),
.Y(n_933)
);

OAI22x1_ASAP7_75t_L g934 ( 
.A1(n_715),
.A2(n_482),
.B1(n_509),
.B2(n_417),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_718),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_694),
.B(n_805),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_719),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_719),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_720),
.Y(n_939)
);

AND2x4_ASAP7_75t_SL g940 ( 
.A(n_821),
.B(n_604),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_720),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_823),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_721),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_721),
.Y(n_944)
);

CKINVDCx6p67_ASAP7_75t_R g945 ( 
.A(n_828),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_722),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_722),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_827),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_727),
.B(n_404),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_727),
.Y(n_950)
);

INVxp33_ASAP7_75t_SL g951 ( 
.A(n_744),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_729),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_729),
.B(n_404),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_732),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_921),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_921),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_921),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_897),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_897),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_895),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_868),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_921),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_888),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_895),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_950),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_854),
.B(n_949),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_904),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_904),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_888),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_950),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_895),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_906),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_950),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_919),
.B(n_815),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_860),
.A2(n_734),
.B(n_732),
.Y(n_975)
);

OA21x2_ASAP7_75t_L g976 ( 
.A1(n_860),
.A2(n_735),
.B(n_734),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_861),
.A2(n_736),
.B(n_735),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_906),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_907),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_950),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_854),
.B(n_736),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_857),
.B(n_798),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_840),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_907),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_874),
.B(n_730),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_840),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_893),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_911),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_919),
.B(n_804),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_840),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_840),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_914),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_914),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_883),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_949),
.B(n_739),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_914),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_914),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_911),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_911),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_948),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_895),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_895),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_903),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_903),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_857),
.B(n_819),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_903),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_903),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_903),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_911),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_922),
.B(n_749),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_911),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_920),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_843),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_868),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_933),
.B(n_762),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_949),
.B(n_739),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_920),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_920),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_920),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_920),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_949),
.B(n_740),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_938),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_879),
.B(n_819),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_938),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_857),
.B(n_744),
.Y(n_1025)
);

AND2x2_ASAP7_75t_SL g1026 ( 
.A(n_858),
.B(n_399),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_938),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_843),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_938),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_834),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_938),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_953),
.B(n_740),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_941),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_869),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_869),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_941),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_918),
.B(n_742),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_941),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_953),
.B(n_742),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_890),
.A2(n_764),
.B1(n_776),
.B2(n_724),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_941),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_885),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_941),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_953),
.B(n_794),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_943),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_918),
.B(n_794),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_845),
.B(n_715),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_943),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_885),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_917),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_878),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_878),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_913),
.B(n_795),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_943),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_917),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_892),
.Y(n_1056)
);

AND2x6_ASAP7_75t_L g1057 ( 
.A(n_887),
.B(n_399),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_861),
.A2(n_802),
.B(n_799),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_943),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_943),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_953),
.B(n_799),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_881),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_922),
.B(n_802),
.Y(n_1063)
);

AND2x2_ASAP7_75t_SL g1064 ( 
.A(n_858),
.B(n_428),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_892),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_881),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_901),
.B(n_803),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_922),
.B(n_803),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_944),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_873),
.B(n_807),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_944),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_873),
.B(n_807),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_896),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_896),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_898),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_944),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_944),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_922),
.B(n_873),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_923),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_901),
.B(n_808),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_912),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_946),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_946),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_901),
.B(n_808),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_946),
.Y(n_1086)
);

NAND2x1_ASAP7_75t_L g1087 ( 
.A(n_901),
.B(n_829),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_946),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_946),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_923),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_947),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_947),
.Y(n_1092)
);

BUFx8_ASAP7_75t_L g1093 ( 
.A(n_856),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_873),
.B(n_809),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_898),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_947),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_947),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_899),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_899),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_908),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_947),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_908),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_924),
.B(n_809),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_924),
.B(n_810),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_928),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_891),
.A2(n_894),
.B(n_925),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_925),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_926),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_924),
.B(n_929),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_926),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_833),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_832),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_935),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_935),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_937),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_833),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_879),
.A2(n_594),
.B1(n_512),
.B2(n_415),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_937),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_939),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_922),
.B(n_810),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_939),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_952),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_952),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_832),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_837),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1047),
.B(n_867),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1107),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1057),
.A2(n_916),
.B1(n_900),
.B2(n_909),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1026),
.A2(n_858),
.B1(n_934),
.B2(n_861),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_958),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_958),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1026),
.A2(n_858),
.B1(n_934),
.B2(n_861),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_958),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1057),
.A2(n_902),
.B1(n_915),
.B2(n_826),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_959),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_969),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1107),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1108),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1026),
.A2(n_876),
.B1(n_910),
.B2(n_836),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_960),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1108),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1015),
.B(n_981),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_981),
.B(n_887),
.Y(n_1143)
);

BUFx8_ASAP7_75t_SL g1144 ( 
.A(n_994),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1110),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1000),
.Y(n_1146)
);

INVx4_ASAP7_75t_SL g1147 ( 
.A(n_1057),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1057),
.B(n_889),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_969),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_969),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_959),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_959),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_L g1153 ( 
.A(n_960),
.B(n_954),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1090),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1057),
.B(n_1071),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_967),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_963),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1090),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_967),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_982),
.B(n_1005),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1064),
.A2(n_876),
.B1(n_910),
.B2(n_836),
.Y(n_1161)
);

INVxp67_ASAP7_75t_SL g1162 ( 
.A(n_963),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1065),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_960),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1110),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1113),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1113),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_967),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1114),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_968),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1093),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1025),
.B(n_913),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1114),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1057),
.B(n_889),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1057),
.B(n_936),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_963),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_987),
.B(n_928),
.Y(n_1177)
);

INVxp33_ASAP7_75t_L g1178 ( 
.A(n_961),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1093),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1052),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1109),
.B(n_936),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_1053),
.Y(n_1182)
);

NOR2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1047),
.B(n_945),
.Y(n_1183)
);

INVx4_ASAP7_75t_SL g1184 ( 
.A(n_1057),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1115),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1052),
.B(n_951),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1052),
.B(n_922),
.Y(n_1187)
);

AND2x6_ASAP7_75t_L g1188 ( 
.A(n_992),
.B(n_924),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1063),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1071),
.B(n_954),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1056),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1080),
.B(n_1105),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1030),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1042),
.Y(n_1194)
);

NAND2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1087),
.B(n_849),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_1049),
.B(n_825),
.C(n_849),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1082),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_968),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1115),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1079),
.B(n_927),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1073),
.B(n_844),
.Y(n_1201)
);

INVx4_ASAP7_75t_SL g1202 ( 
.A(n_1079),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1073),
.B(n_1094),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1118),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1064),
.A2(n_876),
.B1(n_910),
.B2(n_836),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_974),
.A2(n_913),
.B1(n_929),
.B2(n_856),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_L g1207 ( 
.A(n_960),
.B(n_836),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1030),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1118),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1064),
.A2(n_876),
.B1(n_910),
.B2(n_836),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1079),
.B(n_927),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1119),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1119),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1093),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1094),
.B(n_1103),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1121),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_985),
.B(n_913),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_992),
.A2(n_876),
.B1(n_910),
.B2(n_836),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1103),
.B(n_877),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1079),
.B(n_931),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_974),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_968),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1104),
.B(n_929),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_972),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_972),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1121),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_960),
.B(n_931),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_972),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1122),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_974),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1104),
.B(n_929),
.Y(n_1231)
);

AND2x6_ASAP7_75t_L g1232 ( 
.A(n_993),
.B(n_841),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_963),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1040),
.A2(n_1117),
.B1(n_875),
.B2(n_1055),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1045),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_993),
.A2(n_876),
.B1(n_910),
.B2(n_836),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_974),
.B(n_841),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1122),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_966),
.B(n_1109),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1050),
.B(n_930),
.Y(n_1240)
);

INVx4_ASAP7_75t_SL g1241 ( 
.A(n_1063),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_996),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1123),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1045),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_978),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1063),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_996),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_997),
.A2(n_910),
.B1(n_876),
.B2(n_814),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_997),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_960),
.Y(n_1250)
);

CKINVDCx8_ASAP7_75t_R g1251 ( 
.A(n_989),
.Y(n_1251)
);

NAND2xp33_ASAP7_75t_L g1252 ( 
.A(n_964),
.B(n_859),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1123),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_978),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_955),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1014),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_978),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_964),
.B(n_930),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_966),
.A2(n_875),
.B1(n_845),
.B2(n_867),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_995),
.B(n_841),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_955),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_979),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_964),
.B(n_841),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_956),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_L g1265 ( 
.A(n_989),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1063),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_956),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1045),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_989),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_957),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_957),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_979),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_979),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_995),
.B(n_842),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_962),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1013),
.A2(n_814),
.B1(n_817),
.B2(n_812),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_962),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_964),
.B(n_842),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1013),
.A2(n_817),
.B1(n_820),
.B2(n_812),
.Y(n_1279)
);

INVx4_ASAP7_75t_SL g1280 ( 
.A(n_1069),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1069),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_965),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_989),
.B(n_912),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_984),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1069),
.B(n_839),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1016),
.Y(n_1286)
);

INVx4_ASAP7_75t_SL g1287 ( 
.A(n_1069),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_964),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_965),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1087),
.A2(n_416),
.B1(n_418),
.B2(n_413),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1045),
.Y(n_1291)
);

AO22x2_ASAP7_75t_L g1292 ( 
.A1(n_1016),
.A2(n_847),
.B1(n_870),
.B2(n_842),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_984),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_SL g1294 ( 
.A(n_1093),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_984),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1023),
.B(n_942),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1067),
.B(n_905),
.Y(n_1297)
);

NOR2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1021),
.B(n_945),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_1021),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1032),
.B(n_940),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1028),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1032),
.B(n_940),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1001),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1039),
.B(n_842),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_970),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1028),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_970),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1045),
.Y(n_1308)
);

INVxp33_ASAP7_75t_SL g1309 ( 
.A(n_1039),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1045),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_964),
.B(n_847),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1044),
.B(n_859),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1044),
.B(n_942),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_973),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1061),
.B(n_847),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_988),
.Y(n_1316)
);

INVxp67_ASAP7_75t_SL g1317 ( 
.A(n_971),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1001),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_973),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1061),
.B(n_847),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1010),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1301),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1301),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1160),
.A2(n_1058),
.B(n_977),
.C(n_1034),
.Y(n_1324)
);

AND2x6_ASAP7_75t_L g1325 ( 
.A(n_1147),
.B(n_1010),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1181),
.B(n_870),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1127),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1306),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1306),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1160),
.A2(n_915),
.B1(n_902),
.B2(n_1010),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1130),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1208),
.B(n_902),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1142),
.B(n_1037),
.Y(n_1333)
);

O2A1O1Ixp5_ASAP7_75t_L g1334 ( 
.A1(n_1263),
.A2(n_1074),
.B(n_1075),
.C(n_1066),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1201),
.B(n_1046),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1265),
.B(n_971),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1309),
.B(n_902),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1180),
.B(n_988),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1146),
.B(n_712),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1157),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1181),
.A2(n_1010),
.B1(n_1074),
.B2(n_1066),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1219),
.B(n_1081),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1221),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1297),
.B(n_1085),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1137),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1265),
.B(n_971),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1138),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1297),
.B(n_980),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1130),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1242),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1247),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1143),
.B(n_1181),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_SL g1353 ( 
.A(n_1163),
.B(n_932),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1141),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1234),
.A2(n_980),
.B(n_986),
.C(n_983),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1221),
.A2(n_1075),
.B1(n_870),
.B2(n_648),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1237),
.B(n_870),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1239),
.B(n_1028),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1221),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1203),
.B(n_1034),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1215),
.B(n_1034),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1299),
.B(n_977),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1230),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1223),
.B(n_1035),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1145),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1180),
.B(n_971),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1136),
.B(n_988),
.Y(n_1367)
);

NAND2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1163),
.B(n_1035),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1155),
.B(n_971),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1165),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1166),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1309),
.B(n_932),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1230),
.A2(n_1098),
.B1(n_1099),
.B2(n_1095),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1197),
.B(n_470),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1167),
.A2(n_1058),
.B(n_1051),
.C(n_1035),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1230),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1131),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1231),
.B(n_1051),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1269),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1131),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1260),
.B(n_1051),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1274),
.B(n_1062),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1128),
.B(n_971),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1304),
.B(n_1062),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1134),
.A2(n_1102),
.B1(n_1100),
.B2(n_1062),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1269),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1315),
.B(n_1076),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1133),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1169),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1133),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1320),
.B(n_1076),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1173),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1185),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1193),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1259),
.A2(n_1102),
.B1(n_1076),
.B2(n_1098),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1135),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1299),
.B(n_692),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1190),
.B(n_1095),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1286),
.B(n_1095),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1199),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1135),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_1249),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1204),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1209),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1182),
.B(n_1098),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1212),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1196),
.B(n_1009),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1151),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1151),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_1149),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1152),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1182),
.B(n_1099),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1152),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1182),
.B(n_1099),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1157),
.B(n_1008),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1213),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1157),
.B(n_1008),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1172),
.B(n_1100),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1172),
.B(n_1100),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1216),
.B(n_1102),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1226),
.B(n_983),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1176),
.B(n_1008),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1229),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1269),
.B(n_975),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1238),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1186),
.A2(n_988),
.B1(n_1017),
.B2(n_1011),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1256),
.B(n_726),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1243),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1144),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1156),
.Y(n_1430)
);

AO221x1_ASAP7_75t_L g1431 ( 
.A1(n_1292),
.A2(n_607),
.B1(n_666),
.B2(n_552),
.C(n_539),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_SL g1432 ( 
.A(n_1191),
.B(n_723),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1253),
.A2(n_990),
.B1(n_991),
.B2(n_986),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1255),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1140),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1251),
.B(n_831),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1261),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1217),
.B(n_990),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1175),
.A2(n_1111),
.B1(n_1125),
.B2(n_1116),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1217),
.B(n_1148),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1156),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1178),
.B(n_831),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1154),
.Y(n_1443)
);

AND2x6_ASAP7_75t_SL g1444 ( 
.A(n_1240),
.B(n_539),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1174),
.B(n_991),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1159),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1177),
.B(n_975),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1264),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1129),
.A2(n_1111),
.B1(n_1125),
.B2(n_1116),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1171),
.B(n_1179),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1176),
.B(n_1147),
.Y(n_1451)
);

NOR3xp33_ASAP7_75t_L g1452 ( 
.A(n_1186),
.B(n_603),
.C(n_531),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_SL g1453 ( 
.A(n_1171),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1158),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1159),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1267),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1292),
.B(n_1001),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1270),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1149),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1126),
.B(n_723),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1292),
.B(n_1001),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1168),
.Y(n_1462)
);

NOR3xp33_ASAP7_75t_L g1463 ( 
.A(n_1194),
.B(n_1192),
.C(n_1312),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1168),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1271),
.A2(n_1003),
.B(n_1002),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_L g1466 ( 
.A(n_1179),
.B(n_1009),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1170),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1176),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1276),
.B(n_1019),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1170),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1276),
.B(n_1019),
.Y(n_1471)
);

NOR2xp67_ASAP7_75t_L g1472 ( 
.A(n_1214),
.B(n_1009),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1178),
.B(n_1017),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1429),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1327),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1337),
.A2(n_1191),
.B1(n_1302),
.B2(n_1300),
.Y(n_1476)
);

BUFx4f_ASAP7_75t_L g1477 ( 
.A(n_1450),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1350),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1443),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1345),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1450),
.B(n_1202),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1344),
.B(n_1188),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1429),
.Y(n_1483)
);

O2A1O1Ixp5_ASAP7_75t_L g1484 ( 
.A1(n_1368),
.A2(n_1258),
.B(n_1227),
.C(n_1136),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1450),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1460),
.B(n_1283),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1397),
.B(n_1313),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1335),
.B(n_1188),
.Y(n_1488)
);

O2A1O1Ixp5_ASAP7_75t_L g1489 ( 
.A1(n_1368),
.A2(n_1258),
.B(n_1227),
.C(n_1136),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1333),
.B(n_1188),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1347),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1332),
.B(n_1394),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1323),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1460),
.B(n_1296),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1354),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1463),
.B(n_1206),
.Y(n_1496)
);

AND2x6_ASAP7_75t_L g1497 ( 
.A(n_1424),
.B(n_1214),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1365),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1370),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1454),
.B(n_1240),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1342),
.B(n_1188),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1348),
.B(n_1447),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1343),
.B(n_1150),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1450),
.B(n_1202),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1374),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1323),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1372),
.B(n_1202),
.Y(n_1507)
);

NOR2x2_ASAP7_75t_L g1508 ( 
.A(n_1353),
.B(n_1240),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1324),
.A2(n_1319),
.B(n_1277),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1447),
.B(n_1188),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1328),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1330),
.A2(n_1442),
.B1(n_1356),
.B2(n_1436),
.Y(n_1512)
);

NOR2x2_ASAP7_75t_L g1513 ( 
.A(n_1432),
.B(n_1144),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1435),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1352),
.B(n_1321),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_SL g1516 ( 
.A(n_1397),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1435),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1358),
.B(n_1275),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1325),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1360),
.B(n_1282),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1326),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1435),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1326),
.B(n_1339),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1435),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1343),
.B(n_1298),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1375),
.A2(n_1187),
.B(n_999),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1359),
.B(n_1150),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1371),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1389),
.Y(n_1529)
);

INVx5_ASAP7_75t_L g1530 ( 
.A(n_1325),
.Y(n_1530)
);

NOR2x1_ASAP7_75t_L g1531 ( 
.A(n_1405),
.B(n_1183),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1427),
.B(n_1294),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1361),
.B(n_1289),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1359),
.B(n_1241),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1453),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1412),
.A2(n_1290),
.B(n_1252),
.C(n_1311),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1363),
.B(n_1150),
.Y(n_1537)
);

INVx5_ASAP7_75t_L g1538 ( 
.A(n_1325),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1453),
.Y(n_1539)
);

OAI22x1_ASAP7_75t_L g1540 ( 
.A1(n_1392),
.A2(n_1278),
.B1(n_1311),
.B2(n_1263),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1398),
.B(n_1305),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1457),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1452),
.A2(n_1195),
.B1(n_1294),
.B2(n_1232),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1440),
.A2(n_1195),
.B(n_1314),
.C(n_1307),
.Y(n_1544)
);

AOI22x1_ASAP7_75t_L g1545 ( 
.A1(n_1340),
.A2(n_1162),
.B1(n_1316),
.B2(n_1233),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1328),
.Y(n_1546)
);

AND2x6_ASAP7_75t_SL g1547 ( 
.A(n_1473),
.B(n_499),
.Y(n_1547)
);

O2A1O1Ixp5_ASAP7_75t_L g1548 ( 
.A1(n_1418),
.A2(n_1187),
.B(n_1278),
.C(n_1244),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_L g1549 ( 
.A(n_1325),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1393),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1363),
.B(n_1241),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1453),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1459),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1351),
.A2(n_1189),
.B1(n_1266),
.B2(n_1246),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1400),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1376),
.B(n_1285),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1414),
.B(n_1189),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1376),
.B(n_1241),
.Y(n_1558)
);

INVx5_ASAP7_75t_L g1559 ( 
.A(n_1325),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1403),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1364),
.B(n_1233),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1492),
.B(n_1379),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1476),
.B(n_1379),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_SL g1564 ( 
.A(n_1502),
.B(n_1482),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1487),
.B(n_604),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1554),
.B(n_1386),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1530),
.B(n_1386),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1486),
.B(n_604),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_SL g1569 ( 
.A(n_1482),
.B(n_1435),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_SL g1570 ( 
.A(n_1507),
.B(n_1378),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1494),
.B(n_1404),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1530),
.B(n_1459),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1530),
.B(n_1538),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1530),
.B(n_1395),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1538),
.B(n_1402),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1538),
.B(n_1559),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1479),
.B(n_1406),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1538),
.B(n_1385),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1559),
.B(n_1466),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1559),
.B(n_1472),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1559),
.B(n_1341),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_SL g1582 ( 
.A(n_1490),
.B(n_1416),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1478),
.B(n_1423),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1490),
.B(n_1410),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1488),
.B(n_1288),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1523),
.B(n_1425),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1488),
.B(n_1288),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1512),
.B(n_1428),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1515),
.B(n_1288),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1521),
.B(n_1434),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1549),
.B(n_1543),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_SL g1592 ( 
.A(n_1502),
.B(n_1340),
.Y(n_1592)
);

AND2x4_ASAP7_75t_SL g1593 ( 
.A(n_1481),
.B(n_1246),
.Y(n_1593)
);

NAND2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1474),
.B(n_1340),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1518),
.B(n_1468),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1549),
.B(n_1140),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1475),
.B(n_1399),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1557),
.B(n_1501),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1532),
.B(n_1505),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_SL g1600 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1501),
.B(n_1140),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1500),
.B(n_1553),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1496),
.B(n_1140),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1531),
.B(n_1164),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1520),
.B(n_1164),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1533),
.B(n_1164),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1533),
.B(n_1164),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1541),
.B(n_1288),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1541),
.B(n_1519),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1519),
.B(n_1514),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1514),
.B(n_1336),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1561),
.B(n_1468),
.Y(n_1612)
);

NAND2xp33_ASAP7_75t_SL g1613 ( 
.A(n_1561),
.B(n_1468),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1480),
.B(n_1437),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1612),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1599),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1588),
.A2(n_1431),
.B1(n_1132),
.B2(n_1129),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1600),
.B(n_1542),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1563),
.B(n_1547),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1593),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1585),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1593),
.Y(n_1622)
);

AND3x1_ASAP7_75t_SL g1623 ( 
.A(n_1594),
.B(n_530),
.C(n_506),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1600),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1545),
.Y(n_1626)
);

CKINVDCx8_ASAP7_75t_R g1627 ( 
.A(n_1591),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1497),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1583),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1564),
.A2(n_1536),
.B(n_1544),
.C(n_1355),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1614),
.B(n_1509),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1564),
.B(n_1497),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1571),
.B(n_1509),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1603),
.B(n_1526),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_R g1637 ( 
.A(n_1592),
.B(n_1535),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1605),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1609),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1606),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1607),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1597),
.B(n_1497),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1586),
.B(n_1497),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1592),
.A2(n_1489),
.B(n_1484),
.C(n_1548),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1608),
.B(n_1526),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1582),
.B(n_1491),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1574),
.B(n_1510),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1613),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1584),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1325),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1589),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1565),
.B(n_1362),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1590),
.B(n_1362),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1566),
.B(n_1495),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1573),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1569),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1577),
.B(n_1431),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1568),
.B(n_1424),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1570),
.B(n_1510),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1610),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1575),
.Y(n_1662)
);

AND3x1_ASAP7_75t_SL g1663 ( 
.A(n_1562),
.B(n_530),
.C(n_506),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1578),
.B(n_1540),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1624),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1633),
.B(n_1498),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1616),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1635),
.A2(n_1383),
.B(n_1576),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1629),
.Y(n_1669)
);

AO21x2_ASAP7_75t_L g1670 ( 
.A1(n_1664),
.A2(n_1375),
.B(n_1581),
.Y(n_1670)
);

INVx4_ASAP7_75t_SL g1671 ( 
.A(n_1615),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1629),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1637),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1627),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1499),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1629),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1635),
.A2(n_1383),
.B(n_1334),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1629),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1615),
.B(n_1481),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1644),
.A2(n_1324),
.B(n_1419),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1632),
.A2(n_1465),
.B(n_1572),
.Y(n_1681)
);

INVx6_ASAP7_75t_L g1682 ( 
.A(n_1656),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1633),
.B(n_1528),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1640),
.Y(n_1684)
);

BUFx12f_ASAP7_75t_L g1685 ( 
.A(n_1652),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1644),
.A2(n_1624),
.B(n_1630),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1620),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1620),
.Y(n_1688)
);

NAND2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1656),
.B(n_1477),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1645),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

BUFx8_ASAP7_75t_L g1692 ( 
.A(n_1659),
.Y(n_1692)
);

AO21x1_ASAP7_75t_L g1693 ( 
.A1(n_1646),
.A2(n_1602),
.B(n_822),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1632),
.A2(n_1567),
.B(n_1579),
.Y(n_1694)
);

BUFx2_ASAP7_75t_SL g1695 ( 
.A(n_1656),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1630),
.A2(n_1252),
.B(n_1407),
.Y(n_1696)
);

NAND2x1p5_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1477),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1640),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1664),
.A2(n_1646),
.B(n_1618),
.Y(n_1699)
);

INVx6_ASAP7_75t_L g1700 ( 
.A(n_1656),
.Y(n_1700)
);

BUFx12f_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1615),
.B(n_1634),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1645),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1645),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1640),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1627),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1651),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1627),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1634),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1626),
.A2(n_1451),
.B(n_1596),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1660),
.A2(n_1580),
.B(n_1417),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1631),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1653),
.B(n_1529),
.Y(n_1713)
);

CKINVDCx16_ASAP7_75t_R g1714 ( 
.A(n_1637),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1651),
.Y(n_1715)
);

BUFx4f_ASAP7_75t_SL g1716 ( 
.A(n_1620),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1623),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1621),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1660),
.A2(n_1417),
.B(n_1415),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1631),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1620),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1657),
.Y(n_1722)
);

BUFx10_ASAP7_75t_L g1723 ( 
.A(n_1619),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1631),
.B(n_1550),
.Y(n_1724)
);

CKINVDCx11_ASAP7_75t_R g1725 ( 
.A(n_1662),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1634),
.B(n_1514),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1619),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1621),
.A2(n_1422),
.B(n_1415),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1651),
.Y(n_1729)
);

BUFx12f_ASAP7_75t_L g1730 ( 
.A(n_1652),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1620),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1622),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1621),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1648),
.A2(n_820),
.B(n_824),
.C(n_822),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1618),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1638),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1638),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1622),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1625),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1662),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1625),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1622),
.Y(n_1742)
);

AO21x2_ASAP7_75t_L g1743 ( 
.A1(n_1643),
.A2(n_1461),
.B(n_1438),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1648),
.Y(n_1744)
);

AO21x2_ASAP7_75t_L g1745 ( 
.A1(n_1643),
.A2(n_1369),
.B(n_1420),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1626),
.A2(n_829),
.B(n_824),
.Y(n_1746)
);

INVx8_ASAP7_75t_L g1747 ( 
.A(n_1647),
.Y(n_1747)
);

CKINVDCx14_ASAP7_75t_R g1748 ( 
.A(n_1659),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1625),
.A2(n_1422),
.B(n_1366),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1636),
.A2(n_1366),
.B(n_1369),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1717),
.A2(n_1623),
.B1(n_1663),
.B2(n_1658),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1670),
.A2(n_1647),
.B1(n_1659),
.B2(n_1658),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1718),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1670),
.A2(n_1647),
.B1(n_1658),
.B2(n_1617),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1686),
.A2(n_1648),
.B1(n_1654),
.B2(n_1650),
.Y(n_1755)
);

INVx6_ASAP7_75t_L g1756 ( 
.A(n_1714),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1718),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1676),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1686),
.A2(n_1654),
.B1(n_1650),
.B2(n_1642),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_1708),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1670),
.A2(n_1647),
.B1(n_1617),
.B2(n_1642),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1733),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1746),
.A2(n_1639),
.B(n_1641),
.Y(n_1763)
);

BUFx4_ASAP7_75t_R g1764 ( 
.A(n_1723),
.Y(n_1764)
);

BUFx10_ASAP7_75t_L g1765 ( 
.A(n_1674),
.Y(n_1765)
);

BUFx2_ASAP7_75t_SL g1766 ( 
.A(n_1667),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1736),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1736),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1702),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1685),
.A2(n_1647),
.B1(n_1628),
.B2(n_1653),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1737),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1727),
.A2(n_1647),
.B1(n_1628),
.B2(n_1639),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1733),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1739),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1739),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1737),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1706),
.B(n_1655),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1671),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1722),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_SL g1780 ( 
.A1(n_1686),
.A2(n_1653),
.B1(n_1663),
.B2(n_1647),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1727),
.A2(n_1525),
.B1(n_1649),
.B2(n_1657),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1735),
.Y(n_1782)
);

CKINVDCx6p67_ASAP7_75t_R g1783 ( 
.A(n_1714),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1735),
.Y(n_1784)
);

OAI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1674),
.A2(n_1649),
.B1(n_1622),
.B2(n_1662),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1684),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1671),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1685),
.A2(n_1516),
.B1(n_1506),
.B2(n_1511),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1665),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1665),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1741),
.Y(n_1791)
);

BUFx8_ASAP7_75t_L g1792 ( 
.A(n_1701),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1741),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1723),
.B(n_1655),
.Y(n_1794)
);

BUFx10_ASAP7_75t_L g1795 ( 
.A(n_1726),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1712),
.Y(n_1796)
);

INVx6_ASAP7_75t_L g1797 ( 
.A(n_1706),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1706),
.Y(n_1798)
);

NAND2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1706),
.B(n_1655),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1712),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1671),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1720),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1748),
.A2(n_1661),
.B1(n_1622),
.B2(n_1649),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1706),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1720),
.B(n_1641),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1690),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1701),
.A2(n_1546),
.B1(n_1493),
.B2(n_1232),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1690),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1731),
.Y(n_1809)
);

CKINVDCx6p67_ASAP7_75t_R g1810 ( 
.A(n_1723),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1684),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1703),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1702),
.B(n_1662),
.Y(n_1813)
);

INVx6_ASAP7_75t_L g1814 ( 
.A(n_1692),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1691),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1699),
.Y(n_1816)
);

NAND2x1p5_ASAP7_75t_L g1817 ( 
.A(n_1709),
.B(n_1636),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1686),
.A2(n_641),
.B1(n_672),
.B2(n_1661),
.Y(n_1818)
);

OAI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1679),
.A2(n_1636),
.B1(n_1556),
.B2(n_1525),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1703),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1699),
.B(n_532),
.Y(n_1821)
);

CKINVDCx6p67_ASAP7_75t_R g1822 ( 
.A(n_1723),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1704),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1704),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1724),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1730),
.A2(n_1232),
.B1(n_1485),
.B2(n_1555),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1671),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1691),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1699),
.A2(n_641),
.B1(n_672),
.B2(n_614),
.Y(n_1829)
);

OAI22x1_ASAP7_75t_L g1830 ( 
.A1(n_1702),
.A2(n_1513),
.B1(n_1552),
.B2(n_1539),
.Y(n_1830)
);

BUFx10_ASAP7_75t_L g1831 ( 
.A(n_1726),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1680),
.A2(n_1451),
.B(n_1382),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1725),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1716),
.Y(n_1834)
);

CKINVDCx11_ASAP7_75t_R g1835 ( 
.A(n_1673),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1724),
.Y(n_1836)
);

CKINVDCx8_ASAP7_75t_R g1837 ( 
.A(n_1695),
.Y(n_1837)
);

BUFx12f_ASAP7_75t_L g1838 ( 
.A(n_1730),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1679),
.A2(n_1556),
.B1(n_1525),
.B2(n_542),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1702),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1679),
.A2(n_1556),
.B1(n_1560),
.B2(n_542),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1743),
.A2(n_1232),
.B1(n_1329),
.B2(n_1322),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1743),
.A2(n_1232),
.B1(n_1329),
.B2(n_1322),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1709),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1698),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1713),
.A2(n_1666),
.B1(n_1683),
.B2(n_1675),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1743),
.A2(n_1693),
.B1(n_1747),
.B2(n_1696),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1698),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1679),
.A2(n_552),
.B1(n_572),
.B2(n_532),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1680),
.A2(n_672),
.B1(n_641),
.B2(n_576),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1672),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1693),
.A2(n_1132),
.B1(n_1384),
.B2(n_1381),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1744),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1707),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1747),
.A2(n_1391),
.B1(n_1387),
.B2(n_1349),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1669),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1669),
.Y(n_1857)
);

BUFx12f_ASAP7_75t_L g1858 ( 
.A(n_1731),
.Y(n_1858)
);

BUFx12f_ASAP7_75t_L g1859 ( 
.A(n_1731),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1680),
.A2(n_576),
.B1(n_577),
.B2(n_572),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1680),
.A2(n_598),
.B1(n_599),
.B2(n_577),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1747),
.A2(n_599),
.B1(n_600),
.B2(n_598),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_SL g1863 ( 
.A1(n_1747),
.A2(n_607),
.B1(n_609),
.B2(n_600),
.Y(n_1863)
);

BUFx4_ASAP7_75t_R g1864 ( 
.A(n_1687),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1747),
.A2(n_1349),
.B1(n_1377),
.B2(n_1331),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1687),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1740),
.Y(n_1867)
);

CKINVDCx20_ASAP7_75t_R g1868 ( 
.A(n_1692),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1679),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1740),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1692),
.A2(n_1377),
.B1(n_1380),
.B2(n_1331),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1692),
.A2(n_1380),
.B1(n_1390),
.B2(n_1388),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1707),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1707),
.Y(n_1874)
);

BUFx4f_ASAP7_75t_SL g1875 ( 
.A(n_1688),
.Y(n_1875)
);

BUFx4f_ASAP7_75t_SL g1876 ( 
.A(n_1688),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1678),
.B(n_609),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1715),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1731),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1715),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1709),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1705),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1744),
.Y(n_1883)
);

INVx6_ASAP7_75t_L g1884 ( 
.A(n_1726),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1715),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1729),
.Y(n_1886)
);

BUFx12f_ASAP7_75t_L g1887 ( 
.A(n_1731),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1734),
.A2(n_613),
.B1(n_617),
.B2(n_611),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1729),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1745),
.A2(n_1388),
.B1(n_1396),
.B2(n_1390),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1729),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1744),
.Y(n_1892)
);

INVx6_ASAP7_75t_L g1893 ( 
.A(n_1726),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1745),
.A2(n_1396),
.B1(n_1408),
.B2(n_1401),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1689),
.A2(n_1504),
.B1(n_1604),
.B2(n_1551),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1745),
.A2(n_1401),
.B1(n_1409),
.B2(n_1408),
.Y(n_1896)
);

CKINVDCx11_ASAP7_75t_R g1897 ( 
.A(n_1732),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1705),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1678),
.A2(n_1409),
.B1(n_1413),
.B2(n_1411),
.Y(n_1899)
);

BUFx12f_ASAP7_75t_L g1900 ( 
.A(n_1732),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1738),
.Y(n_1901)
);

CKINVDCx20_ASAP7_75t_R g1902 ( 
.A(n_1738),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1785),
.A2(n_1710),
.B(n_1697),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1754),
.A2(n_1504),
.B1(n_1413),
.B2(n_1430),
.Y(n_1904)
);

AOI222xp33_ASAP7_75t_L g1905 ( 
.A1(n_1849),
.A2(n_619),
.B1(n_613),
.B2(n_623),
.C1(n_617),
.C2(n_611),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1846),
.B(n_1779),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1785),
.A2(n_1697),
.B(n_1689),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1833),
.Y(n_1908)
);

AOI21xp33_ASAP7_75t_L g1909 ( 
.A1(n_1829),
.A2(n_623),
.B(n_619),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1856),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1782),
.B(n_1705),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1756),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1755),
.A2(n_1697),
.B(n_1689),
.Y(n_1913)
);

OA21x2_ASAP7_75t_L g1914 ( 
.A1(n_1821),
.A2(n_1668),
.B(n_1694),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1784),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1857),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1760),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1806),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_L g1919 ( 
.A1(n_1821),
.A2(n_1668),
.B(n_1711),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1818),
.A2(n_1430),
.B1(n_1441),
.B2(n_1411),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1825),
.B(n_1721),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1808),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1812),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1755),
.A2(n_1719),
.B(n_1711),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1805),
.B(n_1695),
.Y(n_1925)
);

AO21x2_ASAP7_75t_L g1926 ( 
.A1(n_1816),
.A2(n_1677),
.B(n_1750),
.Y(n_1926)
);

OAI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1829),
.A2(n_633),
.B1(n_637),
.B2(n_628),
.C(n_624),
.Y(n_1927)
);

OA21x2_ASAP7_75t_L g1928 ( 
.A1(n_1816),
.A2(n_1694),
.B(n_1719),
.Y(n_1928)
);

OAI211xp5_ASAP7_75t_L g1929 ( 
.A1(n_1850),
.A2(n_628),
.B(n_633),
.C(n_624),
.Y(n_1929)
);

OA21x2_ASAP7_75t_L g1930 ( 
.A1(n_1805),
.A2(n_1677),
.B(n_1681),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1756),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1756),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1836),
.B(n_1682),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1753),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1757),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1762),
.Y(n_1936)
);

OAI21xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1787),
.A2(n_1681),
.B(n_1728),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1794),
.A2(n_1728),
.B(n_1749),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1820),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1823),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1763),
.A2(n_1847),
.B(n_1832),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1824),
.Y(n_1942)
);

CKINVDCx11_ASAP7_75t_R g1943 ( 
.A(n_1835),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1850),
.A2(n_642),
.B(n_637),
.Y(n_1944)
);

INVx4_ASAP7_75t_L g1945 ( 
.A(n_1864),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1851),
.B(n_1742),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1763),
.A2(n_1749),
.B(n_1750),
.Y(n_1947)
);

BUFx3_ASAP7_75t_L g1948 ( 
.A(n_1758),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1818),
.A2(n_1446),
.B1(n_1455),
.B2(n_1441),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1773),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1840),
.B(n_1682),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1751),
.A2(n_649),
.B(n_653),
.C(n_642),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1849),
.A2(n_451),
.B1(n_463),
.B2(n_449),
.C(n_443),
.Y(n_1953)
);

OAI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1860),
.A2(n_653),
.B(n_649),
.Y(n_1954)
);

NAND2x1p5_ASAP7_75t_L g1955 ( 
.A(n_1869),
.B(n_1742),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1789),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1790),
.B(n_1682),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1774),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1752),
.A2(n_670),
.B(n_684),
.C(n_656),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1772),
.A2(n_1732),
.B(n_1558),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1772),
.A2(n_1732),
.B(n_1534),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1769),
.B(n_1682),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1796),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1860),
.A2(n_1732),
.B(n_1346),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1800),
.B(n_656),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1802),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1765),
.B(n_1483),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1767),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1869),
.B(n_1700),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1877),
.B(n_1768),
.Y(n_1970)
);

NOR2xp67_ASAP7_75t_R g1971 ( 
.A(n_1814),
.B(n_1700),
.Y(n_1971)
);

INVx1_ASAP7_75t_SL g1972 ( 
.A(n_1853),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1780),
.A2(n_1455),
.B1(n_1462),
.B2(n_1446),
.Y(n_1973)
);

AO21x1_ASAP7_75t_L g1974 ( 
.A1(n_1877),
.A2(n_670),
.B(n_666),
.Y(n_1974)
);

A2O1A1Ixp33_ASAP7_75t_L g1975 ( 
.A1(n_1780),
.A2(n_684),
.B(n_677),
.C(n_449),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1867),
.Y(n_1976)
);

OAI21xp33_ASAP7_75t_L g1977 ( 
.A1(n_1861),
.A2(n_677),
.B(n_451),
.Y(n_1977)
);

AOI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1861),
.A2(n_463),
.B(n_443),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1870),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1771),
.B(n_1700),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1832),
.A2(n_1527),
.B(n_1503),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1776),
.B(n_1700),
.Y(n_1982)
);

AND2x4_ASAP7_75t_SL g1983 ( 
.A(n_1783),
.B(n_1517),
.Y(n_1983)
);

AO31x2_ASAP7_75t_L g1984 ( 
.A1(n_1803),
.A2(n_1848),
.A3(n_1775),
.B(n_1793),
.Y(n_1984)
);

OAI211xp5_ASAP7_75t_L g1985 ( 
.A1(n_1781),
.A2(n_647),
.B(n_536),
.C(n_436),
.Y(n_1985)
);

OR2x6_ASAP7_75t_L g1986 ( 
.A(n_1778),
.B(n_1517),
.Y(n_1986)
);

INVx3_ASAP7_75t_L g1987 ( 
.A(n_1769),
.Y(n_1987)
);

AO31x2_ASAP7_75t_L g1988 ( 
.A1(n_1803),
.A2(n_647),
.A3(n_536),
.B(n_837),
.Y(n_1988)
);

AO31x2_ASAP7_75t_L g1989 ( 
.A1(n_1791),
.A2(n_850),
.A3(n_851),
.B(n_848),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1786),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1761),
.A2(n_1464),
.B1(n_1467),
.B2(n_1462),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1766),
.Y(n_1992)
);

OAI21x1_ASAP7_75t_L g1993 ( 
.A1(n_1777),
.A2(n_1527),
.B(n_1503),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1811),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1888),
.A2(n_457),
.B(n_754),
.C(n_752),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1765),
.Y(n_1996)
);

AO31x2_ASAP7_75t_L g1997 ( 
.A1(n_1815),
.A2(n_850),
.A3(n_851),
.B(n_848),
.Y(n_1997)
);

AO21x2_ASAP7_75t_L g1998 ( 
.A1(n_1819),
.A2(n_756),
.B(n_755),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1792),
.Y(n_1999)
);

OAI21x1_ASAP7_75t_L g2000 ( 
.A1(n_1777),
.A2(n_1537),
.B(n_1346),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1828),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1845),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1862),
.A2(n_457),
.B(n_484),
.Y(n_2003)
);

AO21x2_ASAP7_75t_L g2004 ( 
.A1(n_1819),
.A2(n_1874),
.B(n_1873),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1878),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1787),
.A2(n_1336),
.B(n_1537),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1880),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1842),
.A2(n_1467),
.B1(n_1470),
.B2(n_1464),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1886),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1854),
.Y(n_2010)
);

AOI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1827),
.A2(n_1524),
.B(n_1522),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1813),
.B(n_757),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1827),
.A2(n_1524),
.B(n_1522),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1844),
.B(n_759),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1882),
.B(n_761),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1885),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1898),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1889),
.Y(n_2018)
);

AO21x2_ASAP7_75t_L g2019 ( 
.A1(n_1891),
.A2(n_766),
.B(n_765),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1882),
.B(n_767),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1801),
.B(n_1517),
.Y(n_2021)
);

OA21x2_ASAP7_75t_L g2022 ( 
.A1(n_1883),
.A2(n_769),
.B(n_768),
.Y(n_2022)
);

NOR2x1_ASAP7_75t_SL g2023 ( 
.A(n_1838),
.B(n_1834),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1892),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1884),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1884),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1853),
.B(n_770),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1759),
.A2(n_1839),
.B(n_1830),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1834),
.B(n_771),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1881),
.B(n_773),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_1888),
.A2(n_440),
.B1(n_458),
.B2(n_437),
.C(n_423),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1881),
.B(n_775),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1884),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1862),
.A2(n_460),
.B1(n_467),
.B2(n_465),
.Y(n_2034)
);

OAI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1863),
.A2(n_514),
.B(n_484),
.Y(n_2035)
);

AO31x2_ASAP7_75t_L g2036 ( 
.A1(n_1759),
.A2(n_853),
.A3(n_855),
.B(n_852),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1893),
.B(n_777),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1792),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1817),
.B(n_779),
.Y(n_2039)
);

OA21x2_ASAP7_75t_L g2040 ( 
.A1(n_1770),
.A2(n_782),
.B(n_781),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1817),
.B(n_1901),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1866),
.B(n_783),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1843),
.A2(n_1470),
.B1(n_469),
.B2(n_511),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_1893),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1893),
.Y(n_2045)
);

AO21x2_ASAP7_75t_L g2046 ( 
.A1(n_1839),
.A2(n_787),
.B(n_785),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1798),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1902),
.B(n_788),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1810),
.B(n_1822),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1855),
.A2(n_1863),
.B1(n_1852),
.B2(n_1807),
.Y(n_2050)
);

INVx2_ASAP7_75t_SL g2051 ( 
.A(n_1795),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1809),
.B(n_789),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1795),
.Y(n_2053)
);

INVxp67_ASAP7_75t_L g2054 ( 
.A(n_1809),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1831),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1841),
.A2(n_1524),
.B(n_1522),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1865),
.A2(n_469),
.B1(n_511),
.B2(n_1448),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_SL g2058 ( 
.A1(n_2028),
.A2(n_1764),
.B(n_1826),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1941),
.A2(n_1868),
.B1(n_1814),
.B2(n_1875),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1943),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_2050),
.A2(n_1814),
.B1(n_1837),
.B2(n_1876),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1998),
.A2(n_1909),
.B1(n_2046),
.B2(n_1904),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1956),
.Y(n_2063)
);

OA21x2_ASAP7_75t_L g2064 ( 
.A1(n_1906),
.A2(n_1894),
.B(n_1890),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_1998),
.A2(n_1788),
.B1(n_1872),
.B2(n_1871),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1945),
.B(n_1809),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1903),
.A2(n_1799),
.B(n_1896),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1968),
.Y(n_2068)
);

OAI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1945),
.A2(n_1913),
.B1(n_1907),
.B2(n_2040),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1909),
.A2(n_1899),
.B1(n_1895),
.B2(n_1831),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_SL g2071 ( 
.A1(n_2004),
.A2(n_1985),
.B1(n_2046),
.B2(n_2040),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1952),
.A2(n_1799),
.B(n_588),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1917),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1991),
.A2(n_1456),
.B1(n_1458),
.B2(n_1797),
.Y(n_2074)
);

BUFx4f_ASAP7_75t_SL g2075 ( 
.A(n_1948),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1915),
.Y(n_2076)
);

NAND3xp33_ASAP7_75t_L g2077 ( 
.A(n_1937),
.B(n_1879),
.C(n_1804),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1931),
.Y(n_2078)
);

OAI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2022),
.A2(n_1804),
.B1(n_1798),
.B2(n_1797),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_2003),
.A2(n_1797),
.B1(n_1804),
.B2(n_1798),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2003),
.A2(n_567),
.B1(n_588),
.B2(n_514),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_SL g2082 ( 
.A1(n_2004),
.A2(n_1859),
.B1(n_1887),
.B2(n_1858),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2005),
.B(n_1879),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2007),
.B(n_2009),
.Y(n_2084)
);

AOI221xp5_ASAP7_75t_SL g2085 ( 
.A1(n_1924),
.A2(n_791),
.B1(n_790),
.B2(n_1879),
.C(n_3),
.Y(n_2085)
);

OAI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2022),
.A2(n_1900),
.B1(n_1508),
.B2(n_1444),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1944),
.A2(n_567),
.B1(n_853),
.B2(n_852),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2017),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_2038),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1919),
.A2(n_1897),
.B(n_1433),
.Y(n_2090)
);

AOI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_1927),
.A2(n_473),
.B1(n_483),
.B2(n_477),
.C(n_468),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_1975),
.A2(n_498),
.B1(n_503),
.B2(n_501),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1911),
.B(n_504),
.Y(n_2093)
);

OAI221xp5_ASAP7_75t_L g2094 ( 
.A1(n_1944),
.A2(n_508),
.B1(n_517),
.B2(n_515),
.C(n_510),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1973),
.A2(n_567),
.B1(n_864),
.B2(n_855),
.Y(n_2095)
);

NAND2x1_ASAP7_75t_L g2096 ( 
.A(n_1912),
.B(n_452),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1932),
.B(n_1),
.Y(n_2097)
);

OAI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1960),
.A2(n_520),
.B1(n_524),
.B2(n_521),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1912),
.B(n_2),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1910),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1992),
.Y(n_2101)
);

OAI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_1961),
.A2(n_527),
.B1(n_537),
.B2(n_525),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1918),
.Y(n_2103)
);

INVx4_ASAP7_75t_L g2104 ( 
.A(n_1996),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_1905),
.A2(n_865),
.B1(n_871),
.B2(n_864),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1969),
.B(n_2),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1922),
.Y(n_2107)
);

NAND4xp25_ASAP7_75t_L g2108 ( 
.A(n_2029),
.B(n_2014),
.C(n_2032),
.D(n_2030),
.Y(n_2108)
);

AOI31xp33_ASAP7_75t_L g2109 ( 
.A1(n_1999),
.A2(n_544),
.A3(n_545),
.B(n_538),
.Y(n_2109)
);

OAI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1964),
.A2(n_551),
.B1(n_557),
.B2(n_548),
.Y(n_2110)
);

INVx1_ASAP7_75t_SL g2111 ( 
.A(n_2048),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1951),
.B(n_3),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_1976),
.Y(n_2113)
);

OAI21xp33_ASAP7_75t_L g2114 ( 
.A1(n_1925),
.A2(n_561),
.B(n_558),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1923),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_1911),
.B(n_4),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2024),
.B(n_4),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_1908),
.Y(n_2118)
);

INVx8_ASAP7_75t_L g2119 ( 
.A(n_2037),
.Y(n_2119)
);

OAI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_2012),
.A2(n_564),
.B1(n_569),
.B2(n_563),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1905),
.A2(n_871),
.B1(n_872),
.B2(n_865),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1979),
.B(n_570),
.Y(n_2122)
);

INVxp67_ASAP7_75t_L g2123 ( 
.A(n_2042),
.Y(n_2123)
);

OA21x2_ASAP7_75t_L g2124 ( 
.A1(n_1925),
.A2(n_578),
.B(n_573),
.Y(n_2124)
);

AOI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_2034),
.A2(n_590),
.B1(n_608),
.B2(n_589),
.C(n_581),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1939),
.Y(n_2126)
);

OAI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_2015),
.A2(n_620),
.B(n_626),
.C(n_612),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2034),
.A2(n_634),
.B1(n_639),
.B2(n_631),
.C(n_630),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1972),
.B(n_650),
.Y(n_2129)
);

O2A1O1Ixp33_ASAP7_75t_L g2130 ( 
.A1(n_1959),
.A2(n_541),
.B(n_507),
.C(n_1357),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1972),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1962),
.B(n_5),
.Y(n_2132)
);

AOI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2031),
.A2(n_659),
.B1(n_662),
.B2(n_655),
.C(n_652),
.Y(n_2133)
);

OR2x6_ASAP7_75t_L g2134 ( 
.A(n_1947),
.B(n_1367),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1974),
.A2(n_664),
.B1(n_665),
.B2(n_663),
.Y(n_2135)
);

AOI221xp5_ASAP7_75t_L g2136 ( 
.A1(n_1954),
.A2(n_674),
.B1(n_675),
.B2(n_673),
.C(n_669),
.Y(n_2136)
);

AOI21xp33_ASAP7_75t_L g2137 ( 
.A1(n_2015),
.A2(n_680),
.B(n_679),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1940),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1942),
.Y(n_2139)
);

AOI33xp33_ASAP7_75t_L g2140 ( 
.A1(n_1963),
.A2(n_685),
.A3(n_682),
.B1(n_688),
.B2(n_683),
.B3(n_681),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_1954),
.A2(n_1426),
.B1(n_522),
.B2(n_566),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2035),
.A2(n_882),
.B1(n_886),
.B2(n_872),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_2018),
.Y(n_2143)
);

CKINVDCx20_ASAP7_75t_R g2144 ( 
.A(n_1967),
.Y(n_2144)
);

AOI221xp5_ASAP7_75t_L g2145 ( 
.A1(n_1953),
.A2(n_566),
.B1(n_522),
.B2(n_452),
.C(n_406),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_1965),
.Y(n_2146)
);

OAI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_2044),
.A2(n_522),
.B1(n_566),
.B2(n_452),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1966),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2035),
.A2(n_886),
.B1(n_882),
.B2(n_1198),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_2041),
.Y(n_2150)
);

OAI221xp5_ASAP7_75t_SL g2151 ( 
.A1(n_1929),
.A2(n_1279),
.B1(n_1205),
.B2(n_1210),
.C(n_1161),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1987),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1987),
.B(n_5),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_2023),
.B(n_6),
.Y(n_2154)
);

OAI221xp5_ASAP7_75t_L g2155 ( 
.A1(n_1970),
.A2(n_1279),
.B1(n_566),
.B2(n_522),
.C(n_1161),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_SL g2156 ( 
.A1(n_1914),
.A2(n_566),
.B1(n_522),
.B2(n_394),
.Y(n_2156)
);

AO31x2_ASAP7_75t_L g2157 ( 
.A1(n_1916),
.A2(n_894),
.A3(n_891),
.B(n_1421),
.Y(n_2157)
);

AOI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_1971),
.A2(n_1938),
.B(n_2011),
.Y(n_2158)
);

OAI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_2044),
.A2(n_1471),
.B1(n_1469),
.B2(n_1445),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1977),
.A2(n_1222),
.B1(n_1224),
.B2(n_1198),
.Y(n_2160)
);

OR2x6_ASAP7_75t_L g2161 ( 
.A(n_2013),
.B(n_1367),
.Y(n_2161)
);

OAI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_1978),
.A2(n_419),
.B1(n_425),
.B2(n_409),
.C(n_383),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2020),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2010),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_2049),
.B(n_1235),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1969),
.B(n_7),
.Y(n_2166)
);

OAI221xp5_ASAP7_75t_L g2167 ( 
.A1(n_1978),
.A2(n_429),
.B1(n_430),
.B2(n_427),
.C(n_426),
.Y(n_2167)
);

OAI21x1_ASAP7_75t_L g2168 ( 
.A1(n_2020),
.A2(n_1449),
.B(n_1367),
.Y(n_2168)
);

BUFx12f_ASAP7_75t_L g2169 ( 
.A(n_2047),
.Y(n_2169)
);

OA21x2_ASAP7_75t_L g2170 ( 
.A1(n_2041),
.A2(n_999),
.B(n_998),
.Y(n_2170)
);

INVx3_ASAP7_75t_SL g2171 ( 
.A(n_1983),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2016),
.Y(n_2172)
);

AOI221xp5_ASAP7_75t_L g2173 ( 
.A1(n_1995),
.A2(n_2042),
.B1(n_2027),
.B2(n_2039),
.C(n_2052),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2027),
.B(n_7),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1990),
.Y(n_2175)
);

INVxp67_ASAP7_75t_SL g2176 ( 
.A(n_1957),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_L g2177 ( 
.A1(n_2019),
.A2(n_1224),
.B1(n_1225),
.B2(n_1222),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_1971),
.A2(n_1153),
.B(n_1207),
.Y(n_2178)
);

CKINVDCx20_ASAP7_75t_R g2179 ( 
.A(n_2045),
.Y(n_2179)
);

OAI33xp33_ASAP7_75t_L g2180 ( 
.A1(n_2030),
.A2(n_835),
.A3(n_830),
.B1(n_442),
.B2(n_433),
.B3(n_444),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_2047),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_1921),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2019),
.A2(n_1228),
.B1(n_1245),
.B2(n_1225),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_1920),
.A2(n_1949),
.B1(n_2008),
.B2(n_2002),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1994),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2057),
.A2(n_1245),
.B1(n_1254),
.B2(n_1228),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1984),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2025),
.B(n_8),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1957),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2026),
.B(n_9),
.Y(n_2190)
);

AOI21x1_ASAP7_75t_L g2191 ( 
.A1(n_2039),
.A2(n_1120),
.B(n_1012),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_2053),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_1933),
.B(n_10),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_1980),
.A2(n_447),
.B1(n_459),
.B2(n_441),
.C(n_432),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2043),
.A2(n_1257),
.B1(n_1262),
.B2(n_1254),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2001),
.A2(n_1262),
.B1(n_1272),
.B2(n_1257),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_SL g2197 ( 
.A1(n_1955),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2197)
);

OAI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_2032),
.A2(n_1373),
.B1(n_1205),
.B2(n_1210),
.Y(n_2198)
);

CKINVDCx20_ASAP7_75t_R g2199 ( 
.A(n_2033),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1984),
.B(n_11),
.Y(n_2200)
);

AOI221xp5_ASAP7_75t_L g2201 ( 
.A1(n_1980),
.A2(n_474),
.B1(n_478),
.B2(n_466),
.C(n_461),
.Y(n_2201)
);

AOI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_1934),
.A2(n_1935),
.B1(n_1950),
.B2(n_1936),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_L g2203 ( 
.A1(n_1928),
.A2(n_1338),
.B(n_1211),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1984),
.Y(n_2204)
);

AOI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_1958),
.A2(n_1273),
.B1(n_1284),
.B2(n_1272),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2055),
.B(n_12),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_2021),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1930),
.B(n_14),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1982),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_1926),
.A2(n_481),
.B1(n_486),
.B2(n_480),
.C(n_479),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_1955),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2051),
.B(n_14),
.Y(n_2212)
);

OAI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2056),
.A2(n_490),
.B1(n_491),
.B2(n_487),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2187),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_2176),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2150),
.B(n_2054),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2204),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2084),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2084),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2123),
.B(n_2163),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2189),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_2113),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2200),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_2060),
.B(n_1946),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2152),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_2090),
.B(n_1986),
.Y(n_2226)
);

BUFx2_ASAP7_75t_L g2227 ( 
.A(n_2208),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2182),
.B(n_1930),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2063),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2078),
.B(n_2047),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2208),
.B(n_1988),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2200),
.Y(n_2232)
);

INVx4_ASAP7_75t_L g2233 ( 
.A(n_2060),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2068),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2146),
.B(n_1988),
.Y(n_2235)
);

INVx4_ASAP7_75t_L g2236 ( 
.A(n_2060),
.Y(n_2236)
);

AND2x4_ASAP7_75t_SL g2237 ( 
.A(n_2066),
.B(n_1986),
.Y(n_2237)
);

BUFx12f_ASAP7_75t_L g2238 ( 
.A(n_2089),
.Y(n_2238)
);

OAI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2085),
.A2(n_2006),
.B(n_1981),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2076),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2088),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2164),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2152),
.B(n_1986),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2131),
.B(n_1988),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2103),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_2143),
.Y(n_2246)
);

HB1xp67_ASAP7_75t_L g2247 ( 
.A(n_2107),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_2066),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2192),
.B(n_2209),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2172),
.Y(n_2250)
);

OR2x2_ASAP7_75t_L g2251 ( 
.A(n_2116),
.B(n_1928),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2086),
.A2(n_1914),
.B1(n_1926),
.B2(n_2021),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2059),
.B(n_2036),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2211),
.B(n_2036),
.Y(n_2254)
);

INVxp67_ASAP7_75t_SL g2255 ( 
.A(n_2124),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2211),
.B(n_2036),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_2158),
.B(n_1993),
.Y(n_2257)
);

OAI332xp33_ASAP7_75t_L g2258 ( 
.A1(n_2110),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_20),
.B3(n_23),
.C1(n_24),
.C2(n_25),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_SL g2259 ( 
.A(n_2073),
.B(n_2000),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_2179),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2082),
.B(n_1989),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_2077),
.B(n_2207),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_2169),
.Y(n_2263)
);

NOR2x1_ASAP7_75t_L g2264 ( 
.A(n_2104),
.B(n_1153),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2115),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2126),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2138),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2093),
.B(n_1989),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2139),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2061),
.A2(n_1338),
.B1(n_1139),
.B2(n_1233),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2118),
.B(n_1989),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2100),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2148),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2106),
.Y(n_2274)
);

OR2x2_ASAP7_75t_L g2275 ( 
.A(n_2093),
.B(n_2108),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2175),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2185),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2117),
.B(n_1997),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2170),
.Y(n_2279)
);

NAND2x1_ASAP7_75t_L g2280 ( 
.A(n_2106),
.B(n_975),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_2096),
.Y(n_2281)
);

AND2x2_ASAP7_75t_SL g2282 ( 
.A(n_2166),
.B(n_17),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_2124),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2112),
.B(n_1997),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_2083),
.B(n_1997),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2111),
.B(n_18),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2083),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2181),
.B(n_20),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2170),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_2119),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2173),
.B(n_24),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2174),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2134),
.B(n_2166),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2174),
.B(n_28),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2132),
.B(n_28),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2153),
.B(n_29),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2071),
.A2(n_2064),
.B1(n_2069),
.B2(n_2062),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2206),
.B(n_29),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2097),
.B(n_30),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2193),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2064),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2154),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2171),
.B(n_30),
.Y(n_2303)
);

INVx3_ASAP7_75t_L g2304 ( 
.A(n_2104),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2188),
.B(n_2190),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2122),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2157),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2199),
.B(n_31),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2099),
.B(n_31),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_2119),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2212),
.B(n_32),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2122),
.Y(n_2312)
);

INVx2_ASAP7_75t_R g2313 ( 
.A(n_2075),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2157),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2180),
.A2(n_1284),
.B1(n_1293),
.B2(n_1273),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2191),
.Y(n_2316)
);

AOI211xp5_ASAP7_75t_L g2317 ( 
.A1(n_2058),
.A2(n_35),
.B(n_32),
.C(n_34),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2134),
.B(n_34),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_2119),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2129),
.B(n_35),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2129),
.B(n_2079),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2134),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2168),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2157),
.Y(n_2324)
);

CKINVDCx20_ASAP7_75t_R g2325 ( 
.A(n_2101),
.Y(n_2325)
);

HB1xp67_ASAP7_75t_L g2326 ( 
.A(n_2061),
.Y(n_2326)
);

AND2x4_ASAP7_75t_L g2327 ( 
.A(n_2161),
.B(n_36),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2144),
.B(n_37),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_2161),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2067),
.B(n_1235),
.Y(n_2330)
);

BUFx3_ASAP7_75t_L g2331 ( 
.A(n_2197),
.Y(n_2331)
);

AOI21xp33_ASAP7_75t_L g2332 ( 
.A1(n_2098),
.A2(n_38),
.B(n_40),
.Y(n_2332)
);

BUFx2_ASAP7_75t_L g2333 ( 
.A(n_2161),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2165),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2203),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2080),
.B(n_40),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2202),
.B(n_41),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2072),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2159),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2072),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2247),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2234),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_2260),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2310),
.B(n_2114),
.Y(n_2344)
);

INVx2_ASAP7_75t_SL g2345 ( 
.A(n_2260),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2234),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2233),
.Y(n_2347)
);

OAI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2252),
.A2(n_2102),
.B1(n_2094),
.B2(n_2155),
.Y(n_2348)
);

OAI21xp33_ASAP7_75t_SL g2349 ( 
.A1(n_2326),
.A2(n_2109),
.B(n_2210),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2274),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2274),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_2255),
.A2(n_2137),
.B(n_2130),
.Y(n_2352)
);

AOI221x1_ASAP7_75t_L g2353 ( 
.A1(n_2304),
.A2(n_2137),
.B1(n_2178),
.B2(n_2092),
.C(n_2198),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2240),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2240),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2218),
.B(n_2120),
.Y(n_2356)
);

OAI22xp33_ASAP7_75t_L g2357 ( 
.A1(n_2259),
.A2(n_2094),
.B1(n_2135),
.B2(n_2147),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_2233),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2274),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_2238),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2245),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2218),
.B(n_2219),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2339),
.B(n_2184),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2216),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2216),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2233),
.B(n_2127),
.Y(n_2366)
);

NAND4xp25_ASAP7_75t_L g2367 ( 
.A(n_2331),
.B(n_2317),
.C(n_2264),
.D(n_2236),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2219),
.B(n_2140),
.Y(n_2368)
);

AND2x6_ASAP7_75t_L g2369 ( 
.A(n_2303),
.B(n_2213),
.Y(n_2369)
);

OA21x2_ASAP7_75t_L g2370 ( 
.A1(n_2301),
.A2(n_2065),
.B(n_2070),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2283),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2245),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2291),
.A2(n_2141),
.B(n_2092),
.Y(n_2373)
);

OA21x2_ASAP7_75t_L g2374 ( 
.A1(n_2301),
.A2(n_2201),
.B(n_2194),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2285),
.Y(n_2375)
);

OAI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2331),
.A2(n_2156),
.B1(n_2081),
.B2(n_2074),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2285),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2310),
.B(n_2177),
.Y(n_2378)
);

A2O1A1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_2297),
.A2(n_2136),
.B(n_2125),
.C(n_2128),
.Y(n_2379)
);

OAI32xp33_ASAP7_75t_L g2380 ( 
.A1(n_2251),
.A2(n_2198),
.A3(n_2167),
.B1(n_2162),
.B2(n_2087),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2321),
.A2(n_2145),
.B(n_2162),
.Y(n_2381)
);

OAI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2275),
.A2(n_2151),
.B1(n_2167),
.B2(n_2091),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2217),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_2236),
.Y(n_2384)
);

NOR2x1_ASAP7_75t_SL g2385 ( 
.A(n_2290),
.B(n_2183),
.Y(n_2385)
);

OAI21xp33_ASAP7_75t_L g2386 ( 
.A1(n_2228),
.A2(n_2275),
.B(n_2339),
.Y(n_2386)
);

AO31x2_ASAP7_75t_L g2387 ( 
.A1(n_2227),
.A2(n_2205),
.A3(n_2196),
.B(n_1295),
.Y(n_2387)
);

OA21x2_ASAP7_75t_L g2388 ( 
.A1(n_2217),
.A2(n_2095),
.B(n_2186),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2327),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2265),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2312),
.Y(n_2391)
);

OAI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2340),
.A2(n_2133),
.B1(n_2195),
.B2(n_2149),
.Y(n_2392)
);

OA21x2_ASAP7_75t_L g2393 ( 
.A1(n_2214),
.A2(n_2160),
.B(n_2142),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2293),
.B(n_41),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2265),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2266),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2327),
.Y(n_2397)
);

AO31x2_ASAP7_75t_L g2398 ( 
.A1(n_2227),
.A2(n_1295),
.A3(n_1293),
.B(n_835),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2266),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2236),
.B(n_2313),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2330),
.A2(n_2121),
.B(n_2105),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2220),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2229),
.Y(n_2403)
);

OAI21xp33_ASAP7_75t_SL g2404 ( 
.A1(n_2308),
.A2(n_42),
.B(n_43),
.Y(n_2404)
);

OAI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_2282),
.A2(n_1139),
.B(n_494),
.Y(n_2405)
);

A2O1A1Ixp33_ASAP7_75t_L g2406 ( 
.A1(n_2223),
.A2(n_495),
.B(n_496),
.C(n_492),
.Y(n_2406)
);

BUFx2_ASAP7_75t_L g2407 ( 
.A(n_2304),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2267),
.Y(n_2408)
);

OAI211xp5_ASAP7_75t_SL g2409 ( 
.A1(n_2302),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_2409)
);

INVxp67_ASAP7_75t_SL g2410 ( 
.A(n_2334),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_2248),
.Y(n_2411)
);

INVxp67_ASAP7_75t_SL g2412 ( 
.A(n_2244),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2292),
.B(n_44),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2269),
.Y(n_2414)
);

INVxp67_ASAP7_75t_L g2415 ( 
.A(n_2222),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2310),
.B(n_46),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2262),
.B(n_1147),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2327),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2231),
.A2(n_1207),
.B(n_1200),
.Y(n_2419)
);

AOI221xp5_ASAP7_75t_L g2420 ( 
.A1(n_2223),
.A2(n_502),
.B1(n_519),
.B2(n_500),
.C(n_497),
.Y(n_2420)
);

AOI222xp33_ASAP7_75t_L g2421 ( 
.A1(n_2306),
.A2(n_523),
.B1(n_535),
.B2(n_547),
.C1(n_555),
.C2(n_556),
.Y(n_2421)
);

O2A1O1Ixp5_ASAP7_75t_L g2422 ( 
.A1(n_2257),
.A2(n_1211),
.B(n_1220),
.C(n_1200),
.Y(n_2422)
);

BUFx2_ASAP7_75t_L g2423 ( 
.A(n_2304),
.Y(n_2423)
);

AO21x2_ASAP7_75t_L g2424 ( 
.A1(n_2286),
.A2(n_1220),
.B(n_1012),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2273),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2232),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2292),
.B(n_46),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2273),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2232),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2248),
.B(n_48),
.Y(n_2430)
);

OAI21x1_ASAP7_75t_L g2431 ( 
.A1(n_2248),
.A2(n_1338),
.B(n_1439),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2313),
.B(n_48),
.Y(n_2432)
);

OAI21x1_ASAP7_75t_L g2433 ( 
.A1(n_2225),
.A2(n_2251),
.B(n_2214),
.Y(n_2433)
);

INVx2_ASAP7_75t_R g2434 ( 
.A(n_2323),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2338),
.A2(n_1018),
.B1(n_1020),
.B2(n_998),
.Y(n_2435)
);

OA21x2_ASAP7_75t_L g2436 ( 
.A1(n_2262),
.A2(n_2215),
.B(n_2257),
.Y(n_2436)
);

AOI211xp5_ASAP7_75t_L g2437 ( 
.A1(n_2258),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_2437)
);

INVxp67_ASAP7_75t_L g2438 ( 
.A(n_2306),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2276),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2238),
.B(n_50),
.Y(n_2440)
);

AO31x2_ASAP7_75t_L g2441 ( 
.A1(n_2268),
.A2(n_830),
.A3(n_1020),
.B(n_1018),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2276),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2277),
.Y(n_2443)
);

AOI21x1_ASAP7_75t_L g2444 ( 
.A1(n_2262),
.A2(n_976),
.B(n_975),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2277),
.Y(n_2445)
);

A2O1A1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2320),
.A2(n_560),
.B(n_562),
.C(n_559),
.Y(n_2446)
);

NAND2x1_ASAP7_75t_L g2447 ( 
.A(n_2215),
.B(n_976),
.Y(n_2447)
);

AOI21xp33_ASAP7_75t_L g2448 ( 
.A1(n_2320),
.A2(n_53),
.B(n_55),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2282),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2246),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2241),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_2300),
.B(n_57),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2300),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2453),
.B(n_2221),
.Y(n_2454)
);

OAI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2437),
.A2(n_2293),
.B1(n_2319),
.B2(n_2290),
.Y(n_2455)
);

AOI22xp33_ASAP7_75t_L g2456 ( 
.A1(n_2374),
.A2(n_2370),
.B1(n_2369),
.B2(n_2386),
.Y(n_2456)
);

OAI211xp5_ASAP7_75t_SL g2457 ( 
.A1(n_2437),
.A2(n_2294),
.B(n_2296),
.C(n_2263),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2342),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_2345),
.Y(n_2459)
);

AOI33xp33_ASAP7_75t_L g2460 ( 
.A1(n_2402),
.A2(n_2328),
.A3(n_2308),
.B1(n_2299),
.B2(n_2311),
.B3(n_2288),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2346),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2343),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2354),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2436),
.Y(n_2464)
);

OR2x6_ASAP7_75t_L g2465 ( 
.A(n_2352),
.B(n_2337),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2436),
.B(n_2249),
.Y(n_2466)
);

HB1xp67_ASAP7_75t_L g2467 ( 
.A(n_2364),
.Y(n_2467)
);

INVxp67_ASAP7_75t_SL g2468 ( 
.A(n_2385),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2410),
.B(n_2249),
.Y(n_2469)
);

INVx4_ASAP7_75t_L g2470 ( 
.A(n_2360),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2355),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2411),
.Y(n_2472)
);

AO21x2_ASAP7_75t_L g2473 ( 
.A1(n_2386),
.A2(n_2337),
.B(n_2328),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2347),
.Y(n_2474)
);

HB1xp67_ASAP7_75t_L g2475 ( 
.A(n_2365),
.Y(n_2475)
);

OAI211xp5_ASAP7_75t_L g2476 ( 
.A1(n_2349),
.A2(n_2353),
.B(n_2367),
.C(n_2404),
.Y(n_2476)
);

OR2x2_ASAP7_75t_L g2477 ( 
.A(n_2391),
.B(n_2221),
.Y(n_2477)
);

OAI221xp5_ASAP7_75t_SL g2478 ( 
.A1(n_2349),
.A2(n_2318),
.B1(n_2299),
.B2(n_2253),
.C(n_2338),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_2374),
.A2(n_2253),
.B1(n_2340),
.B2(n_2261),
.Y(n_2479)
);

OAI221xp5_ASAP7_75t_L g2480 ( 
.A1(n_2404),
.A2(n_2239),
.B1(n_2235),
.B2(n_2333),
.C(n_2329),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2358),
.B(n_2230),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2350),
.B(n_2351),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2433),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2356),
.A2(n_2293),
.B1(n_2319),
.B2(n_2280),
.Y(n_2484)
);

BUFx2_ASAP7_75t_SL g2485 ( 
.A(n_2394),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2369),
.B(n_2309),
.Y(n_2486)
);

AOI22xp33_ASAP7_75t_L g2487 ( 
.A1(n_2370),
.A2(n_2261),
.B1(n_2316),
.B2(n_2257),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2359),
.B(n_2230),
.Y(n_2488)
);

OR2x2_ASAP7_75t_L g2489 ( 
.A(n_2356),
.B(n_2287),
.Y(n_2489)
);

OR2x6_ASAP7_75t_L g2490 ( 
.A(n_2449),
.B(n_2318),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2411),
.B(n_2287),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2361),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2430),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2425),
.Y(n_2494)
);

OAI22xp5_ASAP7_75t_L g2495 ( 
.A1(n_2415),
.A2(n_2280),
.B1(n_2226),
.B2(n_2224),
.Y(n_2495)
);

BUFx2_ASAP7_75t_L g2496 ( 
.A(n_2384),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2369),
.B(n_2309),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2369),
.B(n_2295),
.Y(n_2498)
);

INVx2_ASAP7_75t_SL g2499 ( 
.A(n_2384),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_2371),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2372),
.Y(n_2501)
);

NAND3xp33_ASAP7_75t_L g2502 ( 
.A(n_2373),
.B(n_2323),
.C(n_2316),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2428),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2442),
.Y(n_2504)
);

OAI21xp5_ASAP7_75t_SL g2505 ( 
.A1(n_2367),
.A2(n_2303),
.B(n_2288),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2407),
.B(n_2225),
.Y(n_2506)
);

OAI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2444),
.A2(n_2225),
.B(n_2335),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2423),
.B(n_2263),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2368),
.B(n_2295),
.Y(n_2509)
);

OR2x6_ASAP7_75t_L g2510 ( 
.A(n_2449),
.B(n_2281),
.Y(n_2510)
);

HB1xp67_ASAP7_75t_L g2511 ( 
.A(n_2450),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2363),
.A2(n_2357),
.B1(n_2348),
.B2(n_2381),
.Y(n_2512)
);

INVx1_ASAP7_75t_SL g2513 ( 
.A(n_2394),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2445),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2390),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2452),
.Y(n_2516)
);

HB1xp67_ASAP7_75t_L g2517 ( 
.A(n_2438),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2400),
.B(n_2263),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2395),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2341),
.B(n_2243),
.Y(n_2520)
);

HB1xp67_ASAP7_75t_L g2521 ( 
.A(n_2403),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2396),
.Y(n_2522)
);

INVx2_ASAP7_75t_SL g2523 ( 
.A(n_2344),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2378),
.B(n_2243),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2426),
.B(n_2429),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2399),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_2447),
.Y(n_2527)
);

AND2x4_ASAP7_75t_L g2528 ( 
.A(n_2408),
.B(n_2279),
.Y(n_2528)
);

AND2x2_ASAP7_75t_SL g2529 ( 
.A(n_2432),
.B(n_2281),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2414),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2368),
.B(n_2279),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2413),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_SL g2533 ( 
.A1(n_2379),
.A2(n_2311),
.B(n_2298),
.Y(n_2533)
);

OAI221xp5_ASAP7_75t_SL g2534 ( 
.A1(n_2446),
.A2(n_2298),
.B1(n_2333),
.B2(n_2329),
.C(n_2305),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2383),
.Y(n_2535)
);

HB1xp67_ASAP7_75t_L g2536 ( 
.A(n_2413),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_2416),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2434),
.B(n_2305),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2389),
.B(n_2271),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2427),
.B(n_2271),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2427),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2523),
.B(n_2397),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2462),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2509),
.B(n_2362),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2521),
.Y(n_2545)
);

AND2x4_ASAP7_75t_SL g2546 ( 
.A(n_2508),
.B(n_2325),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2473),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2538),
.B(n_2362),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2538),
.B(n_2366),
.Y(n_2549)
);

INVx2_ASAP7_75t_SL g2550 ( 
.A(n_2518),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2511),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2536),
.B(n_2439),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2460),
.B(n_2418),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2485),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2518),
.B(n_2443),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2508),
.B(n_2412),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2473),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2473),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2476),
.B(n_2448),
.Y(n_2559)
);

HB1xp67_ASAP7_75t_L g2560 ( 
.A(n_2459),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2460),
.B(n_2448),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2458),
.Y(n_2562)
);

INVxp67_ASAP7_75t_SL g2563 ( 
.A(n_2464),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2464),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2523),
.B(n_2382),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2532),
.B(n_2375),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2464),
.Y(n_2567)
);

BUFx3_ASAP7_75t_L g2568 ( 
.A(n_2470),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2493),
.B(n_2537),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2481),
.B(n_2440),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2510),
.Y(n_2571)
);

HB1xp67_ASAP7_75t_L g2572 ( 
.A(n_2459),
.Y(n_2572)
);

OR2x2_ASAP7_75t_L g2573 ( 
.A(n_2541),
.B(n_2531),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2461),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2463),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2481),
.B(n_2377),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2466),
.B(n_2226),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2471),
.Y(n_2578)
);

OR2x2_ASAP7_75t_L g2579 ( 
.A(n_2531),
.B(n_2454),
.Y(n_2579)
);

NAND3xp33_ASAP7_75t_L g2580 ( 
.A(n_2502),
.B(n_2382),
.C(n_2409),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2493),
.B(n_2537),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2469),
.B(n_2289),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2466),
.B(n_2226),
.Y(n_2583)
);

NAND5xp2_ASAP7_75t_L g2584 ( 
.A(n_2505),
.B(n_2405),
.C(n_2421),
.D(n_2401),
.E(n_2420),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2516),
.B(n_2380),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2490),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2488),
.B(n_2520),
.Y(n_2587)
);

OR2x2_ASAP7_75t_L g2588 ( 
.A(n_2489),
.B(n_2289),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2488),
.B(n_2237),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2520),
.B(n_2237),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2454),
.B(n_2424),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2490),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2470),
.B(n_2325),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2468),
.B(n_2278),
.Y(n_2594)
);

AND2x2_ASAP7_75t_SL g2595 ( 
.A(n_2456),
.B(n_2281),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2506),
.B(n_2278),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2492),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2501),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2506),
.B(n_2417),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2482),
.B(n_2281),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2515),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2490),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2482),
.B(n_2281),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2474),
.B(n_2322),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2516),
.B(n_2421),
.Y(n_2605)
);

AND2x4_ASAP7_75t_SL g2606 ( 
.A(n_2470),
.B(n_2467),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2513),
.B(n_2376),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2496),
.B(n_2475),
.Y(n_2608)
);

AND2x4_ASAP7_75t_L g2609 ( 
.A(n_2510),
.B(n_2424),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2519),
.Y(n_2610)
);

AOI21xp33_ASAP7_75t_L g2611 ( 
.A1(n_2465),
.A2(n_2376),
.B(n_2422),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2517),
.B(n_2284),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2490),
.B(n_2284),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2529),
.B(n_2336),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2489),
.B(n_2392),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2465),
.B(n_2406),
.Y(n_2616)
);

HB1xp67_ASAP7_75t_L g2617 ( 
.A(n_2500),
.Y(n_2617)
);

INVxp67_ASAP7_75t_SL g2618 ( 
.A(n_2498),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2510),
.Y(n_2619)
);

INVx2_ASAP7_75t_SL g2620 ( 
.A(n_2472),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2499),
.B(n_2322),
.Y(n_2621)
);

OR2x6_ASAP7_75t_L g2622 ( 
.A(n_2533),
.B(n_2405),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2477),
.B(n_2451),
.Y(n_2623)
);

NAND4xp75_ASAP7_75t_SL g2624 ( 
.A(n_2549),
.B(n_2491),
.C(n_2524),
.D(n_2539),
.Y(n_2624)
);

INVx4_ASAP7_75t_L g2625 ( 
.A(n_2568),
.Y(n_2625)
);

AOI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2559),
.A2(n_2465),
.B1(n_2457),
.B2(n_2510),
.Y(n_2626)
);

NAND4xp75_ASAP7_75t_SL g2627 ( 
.A(n_2549),
.B(n_2491),
.C(n_2524),
.D(n_2539),
.Y(n_2627)
);

XNOR2xp5_ASAP7_75t_L g2628 ( 
.A(n_2570),
.B(n_2529),
.Y(n_2628)
);

NAND4xp75_ASAP7_75t_SL g2629 ( 
.A(n_2594),
.B(n_2534),
.C(n_2484),
.D(n_2455),
.Y(n_2629)
);

XNOR2xp5_ASAP7_75t_L g2630 ( 
.A(n_2570),
.B(n_2512),
.Y(n_2630)
);

NAND4xp75_ASAP7_75t_L g2631 ( 
.A(n_2559),
.B(n_2486),
.C(n_2497),
.D(n_2483),
.Y(n_2631)
);

INVx2_ASAP7_75t_SL g2632 ( 
.A(n_2546),
.Y(n_2632)
);

XNOR2xp5_ASAP7_75t_L g2633 ( 
.A(n_2546),
.B(n_2465),
.Y(n_2633)
);

AND2x4_ASAP7_75t_SL g2634 ( 
.A(n_2593),
.B(n_2472),
.Y(n_2634)
);

NAND4xp75_ASAP7_75t_L g2635 ( 
.A(n_2595),
.B(n_2483),
.C(n_2540),
.D(n_2535),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2587),
.B(n_2533),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2587),
.B(n_2499),
.Y(n_2637)
);

AO22x2_ASAP7_75t_L g2638 ( 
.A1(n_2547),
.A2(n_2530),
.B1(n_2535),
.B2(n_2526),
.Y(n_2638)
);

NAND2xp33_ASAP7_75t_R g2639 ( 
.A(n_2622),
.B(n_2472),
.Y(n_2639)
);

INVxp67_ASAP7_75t_L g2640 ( 
.A(n_2560),
.Y(n_2640)
);

BUFx2_ASAP7_75t_L g2641 ( 
.A(n_2542),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2571),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_2568),
.B(n_2480),
.Y(n_2643)
);

AOI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2580),
.A2(n_2479),
.B1(n_2487),
.B2(n_2388),
.Y(n_2644)
);

NOR2x1_ASAP7_75t_L g2645 ( 
.A(n_2616),
.B(n_2522),
.Y(n_2645)
);

NOR3xp33_ASAP7_75t_L g2646 ( 
.A(n_2611),
.B(n_2478),
.C(n_2495),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2622),
.A2(n_2388),
.B1(n_2336),
.B2(n_2528),
.Y(n_2647)
);

INVx1_ASAP7_75t_SL g2648 ( 
.A(n_2606),
.Y(n_2648)
);

INVxp67_ASAP7_75t_SL g2649 ( 
.A(n_2571),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2617),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2579),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2576),
.B(n_2525),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_SL g2653 ( 
.A1(n_2561),
.A2(n_2477),
.B1(n_2525),
.B2(n_2528),
.Y(n_2653)
);

NOR2x1_ASAP7_75t_L g2654 ( 
.A(n_2565),
.B(n_2525),
.Y(n_2654)
);

XOR2x2_ASAP7_75t_L g2655 ( 
.A(n_2615),
.B(n_2336),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2571),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2606),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2579),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2564),
.Y(n_2659)
);

NAND3xp33_ASAP7_75t_SL g2660 ( 
.A(n_2554),
.B(n_2503),
.C(n_2494),
.Y(n_2660)
);

AOI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2622),
.A2(n_2528),
.B1(n_2332),
.B2(n_2503),
.Y(n_2661)
);

XOR2x2_ASAP7_75t_L g2662 ( 
.A(n_2607),
.B(n_2393),
.Y(n_2662)
);

NOR3xp33_ASAP7_75t_SL g2663 ( 
.A(n_2618),
.B(n_2270),
.C(n_2507),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2564),
.Y(n_2664)
);

OAI31xp33_ASAP7_75t_L g2665 ( 
.A1(n_2584),
.A2(n_2494),
.A3(n_2514),
.B(n_2504),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2542),
.B(n_2527),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2552),
.Y(n_2667)
);

NOR2x1_ASAP7_75t_L g2668 ( 
.A(n_2567),
.B(n_2527),
.Y(n_2668)
);

OR2x2_ASAP7_75t_L g2669 ( 
.A(n_2553),
.B(n_2504),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2576),
.B(n_2527),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2573),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2567),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2544),
.B(n_2514),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2572),
.Y(n_2674)
);

INVx1_ASAP7_75t_SL g2675 ( 
.A(n_2595),
.Y(n_2675)
);

AND2x4_ASAP7_75t_SL g2676 ( 
.A(n_2590),
.B(n_2322),
.Y(n_2676)
);

NAND4xp75_ASAP7_75t_SL g2677 ( 
.A(n_2594),
.B(n_2507),
.C(n_2256),
.D(n_2254),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2567),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2542),
.B(n_2254),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2577),
.Y(n_2680)
);

OR2x2_ASAP7_75t_L g2681 ( 
.A(n_2543),
.B(n_2441),
.Y(n_2681)
);

INVx3_ASAP7_75t_SL g2682 ( 
.A(n_2550),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2577),
.Y(n_2683)
);

OAI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2622),
.A2(n_2435),
.B1(n_2256),
.B2(n_2335),
.Y(n_2684)
);

NAND4xp75_ASAP7_75t_L g2685 ( 
.A(n_2585),
.B(n_2419),
.C(n_2393),
.D(n_2307),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2638),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2641),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2652),
.B(n_2608),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2670),
.B(n_2608),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2637),
.B(n_2590),
.Y(n_2690)
);

NAND4xp25_ASAP7_75t_L g2691 ( 
.A(n_2643),
.B(n_2551),
.C(n_2545),
.D(n_2556),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2674),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2632),
.B(n_2550),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2638),
.Y(n_2694)
);

OAI322xp33_ASAP7_75t_L g2695 ( 
.A1(n_2626),
.A2(n_2547),
.A3(n_2558),
.B1(n_2557),
.B2(n_2573),
.C1(n_2586),
.C2(n_2592),
.Y(n_2695)
);

AOI21xp33_ASAP7_75t_L g2696 ( 
.A1(n_2665),
.A2(n_2605),
.B(n_2592),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2649),
.B(n_2556),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_R g2698 ( 
.A(n_2625),
.B(n_2620),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2682),
.B(n_2654),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2673),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2651),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2654),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2680),
.B(n_2548),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2683),
.B(n_2548),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2635),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2658),
.B(n_2671),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2645),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2659),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2648),
.B(n_2604),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2666),
.B(n_2604),
.Y(n_2710)
);

AND2x4_ASAP7_75t_L g2711 ( 
.A(n_2666),
.B(n_2586),
.Y(n_2711)
);

INVx2_ASAP7_75t_SL g2712 ( 
.A(n_2634),
.Y(n_2712)
);

OAI21xp33_ASAP7_75t_L g2713 ( 
.A1(n_2646),
.A2(n_2612),
.B(n_2613),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2644),
.A2(n_2558),
.B1(n_2557),
.B2(n_2614),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2645),
.B(n_2602),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2664),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2657),
.B(n_2589),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2676),
.B(n_2589),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2626),
.B(n_2602),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2640),
.B(n_2555),
.Y(n_2720)
);

AND2x4_ASAP7_75t_L g2721 ( 
.A(n_2625),
.B(n_2619),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2633),
.B(n_2555),
.Y(n_2722)
);

CKINVDCx16_ASAP7_75t_R g2723 ( 
.A(n_2630),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2650),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2642),
.B(n_2569),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2656),
.B(n_2581),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2655),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2667),
.Y(n_2728)
);

INVx1_ASAP7_75t_SL g2729 ( 
.A(n_2636),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2672),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2678),
.Y(n_2731)
);

INVxp67_ASAP7_75t_L g2732 ( 
.A(n_2639),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2707),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2707),
.Y(n_2734)
);

XNOR2xp5_ASAP7_75t_L g2735 ( 
.A(n_2688),
.B(n_2628),
.Y(n_2735)
);

AOI31xp33_ASAP7_75t_L g2736 ( 
.A1(n_2712),
.A2(n_2660),
.A3(n_2669),
.B(n_2563),
.Y(n_2736)
);

AOI21xp33_ASAP7_75t_L g2737 ( 
.A1(n_2705),
.A2(n_2675),
.B(n_2661),
.Y(n_2737)
);

AOI31xp33_ASAP7_75t_L g2738 ( 
.A1(n_2699),
.A2(n_2692),
.A3(n_2712),
.B(n_2687),
.Y(n_2738)
);

NAND3xp33_ASAP7_75t_L g2739 ( 
.A(n_2705),
.B(n_2661),
.C(n_2663),
.Y(n_2739)
);

OAI211xp5_ASAP7_75t_SL g2740 ( 
.A1(n_2713),
.A2(n_2644),
.B(n_2629),
.C(n_2668),
.Y(n_2740)
);

OAI21xp33_ASAP7_75t_L g2741 ( 
.A1(n_2709),
.A2(n_2621),
.B(n_2599),
.Y(n_2741)
);

AOI31xp33_ASAP7_75t_L g2742 ( 
.A1(n_2699),
.A2(n_2668),
.A3(n_2620),
.B(n_2574),
.Y(n_2742)
);

OAI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2714),
.A2(n_2647),
.B1(n_2614),
.B2(n_2588),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2703),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2690),
.Y(n_2745)
);

INVxp67_ASAP7_75t_SL g2746 ( 
.A(n_2697),
.Y(n_2746)
);

NAND3xp33_ASAP7_75t_L g2747 ( 
.A(n_2732),
.B(n_2702),
.C(n_2694),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2689),
.B(n_2631),
.Y(n_2748)
);

OAI22xp33_ASAP7_75t_R g2749 ( 
.A1(n_2706),
.A2(n_2627),
.B1(n_2624),
.B2(n_2653),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2703),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2695),
.A2(n_2662),
.B(n_2647),
.Y(n_2751)
);

INVxp67_ASAP7_75t_L g2752 ( 
.A(n_2709),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2704),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_2718),
.B(n_2619),
.Y(n_2754)
);

XNOR2xp5_ASAP7_75t_L g2755 ( 
.A(n_2688),
.B(n_2685),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2689),
.B(n_2596),
.Y(n_2756)
);

AOI21xp33_ASAP7_75t_L g2757 ( 
.A1(n_2719),
.A2(n_2681),
.B(n_2684),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2723),
.A2(n_2583),
.B1(n_2599),
.B2(n_2600),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2690),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2704),
.Y(n_2760)
);

INVx1_ASAP7_75t_SL g2761 ( 
.A(n_2698),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2693),
.B(n_2566),
.Y(n_2762)
);

NOR2xp33_ASAP7_75t_L g2763 ( 
.A(n_2718),
.B(n_2600),
.Y(n_2763)
);

OAI22xp33_ASAP7_75t_L g2764 ( 
.A1(n_2686),
.A2(n_2582),
.B1(n_2623),
.B2(n_2583),
.Y(n_2764)
);

OAI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2702),
.A2(n_2603),
.B1(n_2596),
.B2(n_2679),
.Y(n_2765)
);

BUFx2_ASAP7_75t_L g2766 ( 
.A(n_2698),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2706),
.B(n_2562),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2686),
.A2(n_2603),
.B1(n_2623),
.B2(n_2679),
.Y(n_2768)
);

AOI21xp33_ASAP7_75t_SL g2769 ( 
.A1(n_2720),
.A2(n_2578),
.B(n_2575),
.Y(n_2769)
);

AOI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2696),
.A2(n_2729),
.B1(n_2700),
.B2(n_2727),
.Y(n_2770)
);

OAI32xp33_ASAP7_75t_L g2771 ( 
.A1(n_2740),
.A2(n_2715),
.A3(n_2691),
.B1(n_2701),
.B2(n_2725),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2756),
.B(n_2693),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2751),
.A2(n_2727),
.B1(n_2711),
.B2(n_2722),
.Y(n_2773)
);

NAND2xp33_ASAP7_75t_SL g2774 ( 
.A(n_2735),
.B(n_2710),
.Y(n_2774)
);

OAI31xp33_ASAP7_75t_L g2775 ( 
.A1(n_2743),
.A2(n_2708),
.A3(n_2716),
.B(n_2711),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2745),
.Y(n_2776)
);

INVx1_ASAP7_75t_SL g2777 ( 
.A(n_2762),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2741),
.B(n_2710),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2761),
.B(n_2693),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2761),
.B(n_2721),
.Y(n_2780)
);

XNOR2xp5_ASAP7_75t_L g2781 ( 
.A(n_2755),
.B(n_2717),
.Y(n_2781)
);

AOI21xp33_ASAP7_75t_L g2782 ( 
.A1(n_2736),
.A2(n_2726),
.B(n_2711),
.Y(n_2782)
);

INVxp67_ASAP7_75t_SL g2783 ( 
.A(n_2752),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2759),
.B(n_2721),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2748),
.A2(n_2728),
.B1(n_2724),
.B2(n_2722),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2758),
.B(n_2721),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2744),
.B(n_2717),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2739),
.A2(n_2609),
.B1(n_2591),
.B2(n_2730),
.Y(n_2788)
);

INVxp67_ASAP7_75t_L g2789 ( 
.A(n_2754),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2750),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2764),
.A2(n_2731),
.B1(n_2621),
.B2(n_2609),
.Y(n_2791)
);

INVx1_ASAP7_75t_SL g2792 ( 
.A(n_2766),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2770),
.A2(n_2747),
.B1(n_2737),
.B2(n_2768),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2742),
.B(n_2598),
.C(n_2597),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2753),
.Y(n_2795)
);

OR2x2_ASAP7_75t_L g2796 ( 
.A(n_2760),
.B(n_2767),
.Y(n_2796)
);

AOI221xp5_ASAP7_75t_L g2797 ( 
.A1(n_2757),
.A2(n_2601),
.B1(n_2610),
.B2(n_2609),
.C(n_2591),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2738),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2738),
.Y(n_2799)
);

OAI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2742),
.A2(n_2677),
.B(n_2431),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2733),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2746),
.B(n_2441),
.Y(n_2802)
);

OAI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_2793),
.A2(n_2763),
.B(n_2765),
.Y(n_2803)
);

AOI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2773),
.A2(n_2749),
.B1(n_2734),
.B2(n_2307),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2781),
.A2(n_2777),
.B1(n_2786),
.B2(n_2791),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2787),
.Y(n_2806)
);

AOI221xp5_ASAP7_75t_L g2807 ( 
.A1(n_2797),
.A2(n_2769),
.B1(n_2272),
.B2(n_2250),
.C(n_2242),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2772),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2784),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2779),
.B(n_2441),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2780),
.B(n_2398),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2796),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2776),
.A2(n_2272),
.B1(n_2241),
.B2(n_2250),
.Y(n_2813)
);

INVxp67_ASAP7_75t_L g2814 ( 
.A(n_2774),
.Y(n_2814)
);

AOI321xp33_ASAP7_75t_L g2815 ( 
.A1(n_2771),
.A2(n_2785),
.A3(n_2788),
.B1(n_2799),
.B2(n_2798),
.C(n_2782),
.Y(n_2815)
);

OR2x2_ASAP7_75t_L g2816 ( 
.A(n_2792),
.B(n_2398),
.Y(n_2816)
);

INVx1_ASAP7_75t_SL g2817 ( 
.A(n_2790),
.Y(n_2817)
);

AOI21xp33_ASAP7_75t_SL g2818 ( 
.A1(n_2775),
.A2(n_59),
.B(n_60),
.Y(n_2818)
);

AOI22xp33_ASAP7_75t_L g2819 ( 
.A1(n_2789),
.A2(n_2802),
.B1(n_2785),
.B2(n_2800),
.Y(n_2819)
);

NAND3xp33_ASAP7_75t_L g2820 ( 
.A(n_2778),
.B(n_2315),
.C(n_2314),
.Y(n_2820)
);

A2O1A1Ixp33_ASAP7_75t_SL g2821 ( 
.A1(n_2801),
.A2(n_2783),
.B(n_2795),
.C(n_2800),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2794),
.B(n_60),
.Y(n_2822)
);

AOI22xp33_ASAP7_75t_L g2823 ( 
.A1(n_2793),
.A2(n_2314),
.B1(n_2324),
.B2(n_2242),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2787),
.Y(n_2824)
);

OAI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2781),
.A2(n_2324),
.B1(n_2398),
.B2(n_2387),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2787),
.B(n_2387),
.Y(n_2826)
);

O2A1O1Ixp33_ASAP7_75t_SL g2827 ( 
.A1(n_2772),
.A2(n_66),
.B(n_62),
.C(n_65),
.Y(n_2827)
);

NAND3xp33_ASAP7_75t_L g2828 ( 
.A(n_2815),
.B(n_568),
.C(n_565),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2808),
.B(n_2387),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2806),
.B(n_62),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2824),
.B(n_65),
.Y(n_2831)
);

INVx1_ASAP7_75t_SL g2832 ( 
.A(n_2817),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2814),
.B(n_66),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2812),
.Y(n_2834)
);

INVx1_ASAP7_75t_SL g2835 ( 
.A(n_2809),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2814),
.B(n_68),
.Y(n_2836)
);

NAND4xp25_ASAP7_75t_L g2837 ( 
.A(n_2804),
.B(n_72),
.C(n_69),
.D(n_71),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2827),
.B(n_73),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2819),
.A2(n_2805),
.B1(n_2822),
.B2(n_2803),
.Y(n_2839)
);

AOI221xp5_ASAP7_75t_L g2840 ( 
.A1(n_2821),
.A2(n_575),
.B1(n_585),
.B2(n_574),
.C(n_571),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_2818),
.B(n_2816),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_SL g2842 ( 
.A(n_2810),
.B(n_1285),
.Y(n_2842)
);

NAND3xp33_ASAP7_75t_L g2843 ( 
.A(n_2811),
.B(n_593),
.C(n_587),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2826),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2820),
.Y(n_2845)
);

NAND2x1p5_ASAP7_75t_L g2846 ( 
.A(n_2807),
.B(n_1266),
.Y(n_2846)
);

AOI321xp33_ASAP7_75t_L g2847 ( 
.A1(n_2839),
.A2(n_2823),
.A3(n_2807),
.B1(n_2825),
.B2(n_2813),
.C(n_1236),
.Y(n_2847)
);

AOI221xp5_ASAP7_75t_L g2848 ( 
.A1(n_2828),
.A2(n_606),
.B1(n_610),
.B2(n_605),
.C(n_595),
.Y(n_2848)
);

NAND3xp33_ASAP7_75t_SL g2849 ( 
.A(n_2832),
.B(n_2835),
.C(n_2838),
.Y(n_2849)
);

OAI21xp5_ASAP7_75t_SL g2850 ( 
.A1(n_2836),
.A2(n_2834),
.B(n_2833),
.Y(n_2850)
);

AOI221x1_ASAP7_75t_L g2851 ( 
.A1(n_2837),
.A2(n_76),
.B1(n_73),
.B2(n_74),
.C(n_78),
.Y(n_2851)
);

AOI221xp5_ASAP7_75t_L g2852 ( 
.A1(n_2841),
.A2(n_621),
.B1(n_625),
.B2(n_618),
.C(n_615),
.Y(n_2852)
);

OAI211xp5_ASAP7_75t_L g2853 ( 
.A1(n_2830),
.A2(n_80),
.B(n_74),
.C(n_78),
.Y(n_2853)
);

O2A1O1Ixp33_ASAP7_75t_L g2854 ( 
.A1(n_2844),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2854)
);

OAI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2840),
.A2(n_1281),
.B1(n_1318),
.B2(n_1303),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2831),
.B(n_2842),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2845),
.A2(n_1281),
.B1(n_1287),
.B2(n_1280),
.Y(n_2857)
);

AOI211xp5_ASAP7_75t_SL g2858 ( 
.A1(n_2829),
.A2(n_85),
.B(n_82),
.C(n_84),
.Y(n_2858)
);

AOI221x1_ASAP7_75t_L g2859 ( 
.A1(n_2843),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C(n_89),
.Y(n_2859)
);

OAI22x1_ASAP7_75t_L g2860 ( 
.A1(n_2857),
.A2(n_2846),
.B1(n_91),
.B2(n_88),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2849),
.Y(n_2861)
);

NAND4xp75_ASAP7_75t_L g2862 ( 
.A(n_2851),
.B(n_2846),
.C(n_94),
.D(n_90),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2856),
.A2(n_1033),
.B1(n_1036),
.B2(n_1024),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2853),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2852),
.A2(n_1033),
.B1(n_1036),
.B2(n_1024),
.Y(n_2865)
);

INVx1_ASAP7_75t_SL g2866 ( 
.A(n_2855),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2854),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_2850),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2859),
.Y(n_2869)
);

AOI22xp33_ASAP7_75t_L g2870 ( 
.A1(n_2848),
.A2(n_1041),
.B1(n_1043),
.B2(n_1038),
.Y(n_2870)
);

AO22x2_ASAP7_75t_L g2871 ( 
.A1(n_2858),
.A2(n_96),
.B1(n_90),
.B2(n_91),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2847),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2861),
.A2(n_1280),
.B1(n_1287),
.B2(n_1184),
.Y(n_2873)
);

AOI222xp33_ASAP7_75t_L g2874 ( 
.A1(n_2869),
.A2(n_1184),
.B1(n_632),
.B2(n_636),
.C1(n_638),
.C2(n_640),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2871),
.B(n_102),
.Y(n_2875)
);

OAI211xp5_ASAP7_75t_SL g2876 ( 
.A1(n_2864),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_2876)
);

OAI32xp33_ASAP7_75t_L g2877 ( 
.A1(n_2867),
.A2(n_103),
.A3(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_2877)
);

AOI211xp5_ASAP7_75t_SL g2878 ( 
.A1(n_2872),
.A2(n_113),
.B(n_108),
.C(n_112),
.Y(n_2878)
);

A2O1A1Ixp33_ASAP7_75t_L g2879 ( 
.A1(n_2868),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2879)
);

NOR3xp33_ASAP7_75t_L g2880 ( 
.A(n_2862),
.B(n_643),
.C(n_627),
.Y(n_2880)
);

AOI221xp5_ASAP7_75t_L g2881 ( 
.A1(n_2860),
.A2(n_644),
.B1(n_654),
.B2(n_658),
.C(n_667),
.Y(n_2881)
);

OAI211xp5_ASAP7_75t_SL g2882 ( 
.A1(n_2866),
.A2(n_117),
.B(n_114),
.C(n_115),
.Y(n_2882)
);

AOI221xp5_ASAP7_75t_L g2883 ( 
.A1(n_2871),
.A2(n_676),
.B1(n_687),
.B2(n_120),
.C(n_121),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2863),
.B(n_2870),
.Y(n_2884)
);

INVx2_ASAP7_75t_SL g2885 ( 
.A(n_2865),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2861),
.A2(n_1280),
.B1(n_1287),
.B2(n_1184),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2861),
.A2(n_1303),
.B1(n_1318),
.B2(n_1011),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_SL g2888 ( 
.A1(n_2861),
.A2(n_117),
.B(n_119),
.Y(n_2888)
);

AOI211x1_ASAP7_75t_L g2889 ( 
.A1(n_2861),
.A2(n_122),
.B(n_119),
.C(n_121),
.Y(n_2889)
);

AOI211xp5_ASAP7_75t_L g2890 ( 
.A1(n_2888),
.A2(n_125),
.B(n_122),
.C(n_123),
.Y(n_2890)
);

NAND3xp33_ASAP7_75t_L g2891 ( 
.A(n_2880),
.B(n_1248),
.C(n_1236),
.Y(n_2891)
);

AO22x2_ASAP7_75t_L g2892 ( 
.A1(n_2889),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_2892)
);

AOI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2884),
.A2(n_1316),
.B1(n_1011),
.B2(n_1019),
.Y(n_2893)
);

OAI222xp33_ASAP7_75t_L g2894 ( 
.A1(n_2875),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.C1(n_133),
.C2(n_134),
.Y(n_2894)
);

NAND4xp25_ASAP7_75t_L g2895 ( 
.A(n_2883),
.B(n_135),
.C(n_131),
.D(n_133),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2882),
.Y(n_2896)
);

NOR3xp33_ASAP7_75t_L g2897 ( 
.A(n_2881),
.B(n_839),
.C(n_1009),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2887),
.A2(n_1218),
.B1(n_1248),
.B2(n_1011),
.Y(n_2898)
);

OAI21xp33_ASAP7_75t_L g2899 ( 
.A1(n_2876),
.A2(n_839),
.B(n_135),
.Y(n_2899)
);

HB1xp67_ASAP7_75t_L g2900 ( 
.A(n_2878),
.Y(n_2900)
);

AOI22xp33_ASAP7_75t_L g2901 ( 
.A1(n_2885),
.A2(n_1038),
.B1(n_1043),
.B2(n_1041),
.Y(n_2901)
);

AOI221xp5_ASAP7_75t_L g2902 ( 
.A1(n_2877),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.C(n_145),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2879),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2874),
.Y(n_2904)
);

NOR3xp33_ASAP7_75t_L g2905 ( 
.A(n_2894),
.B(n_2886),
.C(n_2873),
.Y(n_2905)
);

NAND4xp75_ASAP7_75t_L g2906 ( 
.A(n_2904),
.B(n_976),
.C(n_141),
.D(n_145),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2900),
.B(n_139),
.Y(n_2907)
);

A2O1A1Ixp33_ASAP7_75t_SL g2908 ( 
.A1(n_2897),
.A2(n_147),
.B(n_148),
.C(n_149),
.Y(n_2908)
);

AOI21xp33_ASAP7_75t_SL g2909 ( 
.A1(n_2892),
.A2(n_147),
.B(n_149),
.Y(n_2909)
);

OAI22xp33_ASAP7_75t_SL g2910 ( 
.A1(n_2896),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_2910)
);

HB1xp67_ASAP7_75t_L g2911 ( 
.A(n_2892),
.Y(n_2911)
);

OAI321xp33_ASAP7_75t_L g2912 ( 
.A1(n_2893),
.A2(n_1218),
.A3(n_151),
.B1(n_152),
.B2(n_154),
.C(n_155),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2890),
.B(n_2903),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2899),
.B(n_150),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_2895),
.B(n_155),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2902),
.Y(n_2916)
);

AOI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2911),
.A2(n_2901),
.B1(n_2898),
.B2(n_2891),
.Y(n_2917)
);

AND2x4_ASAP7_75t_L g2918 ( 
.A(n_2913),
.B(n_156),
.Y(n_2918)
);

NOR2x1_ASAP7_75t_L g2919 ( 
.A(n_2907),
.B(n_2916),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2909),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2908),
.B(n_2915),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2910),
.B(n_157),
.Y(n_2922)
);

NOR3xp33_ASAP7_75t_L g2923 ( 
.A(n_2914),
.B(n_839),
.C(n_162),
.Y(n_2923)
);

NAND5xp2_ASAP7_75t_L g2924 ( 
.A(n_2905),
.B(n_162),
.C(n_163),
.D(n_166),
.E(n_167),
.Y(n_2924)
);

NOR3xp33_ASAP7_75t_SL g2925 ( 
.A(n_2906),
.B(n_163),
.C(n_166),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2912),
.Y(n_2926)
);

OAI22xp33_ASAP7_75t_SL g2927 ( 
.A1(n_2911),
.A2(n_168),
.B1(n_169),
.B2(n_172),
.Y(n_2927)
);

OR3x1_ASAP7_75t_L g2928 ( 
.A(n_2924),
.B(n_168),
.C(n_173),
.Y(n_2928)
);

AOI211xp5_ASAP7_75t_L g2929 ( 
.A1(n_2920),
.A2(n_173),
.B(n_174),
.C(n_175),
.Y(n_2929)
);

OAI211xp5_ASAP7_75t_L g2930 ( 
.A1(n_2921),
.A2(n_175),
.B(n_178),
.C(n_179),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2918),
.Y(n_2931)
);

AND4x1_ASAP7_75t_L g2932 ( 
.A(n_2919),
.B(n_178),
.C(n_179),
.D(n_180),
.Y(n_2932)
);

NOR2xp67_ASAP7_75t_L g2933 ( 
.A(n_2922),
.B(n_180),
.Y(n_2933)
);

NOR3xp33_ASAP7_75t_L g2934 ( 
.A(n_2927),
.B(n_182),
.C(n_183),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2925),
.Y(n_2935)
);

NAND3x1_ASAP7_75t_L g2936 ( 
.A(n_2923),
.B(n_183),
.C(n_184),
.Y(n_2936)
);

AOI211xp5_ASAP7_75t_L g2937 ( 
.A1(n_2926),
.A2(n_184),
.B(n_185),
.C(n_186),
.Y(n_2937)
);

AOI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_2917),
.A2(n_976),
.B1(n_1068),
.B2(n_1019),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2918),
.Y(n_2939)
);

NOR4xp25_ASAP7_75t_L g2940 ( 
.A(n_2920),
.B(n_186),
.C(n_187),
.D(n_188),
.Y(n_2940)
);

NAND3xp33_ASAP7_75t_L g2941 ( 
.A(n_2935),
.B(n_1017),
.C(n_1054),
.Y(n_2941)
);

XNOR2x1_ASAP7_75t_L g2942 ( 
.A(n_2931),
.B(n_188),
.Y(n_2942)
);

AND3x4_ASAP7_75t_L g2943 ( 
.A(n_2932),
.B(n_189),
.C(n_190),
.Y(n_2943)
);

NOR2x1p5_ASAP7_75t_L g2944 ( 
.A(n_2939),
.B(n_189),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2928),
.Y(n_2945)
);

AND3x4_ASAP7_75t_L g2946 ( 
.A(n_2934),
.B(n_190),
.C(n_191),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2933),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2940),
.B(n_191),
.Y(n_2948)
);

XNOR2x1_ASAP7_75t_L g2949 ( 
.A(n_2938),
.B(n_192),
.Y(n_2949)
);

AO22x2_ASAP7_75t_L g2950 ( 
.A1(n_2942),
.A2(n_2930),
.B1(n_2936),
.B2(n_2937),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2944),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_SL g2952 ( 
.A1(n_2945),
.A2(n_2929),
.B1(n_193),
.B2(n_194),
.Y(n_2952)
);

NOR4xp25_ASAP7_75t_L g2953 ( 
.A(n_2947),
.B(n_192),
.C(n_193),
.D(n_194),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2943),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_2954)
);

AO22x2_ASAP7_75t_L g2955 ( 
.A1(n_2946),
.A2(n_198),
.B1(n_200),
.B2(n_202),
.Y(n_2955)
);

AOI22xp5_ASAP7_75t_L g2956 ( 
.A1(n_2948),
.A2(n_1072),
.B1(n_1068),
.B2(n_1031),
.Y(n_2956)
);

AO22x2_ASAP7_75t_L g2957 ( 
.A1(n_2949),
.A2(n_200),
.B1(n_1017),
.B2(n_1048),
.Y(n_2957)
);

AOI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2941),
.A2(n_1068),
.B1(n_1072),
.B2(n_1031),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2943),
.A2(n_1068),
.B1(n_1072),
.B2(n_1031),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2944),
.Y(n_2960)
);

AOI22xp5_ASAP7_75t_L g2961 ( 
.A1(n_2943),
.A2(n_1072),
.B1(n_1031),
.B2(n_1029),
.Y(n_2961)
);

AOI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2943),
.A2(n_1029),
.B1(n_1022),
.B2(n_1027),
.Y(n_2962)
);

BUFx6f_ASAP7_75t_L g2963 ( 
.A(n_2945),
.Y(n_2963)
);

HB1xp67_ASAP7_75t_L g2964 ( 
.A(n_2944),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2943),
.A2(n_1029),
.B1(n_1022),
.B2(n_1027),
.Y(n_2965)
);

HB1xp67_ASAP7_75t_L g2966 ( 
.A(n_2944),
.Y(n_2966)
);

HB1xp67_ASAP7_75t_L g2967 ( 
.A(n_2944),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2944),
.Y(n_2968)
);

AOI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2943),
.A2(n_1029),
.B1(n_1022),
.B2(n_1027),
.Y(n_2969)
);

OAI31xp33_ASAP7_75t_L g2970 ( 
.A1(n_2954),
.A2(n_1027),
.A3(n_1022),
.B(n_1089),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2963),
.A2(n_1235),
.B1(n_1310),
.B2(n_1308),
.Y(n_2971)
);

AOI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2952),
.A2(n_1244),
.B1(n_1310),
.B2(n_1308),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2955),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2950),
.A2(n_1244),
.B1(n_1310),
.B2(n_1308),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2964),
.A2(n_1088),
.B1(n_1059),
.B2(n_1054),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2966),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2967),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2951),
.A2(n_1088),
.B1(n_1059),
.B2(n_1054),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2960),
.Y(n_2979)
);

CKINVDCx20_ASAP7_75t_R g2980 ( 
.A(n_2968),
.Y(n_2980)
);

AOI22xp5_ASAP7_75t_L g2981 ( 
.A1(n_2959),
.A2(n_1268),
.B1(n_1291),
.B2(n_1078),
.Y(n_2981)
);

AOI22xp33_ASAP7_75t_L g2982 ( 
.A1(n_2957),
.A2(n_1088),
.B1(n_1059),
.B2(n_1054),
.Y(n_2982)
);

AOI31xp33_ASAP7_75t_L g2983 ( 
.A1(n_2956),
.A2(n_1101),
.A3(n_1097),
.B(n_1096),
.Y(n_2983)
);

AOI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_2961),
.A2(n_1088),
.B1(n_1059),
.B2(n_1054),
.Y(n_2984)
);

OAI22xp5_ASAP7_75t_L g2985 ( 
.A1(n_2962),
.A2(n_1291),
.B1(n_1268),
.B2(n_1250),
.Y(n_2985)
);

NOR2x1_ASAP7_75t_L g2986 ( 
.A(n_2953),
.B(n_1048),
.Y(n_2986)
);

INVx5_ASAP7_75t_L g2987 ( 
.A(n_2965),
.Y(n_2987)
);

AOI31xp33_ASAP7_75t_L g2988 ( 
.A1(n_2969),
.A2(n_1101),
.A3(n_1097),
.B(n_1096),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2958),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2964),
.B(n_203),
.Y(n_2990)
);

AOI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2963),
.A2(n_1268),
.B1(n_1291),
.B2(n_1070),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2964),
.Y(n_2992)
);

BUFx2_ASAP7_75t_L g2993 ( 
.A(n_2955),
.Y(n_2993)
);

AOI22xp33_ASAP7_75t_L g2994 ( 
.A1(n_2963),
.A2(n_1088),
.B1(n_1059),
.B2(n_1054),
.Y(n_2994)
);

AOI31xp33_ASAP7_75t_L g2995 ( 
.A1(n_2964),
.A2(n_1092),
.A3(n_1091),
.B(n_1089),
.Y(n_2995)
);

XOR2xp5_ASAP7_75t_L g2996 ( 
.A(n_2980),
.B(n_208),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2976),
.B(n_219),
.Y(n_2997)
);

NAND4xp25_ASAP7_75t_L g2998 ( 
.A(n_2977),
.B(n_1092),
.C(n_1091),
.D(n_1086),
.Y(n_2998)
);

AOI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2992),
.A2(n_1078),
.B1(n_1060),
.B2(n_1070),
.Y(n_2999)
);

NOR2x1p5_ASAP7_75t_L g3000 ( 
.A(n_2973),
.B(n_832),
.Y(n_3000)
);

AOI222xp33_ASAP7_75t_L g3001 ( 
.A1(n_2993),
.A2(n_1060),
.B1(n_1077),
.B2(n_1083),
.C1(n_1084),
.C2(n_1086),
.Y(n_3001)
);

NAND5xp2_ASAP7_75t_L g3002 ( 
.A(n_2979),
.B(n_221),
.C(n_222),
.D(n_226),
.E(n_228),
.Y(n_3002)
);

OAI22xp5_ASAP7_75t_L g3003 ( 
.A1(n_2972),
.A2(n_1317),
.B1(n_1084),
.B2(n_1083),
.Y(n_3003)
);

OAI22x1_ASAP7_75t_L g3004 ( 
.A1(n_2987),
.A2(n_2990),
.B1(n_2986),
.B2(n_2989),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2987),
.B(n_235),
.Y(n_3005)
);

NOR2x1p5_ASAP7_75t_L g3006 ( 
.A(n_2987),
.B(n_832),
.Y(n_3006)
);

AOI221xp5_ASAP7_75t_L g3007 ( 
.A1(n_2995),
.A2(n_1059),
.B1(n_1088),
.B2(n_838),
.C(n_884),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2974),
.A2(n_1077),
.B1(n_1124),
.B2(n_1112),
.Y(n_3008)
);

OAI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2970),
.A2(n_1002),
.B(n_1003),
.Y(n_3009)
);

AOI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_2985),
.A2(n_1112),
.B1(n_1124),
.B2(n_1002),
.Y(n_3010)
);

AOI211xp5_ASAP7_75t_L g3011 ( 
.A1(n_2971),
.A2(n_2991),
.B(n_2981),
.C(n_2988),
.Y(n_3011)
);

OAI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2982),
.A2(n_1112),
.B1(n_1124),
.B2(n_838),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_SL g3013 ( 
.A1(n_2984),
.A2(n_1007),
.B1(n_1006),
.B2(n_1004),
.Y(n_3013)
);

AOI211xp5_ASAP7_75t_L g3014 ( 
.A1(n_2983),
.A2(n_884),
.B(n_838),
.C(n_846),
.Y(n_3014)
);

NOR4xp25_ASAP7_75t_L g3015 ( 
.A(n_2994),
.B(n_2975),
.C(n_2978),
.D(n_1124),
.Y(n_3015)
);

XOR2xp5_ASAP7_75t_L g3016 ( 
.A(n_2980),
.B(n_236),
.Y(n_3016)
);

NAND5xp2_ASAP7_75t_L g3017 ( 
.A(n_2976),
.B(n_237),
.C(n_248),
.D(n_250),
.E(n_253),
.Y(n_3017)
);

AOI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2980),
.A2(n_1112),
.B1(n_1004),
.B2(n_1003),
.Y(n_3018)
);

AOI221xp5_ASAP7_75t_L g3019 ( 
.A1(n_2993),
.A2(n_884),
.B1(n_838),
.B2(n_846),
.C(n_862),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2980),
.A2(n_1004),
.B1(n_1006),
.B2(n_1007),
.Y(n_3020)
);

AOI31xp33_ASAP7_75t_L g3021 ( 
.A1(n_3005),
.A2(n_2997),
.A3(n_3004),
.B(n_2996),
.Y(n_3021)
);

AOI31xp33_ASAP7_75t_L g3022 ( 
.A1(n_3016),
.A2(n_1007),
.A3(n_1006),
.B(n_259),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_3000),
.A2(n_880),
.B1(n_838),
.B2(n_846),
.Y(n_3023)
);

AOI31xp33_ASAP7_75t_L g3024 ( 
.A1(n_3011),
.A2(n_256),
.A3(n_258),
.B(n_261),
.Y(n_3024)
);

AOI31xp33_ASAP7_75t_L g3025 ( 
.A1(n_3014),
.A2(n_263),
.A3(n_264),
.B(n_266),
.Y(n_3025)
);

AOI31xp33_ASAP7_75t_L g3026 ( 
.A1(n_3019),
.A2(n_267),
.A3(n_269),
.B(n_271),
.Y(n_3026)
);

AOI31xp33_ASAP7_75t_L g3027 ( 
.A1(n_3020),
.A2(n_273),
.A3(n_275),
.B(n_276),
.Y(n_3027)
);

AOI31xp33_ASAP7_75t_L g3028 ( 
.A1(n_3001),
.A2(n_280),
.A3(n_282),
.B(n_284),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_3017),
.A2(n_880),
.B1(n_846),
.B2(n_862),
.Y(n_3029)
);

AOI31xp33_ASAP7_75t_L g3030 ( 
.A1(n_2999),
.A2(n_285),
.A3(n_292),
.B(n_298),
.Y(n_3030)
);

AOI22xp33_ASAP7_75t_L g3031 ( 
.A1(n_3002),
.A2(n_3006),
.B1(n_2998),
.B2(n_3013),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_3007),
.A2(n_880),
.B1(n_846),
.B2(n_862),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_3010),
.A2(n_884),
.B1(n_862),
.B2(n_863),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_3003),
.A2(n_884),
.B1(n_862),
.B2(n_863),
.Y(n_3034)
);

AOI22xp33_ASAP7_75t_L g3035 ( 
.A1(n_3012),
.A2(n_832),
.B1(n_863),
.B2(n_866),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_SL g3036 ( 
.A1(n_3031),
.A2(n_3015),
.B1(n_3018),
.B2(n_3008),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_3021),
.Y(n_3037)
);

AOI221xp5_ASAP7_75t_L g3038 ( 
.A1(n_3028),
.A2(n_3009),
.B1(n_880),
.B2(n_866),
.C(n_863),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_3033),
.A2(n_863),
.B1(n_866),
.B2(n_880),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_3034),
.A2(n_866),
.B1(n_1008),
.B2(n_1106),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_3022),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_3029),
.A2(n_866),
.B1(n_1008),
.B2(n_1106),
.Y(n_3042)
);

XOR2xp5_ASAP7_75t_L g3043 ( 
.A(n_3023),
.B(n_301),
.Y(n_3043)
);

OAI221xp5_ASAP7_75t_L g3044 ( 
.A1(n_3030),
.A2(n_1008),
.B1(n_304),
.B2(n_305),
.C(n_307),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_3025),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_3024),
.Y(n_3046)
);

OAI22xp5_ASAP7_75t_L g3047 ( 
.A1(n_3037),
.A2(n_3032),
.B1(n_3035),
.B2(n_3027),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_3041),
.Y(n_3048)
);

AOI21xp5_ASAP7_75t_L g3049 ( 
.A1(n_3045),
.A2(n_3026),
.B(n_1125),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_3046),
.B(n_302),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_3044),
.A2(n_1106),
.B1(n_1116),
.B2(n_1111),
.Y(n_3051)
);

OAI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_3043),
.A2(n_3038),
.B(n_3042),
.Y(n_3052)
);

AOI22xp5_ASAP7_75t_L g3053 ( 
.A1(n_3036),
.A2(n_1106),
.B1(n_311),
.B2(n_312),
.Y(n_3053)
);

AOI31xp33_ASAP7_75t_L g3054 ( 
.A1(n_3048),
.A2(n_3039),
.A3(n_3040),
.B(n_314),
.Y(n_3054)
);

OAI21x1_ASAP7_75t_L g3055 ( 
.A1(n_3047),
.A2(n_310),
.B(n_313),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_3049),
.A2(n_315),
.B(n_318),
.Y(n_3056)
);

AND2x2_ASAP7_75t_SL g3057 ( 
.A(n_3051),
.B(n_322),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_3057),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3054),
.Y(n_3059)
);

XNOR2xp5_ASAP7_75t_L g3060 ( 
.A(n_3056),
.B(n_3052),
.Y(n_3060)
);

OA21x2_ASAP7_75t_L g3061 ( 
.A1(n_3059),
.A2(n_3055),
.B(n_3050),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_3058),
.A2(n_3060),
.B(n_3053),
.Y(n_3062)
);

AOI221xp5_ASAP7_75t_L g3063 ( 
.A1(n_3062),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.C(n_327),
.Y(n_3063)
);

AOI211xp5_ASAP7_75t_L g3064 ( 
.A1(n_3063),
.A2(n_3061),
.B(n_331),
.C(n_333),
.Y(n_3064)
);


endmodule