module fake_jpeg_12118_n_393 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_56),
.B(n_57),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_64),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_67),
.B(n_69),
.Y(n_160)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_73),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_9),
.C(n_14),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_39),
.C(n_41),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_0),
.Y(n_72)
);

AND2x4_ASAP7_75t_SL g136 ( 
.A(n_72),
.B(n_61),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_74),
.B(n_81),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_77),
.B(n_84),
.Y(n_174)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_5),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_6),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_86),
.B(n_91),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_17),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_17),
.B(n_16),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_25),
.B(n_16),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_94),
.B(n_96),
.Y(n_154)
);

INVx2_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_38),
.B(n_16),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_97),
.B(n_100),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_11),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_104),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_20),
.B(n_11),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_39),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_22),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_113),
.Y(n_168)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_116),
.B(n_162),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_40),
.B1(n_37),
.B2(n_44),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_117),
.A2(n_150),
.B1(n_60),
.B2(n_104),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_136),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_37),
.B1(n_40),
.B2(n_44),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_132),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_33),
.B1(n_42),
.B2(n_30),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_139),
.B1(n_165),
.B2(n_105),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_47),
.B1(n_30),
.B2(n_41),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_65),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_152),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_78),
.B(n_52),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_103),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_59),
.A2(n_52),
.B1(n_46),
.B2(n_1),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_157),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_90),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_90),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_11),
.B1(n_79),
.B2(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_72),
.B(n_106),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_121),
.Y(n_213)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_60),
.B(n_102),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_194),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_99),
.C(n_102),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_182),
.B(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_123),
.A2(n_99),
.B(n_103),
.C(n_104),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_232),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_205),
.B(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_231),
.B1(n_114),
.B2(n_140),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g246 ( 
.A(n_197),
.B(n_202),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_200),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_203),
.B(n_214),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_75),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_75),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_206),
.B(n_207),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_82),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_82),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_145),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_129),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_210),
.B(n_215),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_123),
.B(n_137),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_213),
.B(n_222),
.Y(n_241)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_128),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_217),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_176),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_218),
.B(n_220),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_151),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_146),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_173),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_223),
.Y(n_266)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_165),
.A2(n_130),
.B1(n_117),
.B2(n_141),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_229),
.B1(n_192),
.B2(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_124),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_169),
.A2(n_150),
.B1(n_124),
.B2(n_167),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_125),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

OR2x4_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_125),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_234),
.A2(n_249),
.B(n_272),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_248),
.B1(n_274),
.B2(n_260),
.Y(n_295)
);

OAI22x1_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_114),
.B1(n_158),
.B2(n_169),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_245),
.A2(n_255),
.B1(n_258),
.B2(n_240),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_148),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_257),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_180),
.A2(n_148),
.B1(n_177),
.B2(n_227),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_177),
.B(n_191),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_177),
.B1(n_179),
.B2(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_204),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_211),
.A2(n_227),
.B1(n_229),
.B2(n_194),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_212),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_273),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_208),
.A2(n_192),
.B1(n_212),
.B2(n_183),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_260),
.A2(n_271),
.B1(n_274),
.B2(n_196),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_188),
.B(n_208),
.CI(n_232),
.CON(n_261),
.SN(n_261)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_187),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_193),
.A2(n_219),
.B1(n_226),
.B2(n_197),
.Y(n_271)
);

AOI32xp33_ASAP7_75t_L g272 ( 
.A1(n_202),
.A2(n_231),
.A3(n_218),
.B1(n_229),
.B2(n_181),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_201),
.B(n_190),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_224),
.B1(n_185),
.B2(n_181),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_275),
.A2(n_303),
.B(n_268),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_228),
.B(n_214),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_276),
.A2(n_294),
.B(n_256),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_184),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_281),
.B(n_282),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_254),
.B(n_184),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_199),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_284),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_186),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_293),
.B(n_300),
.Y(n_307)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_291),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_189),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_288),
.B(n_289),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_242),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_200),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_298),
.C(n_262),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_237),
.A2(n_250),
.B(n_243),
.Y(n_294)
);

NAND2x1_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_240),
.Y(n_306)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_301),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_261),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_299),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_247),
.C(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_239),
.B(n_258),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_250),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_242),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_305),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_244),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_270),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_322),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_241),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_323),
.C(n_290),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_315),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_302),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_240),
.B1(n_245),
.B2(n_264),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_317),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_264),
.B1(n_246),
.B2(n_236),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_234),
.B(n_266),
.Y(n_320)
);

AOI221xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_327),
.B1(n_276),
.B2(n_293),
.C(n_300),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_262),
.Y(n_323)
);

AO221x1_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_295),
.B1(n_305),
.B2(n_299),
.C(n_303),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_326),
.B(n_319),
.Y(n_353)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_325),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_298),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_335),
.C(n_337),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_286),
.B1(n_287),
.B2(n_285),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_316),
.B1(n_317),
.B2(n_311),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_294),
.C(n_292),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_301),
.C(n_277),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_340),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_277),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_342),
.C(n_343),
.Y(n_348)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_321),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_297),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_318),
.C(n_315),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_311),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_336),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_309),
.C(n_318),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_353),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_339),
.A2(n_327),
.B(n_336),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

OAI21x1_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_308),
.B(n_295),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_330),
.C(n_335),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_357),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_362),
.A2(n_337),
.B1(n_306),
.B2(n_295),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_351),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_366),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_367),
.B(n_368),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_296),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_348),
.A2(n_308),
.B(n_342),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_343),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_348),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_369),
.B(n_373),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_357),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_371),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_365),
.A2(n_350),
.B(n_355),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_334),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_347),
.C(n_306),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_370),
.B(n_373),
.Y(n_380)
);

AOI322xp5_ASAP7_75t_L g379 ( 
.A1(n_376),
.A2(n_365),
.A3(n_358),
.B1(n_360),
.B2(n_362),
.C1(n_347),
.C2(n_310),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_381),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_369),
.Y(n_385)
);

AOI322xp5_ASAP7_75t_L g381 ( 
.A1(n_375),
.A2(n_310),
.A3(n_314),
.B1(n_279),
.B2(n_278),
.C1(n_269),
.C2(n_268),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_378),
.B(n_374),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_377),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_384),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_380),
.B(n_386),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_388),
.A2(n_389),
.B(n_372),
.C(n_314),
.Y(n_391)
);

AOI211xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_390),
.B(n_279),
.C(n_256),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_279),
.Y(n_393)
);


endmodule