module real_jpeg_11664_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_6),
.A2(n_52),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_52),
.B1(n_59),
.B2(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_52),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_64),
.B1(n_72),
.B2(n_73),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_64),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_13),
.B(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_13),
.B(n_118),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_80),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_26),
.C(n_41),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_13),
.B(n_62),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_13),
.A2(n_104),
.B(n_145),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_58),
.B(n_61),
.C(n_172),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_13),
.A2(n_59),
.B1(n_61),
.B2(n_80),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_14),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_67),
.Y(n_179)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_19),
.B(n_107),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_85),
.B2(n_86),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_23)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_24),
.A2(n_29),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_24),
.B(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_25),
.B(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_29),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_38),
.B1(n_57),
.B2(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_37),
.B(n_135),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_38),
.A2(n_57),
.B(n_80),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_39),
.A2(n_46),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_49),
.B(n_50),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_43),
.A2(n_50),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_43),
.B(n_80),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_46),
.B(n_51),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.C(n_68),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_48),
.B(n_53),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_66),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_54),
.A2(n_90),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_59),
.B(n_77),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_73),
.A3(n_78),
.B1(n_82),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_65),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_69),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_79),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_80),
.B(n_81),
.C(n_83),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_80),
.B(n_106),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_98),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_97),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_106),
.A2(n_151),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_106),
.A2(n_120),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.C(n_113),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_111),
.B(n_113),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.C(n_119),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_198),
.B(n_202),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_183),
.B(n_197),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_167),
.B(n_182),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_147),
.B(n_166),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_136),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_131),
.A2(n_133),
.B(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_144),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_155),
.B(n_165),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_153),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_160),
.B(n_164),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_169),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_177),
.C(n_181),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_173),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_193),
.C(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);


endmodule