module real_aes_3576_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_673;
wire n_386;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_899;
wire n_637;
wire n_928;
wire n_155;
wire n_365;
wire n_243;
wire n_526;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_0), .Y(n_915) );
INVx1_ASAP7_75t_L g574 ( .A(n_1), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_2), .A2(n_15), .B1(n_134), .B2(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g618 ( .A(n_3), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_4), .A2(n_33), .B1(n_162), .B2(n_165), .Y(n_161) );
INVx1_ASAP7_75t_SL g672 ( .A(n_5), .Y(n_672) );
INVxp67_ASAP7_75t_L g110 ( .A(n_6), .Y(n_110) );
INVx1_ASAP7_75t_L g552 ( .A(n_6), .Y(n_552) );
INVx1_ASAP7_75t_L g903 ( .A(n_6), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_7), .A2(n_90), .B1(n_210), .B2(n_211), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_8), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_9), .B(n_156), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_10), .A2(n_34), .B1(n_131), .B2(n_133), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_11), .A2(n_531), .B1(n_532), .B2(n_533), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_11), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g537 ( .A1(n_11), .A2(n_532), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_SL g538 ( .A(n_11), .B(n_532), .Y(n_538) );
INVx2_ASAP7_75t_L g241 ( .A(n_12), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_13), .A2(n_56), .B1(n_147), .B2(n_580), .Y(n_579) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_14), .A2(n_69), .B(n_152), .Y(n_151) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_14), .A2(n_69), .B(n_152), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_16), .B(n_237), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_17), .A2(n_82), .B1(n_144), .B2(n_166), .Y(n_613) );
INVx2_ASAP7_75t_L g660 ( .A(n_18), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_19), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_SL g238 ( .A(n_20), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_21), .B(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_22), .A2(n_24), .B1(n_210), .B2(n_211), .Y(n_624) );
BUFx8_ASAP7_75t_SL g543 ( .A(n_23), .Y(n_543) );
BUFx3_ASAP7_75t_L g919 ( .A(n_23), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_25), .A2(n_64), .B1(n_163), .B2(n_616), .Y(n_615) );
O2A1O1Ixp5_ASAP7_75t_L g656 ( .A1(n_26), .A2(n_141), .B(n_162), .C(n_657), .Y(n_656) );
O2A1O1Ixp5_ASAP7_75t_L g259 ( .A1(n_27), .A2(n_140), .B(n_260), .C(n_263), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_28), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_29), .B(n_171), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_30), .A2(n_83), .B1(n_234), .B2(n_267), .Y(n_585) );
INVx1_ASAP7_75t_L g115 ( .A(n_31), .Y(n_115) );
INVx1_ASAP7_75t_L g653 ( .A(n_32), .Y(n_653) );
AND2x2_ASAP7_75t_L g924 ( .A(n_35), .B(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_36), .B(n_248), .Y(n_570) );
INVx2_ASAP7_75t_L g658 ( .A(n_37), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_38), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_39), .A2(n_44), .B1(n_170), .B2(n_172), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_40), .A2(n_68), .B1(n_172), .B2(n_193), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_41), .B(n_166), .Y(n_246) );
INVx2_ASAP7_75t_L g186 ( .A(n_42), .Y(n_186) );
INVx2_ASAP7_75t_L g632 ( .A(n_43), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_45), .A2(n_67), .B1(n_534), .B2(n_535), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_45), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_46), .B(n_171), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_47), .B(n_150), .Y(n_216) );
INVx1_ASAP7_75t_SL g675 ( .A(n_48), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_49), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_50), .A2(n_137), .B(n_234), .C(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g319 ( .A(n_51), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_52), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g597 ( .A(n_53), .Y(n_597) );
INVx2_ASAP7_75t_L g270 ( .A(n_54), .Y(n_270) );
INVx1_ASAP7_75t_L g152 ( .A(n_55), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_57), .B(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g201 ( .A(n_57), .B(n_154), .Y(n_201) );
INVx2_ASAP7_75t_L g195 ( .A(n_58), .Y(n_195) );
INVx1_ASAP7_75t_L g678 ( .A(n_59), .Y(n_678) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_60), .Y(n_138) );
INVx1_ASAP7_75t_SL g264 ( .A(n_61), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_62), .A2(n_104), .B1(n_920), .B2(n_928), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_63), .A2(n_79), .B1(n_908), .B2(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g909 ( .A(n_63), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_65), .B(n_637), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_66), .Y(n_199) );
CKINVDCx14_ASAP7_75t_R g535 ( .A(n_67), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_70), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_71), .A2(n_137), .B(n_162), .C(n_198), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_72), .Y(n_651) );
OR2x6_ASAP7_75t_L g112 ( .A(n_73), .B(n_113), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_74), .Y(n_305) );
INVx1_ASAP7_75t_L g315 ( .A(n_75), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_76), .B(n_167), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_77), .B(n_131), .Y(n_253) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_78), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g908 ( .A(n_79), .Y(n_908) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_80), .A2(n_190), .B(n_192), .C(n_196), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_80), .A2(n_190), .B(n_192), .C(n_196), .Y(n_295) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_84), .A2(n_96), .B1(n_143), .B2(n_147), .Y(n_142) );
INVx1_ASAP7_75t_L g925 ( .A(n_85), .Y(n_925) );
BUFx5_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_87), .B(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_88), .B(n_637), .Y(n_673) );
INVx2_ASAP7_75t_L g635 ( .A(n_89), .Y(n_635) );
INVx1_ASAP7_75t_L g640 ( .A(n_91), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_92), .A2(n_906), .B1(n_907), .B2(n_910), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_92), .Y(n_910) );
INVx2_ASAP7_75t_L g604 ( .A(n_93), .Y(n_604) );
INVx2_ASAP7_75t_SL g154 ( .A(n_94), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_95), .B(n_255), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_97), .B(n_157), .Y(n_316) );
INVx1_ASAP7_75t_SL g181 ( .A(n_98), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_99), .B(n_202), .Y(n_273) );
AND2x2_ASAP7_75t_L g155 ( .A(n_100), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_SL g268 ( .A(n_101), .Y(n_268) );
AO22x2_ASAP7_75t_L g620 ( .A1(n_102), .A2(n_321), .B1(n_621), .B2(n_625), .Y(n_620) );
AO32x2_ASAP7_75t_L g693 ( .A1(n_102), .A2(n_207), .A3(n_322), .B1(n_621), .B2(n_694), .Y(n_693) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_542), .B(n_544), .Y(n_104) );
OAI21x1_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_116), .B(n_539), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx10_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx8_ASAP7_75t_L g541 ( .A(n_108), .Y(n_541) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_108), .Y(n_927) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_L g902 ( .A(n_111), .B(n_903), .Y(n_902) );
INVx8_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g551 ( .A(n_112), .B(n_552), .Y(n_551) );
OR2x6_ASAP7_75t_L g917 ( .A(n_112), .B(n_552), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_530), .B1(n_536), .B2(n_537), .Y(n_118) );
INVx1_ASAP7_75t_L g536 ( .A(n_119), .Y(n_536) );
INVx2_ASAP7_75t_L g547 ( .A(n_119), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_119), .A2(n_554), .B1(n_899), .B2(n_912), .Y(n_911) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_442), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_362), .C(n_406), .Y(n_120) );
NOR3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_332), .C(n_350), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_285), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_217), .B1(n_274), .B2(n_282), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g418 ( .A(n_125), .Y(n_418) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_182), .Y(n_125) );
NOR2x1p5_ASAP7_75t_L g433 ( .A(n_126), .B(n_338), .Y(n_433) );
NAND2x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_158), .Y(n_126) );
INVx2_ASAP7_75t_L g277 ( .A(n_127), .Y(n_277) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g342 ( .A(n_128), .Y(n_342) );
AO31x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_139), .A3(n_148), .B(n_155), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_136), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_131), .A2(n_137), .B(n_675), .C(n_676), .Y(n_674) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g147 ( .A(n_132), .Y(n_147) );
INVx2_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVx1_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
INVx2_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
NAND2xp33_ASAP7_75t_L g227 ( .A(n_132), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g654 ( .A(n_133), .Y(n_654) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_134), .Y(n_234) );
INVx1_ASAP7_75t_L g269 ( .A(n_134), .Y(n_269) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
INVx2_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
INVx6_ASAP7_75t_L g237 ( .A(n_135), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_136), .A2(n_169), .B(n_173), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_136), .B(n_200), .Y(n_594) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_136), .B(n_200), .C(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_136), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_137), .A2(n_631), .B(n_632), .C(n_633), .Y(n_630) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_138), .Y(n_141) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_138), .Y(n_196) );
INVxp67_ASAP7_75t_L g213 ( .A(n_138), .Y(n_213) );
INVx4_ASAP7_75t_L g249 ( .A(n_138), .Y(n_249) );
INVx1_ASAP7_75t_L g587 ( .A(n_138), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_140), .B(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_140), .B(n_200), .Y(n_599) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_141), .A2(n_566), .B(n_568), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_141), .A2(n_231), .B1(n_622), .B2(n_624), .Y(n_621) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g164 ( .A(n_146), .Y(n_164) );
INVx2_ASAP7_75t_L g313 ( .A(n_147), .Y(n_313) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_149), .B(n_207), .Y(n_292) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_149), .A2(n_590), .B(n_603), .Y(n_589) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_150), .B(n_272), .Y(n_271) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
INVx2_ASAP7_75t_L g240 ( .A(n_151), .Y(n_240) );
INVx3_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_153), .Y(n_207) );
INVx1_ASAP7_75t_L g272 ( .A(n_153), .Y(n_272) );
INVx3_ASAP7_75t_L g576 ( .A(n_153), .Y(n_576) );
AND2x2_ASAP7_75t_L g611 ( .A(n_153), .B(n_223), .Y(n_611) );
AND2x2_ASAP7_75t_L g625 ( .A(n_153), .B(n_626), .Y(n_625) );
BUFx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_157), .B(n_576), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g582 ( .A(n_157), .B(n_576), .Y(n_582) );
INVx1_ASAP7_75t_L g605 ( .A(n_157), .Y(n_605) );
INVx1_ASAP7_75t_L g626 ( .A(n_157), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_157), .B(n_576), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_157), .Y(n_641) );
NOR2x1_ASAP7_75t_L g343 ( .A(n_158), .B(n_291), .Y(n_343) );
INVx1_ASAP7_75t_L g393 ( .A(n_158), .Y(n_393) );
AND2x2_ASAP7_75t_L g453 ( .A(n_158), .B(n_279), .Y(n_453) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g290 ( .A(n_159), .Y(n_290) );
AOI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_168), .B(n_179), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_162), .B(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g637 ( .A(n_164), .Y(n_637) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g211 ( .A(n_167), .Y(n_211) );
INVx1_ASAP7_75t_L g230 ( .A(n_167), .Y(n_230) );
INVx1_ASAP7_75t_L g567 ( .A(n_167), .Y(n_567) );
INVx1_ASAP7_75t_L g580 ( .A(n_167), .Y(n_580) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_172), .B(n_593), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_172), .A2(n_196), .B(n_635), .C(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_177), .Y(n_173) );
AOI21x1_ASAP7_75t_L g279 ( .A1(n_174), .A2(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g224 ( .A(n_176), .Y(n_224) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_177), .A2(n_245), .B(n_250), .Y(n_244) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_178), .A2(n_316), .B(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g202 ( .A(n_180), .Y(n_202) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g410 ( .A(n_183), .B(n_341), .Y(n_410) );
NOR2x1_ASAP7_75t_L g183 ( .A(n_184), .B(n_203), .Y(n_183) );
AND2x2_ASAP7_75t_L g366 ( .A(n_184), .B(n_342), .Y(n_366) );
INVx1_ASAP7_75t_L g432 ( .A(n_184), .Y(n_432) );
AND2x4_ASAP7_75t_L g440 ( .A(n_184), .B(n_277), .Y(n_440) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_184), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_184), .B(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_188), .Y(n_184) );
INVxp67_ASAP7_75t_SL g297 ( .A(n_185), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx1_ASAP7_75t_L g205 ( .A(n_187), .Y(n_205) );
NOR4xp25_ASAP7_75t_L g188 ( .A(n_189), .B(n_197), .C(n_200), .D(n_202), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g571 ( .A(n_191), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_193), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g267 ( .A(n_193), .Y(n_267) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g310 ( .A(n_194), .Y(n_310) );
INVx2_ASAP7_75t_SL g215 ( .A(n_196), .Y(n_215) );
INVx1_ASAP7_75t_L g231 ( .A(n_196), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_196), .B(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_196), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_196), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g614 ( .A(n_196), .Y(n_614) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_196), .A2(n_671), .B(n_672), .C(n_673), .Y(n_670) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_197), .Y(n_296) );
NOR2x1_ASAP7_75t_SL g221 ( .A(n_200), .B(n_222), .Y(n_221) );
AOI221x1_ASAP7_75t_L g647 ( .A1(n_200), .A2(n_648), .B1(n_650), .B2(n_652), .C(n_654), .Y(n_647) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_204), .Y(n_338) );
AND2x2_ASAP7_75t_L g361 ( .A(n_204), .B(n_289), .Y(n_361) );
INVx1_ASAP7_75t_L g489 ( .A(n_204), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_204), .B(n_342), .Y(n_492) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_216), .Y(n_204) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_205), .A2(n_244), .B(n_254), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_212), .B1(n_214), .B2(n_215), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_210), .A2(n_262), .B1(n_601), .B2(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g671 ( .A(n_211), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g265 ( .A1(n_212), .A2(n_266), .B(n_271), .Y(n_265) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g281 ( .A(n_216), .Y(n_281) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_242), .Y(n_217) );
OR2x6_ASAP7_75t_L g348 ( .A(n_218), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g460 ( .A(n_218), .B(n_370), .Y(n_460) );
INVx2_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g401 ( .A(n_219), .B(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_219), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g449 ( .A(n_219), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
OR2x2_ASAP7_75t_L g301 ( .A(n_220), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g356 ( .A(n_220), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g375 ( .A(n_220), .B(n_302), .Y(n_375) );
AND2x2_ASAP7_75t_L g425 ( .A(n_220), .B(n_357), .Y(n_425) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_220), .Y(n_503) );
AO31x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_225), .A3(n_232), .B(n_239), .Y(n_220) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_224), .B(n_576), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_229), .B(n_231), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_231), .A2(n_251), .B(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
INVx1_ASAP7_75t_L g649 ( .A(n_236), .Y(n_649) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g252 ( .A(n_237), .Y(n_252) );
INVx2_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
INVx1_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
INVx1_ASAP7_75t_L g616 ( .A(n_237), .Y(n_616) );
INVx2_ASAP7_75t_SL g623 ( .A(n_237), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx3_ASAP7_75t_L g255 ( .A(n_240), .Y(n_255) );
BUFx3_ASAP7_75t_L g322 ( .A(n_240), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_240), .B(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_240), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_256), .Y(n_242) );
AND2x2_ASAP7_75t_L g284 ( .A(n_243), .B(n_257), .Y(n_284) );
OR2x2_ASAP7_75t_L g408 ( .A(n_243), .B(n_356), .Y(n_408) );
AND2x2_ASAP7_75t_L g450 ( .A(n_243), .B(n_303), .Y(n_450) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_244), .A2(n_254), .B(n_321), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_248), .Y(n_245) );
AND2x2_ASAP7_75t_L g650 ( .A(n_248), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g652 ( .A(n_248), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
O2A1O1Ixp5_ASAP7_75t_SL g304 ( .A1(n_249), .A2(n_305), .B(n_306), .C(n_309), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_249), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g324 ( .A(n_256), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g500 ( .A(n_256), .B(n_283), .Y(n_500) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_257), .B(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g331 ( .A(n_258), .Y(n_331) );
INVx1_ASAP7_75t_L g389 ( .A(n_258), .Y(n_389) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_265), .B(n_273), .Y(n_258) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_262), .B(n_573), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B1(n_269), .B2(n_270), .Y(n_266) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g511 ( .A(n_275), .B(n_343), .Y(n_511) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
BUFx2_ASAP7_75t_SL g287 ( .A(n_277), .Y(n_287) );
INVx1_ASAP7_75t_L g354 ( .A(n_277), .Y(n_354) );
AND2x2_ASAP7_75t_L g394 ( .A(n_277), .B(n_291), .Y(n_394) );
AND2x2_ASAP7_75t_L g416 ( .A(n_278), .B(n_405), .Y(n_416) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g396 ( .A(n_279), .B(n_289), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_282), .B(n_435), .Y(n_434) );
INVxp33_ASAP7_75t_L g441 ( .A(n_282), .Y(n_441) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g379 ( .A(n_283), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_283), .Y(n_382) );
OR2x2_ASAP7_75t_L g461 ( .A(n_283), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g510 ( .A(n_283), .B(n_329), .Y(n_510) );
INVx1_ASAP7_75t_L g402 ( .A(n_284), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_298), .Y(n_285) );
INVx1_ASAP7_75t_L g371 ( .A(n_286), .Y(n_371) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_288), .B(n_338), .Y(n_385) );
INVx3_ASAP7_75t_L g487 ( .A(n_288), .Y(n_487) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g405 ( .A(n_290), .Y(n_405) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_291), .Y(n_528) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_297), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_323), .B(n_327), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g476 ( .A(n_301), .Y(n_476) );
OR2x2_ASAP7_75t_L g507 ( .A(n_301), .B(n_479), .Y(n_507) );
AND2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_302), .B(n_329), .Y(n_370) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g463 ( .A(n_303), .B(n_325), .Y(n_463) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_311), .B(n_320), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_304), .A2(n_311), .B(n_320), .Y(n_357) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_307), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g595 ( .A(n_310), .Y(n_595) );
NAND3x1_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .C(n_317), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AO31x2_ASAP7_75t_L g646 ( .A1(n_322), .A2(n_647), .A3(n_655), .B(n_659), .Y(n_646) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g400 ( .A(n_324), .B(n_375), .Y(n_400) );
INVxp67_ASAP7_75t_L g413 ( .A(n_324), .Y(n_413) );
INVx2_ASAP7_75t_L g329 ( .A(n_325), .Y(n_329) );
AND2x2_ASAP7_75t_L g383 ( .A(n_325), .B(n_331), .Y(n_383) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g419 ( .A(n_327), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx2_ASAP7_75t_L g429 ( .A(n_328), .Y(n_429) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_SL g349 ( .A(n_329), .Y(n_349) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_329), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_330), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g397 ( .A(n_330), .Y(n_397) );
INVx2_ASAP7_75t_SL g347 ( .A(n_331), .Y(n_347) );
BUFx2_ASAP7_75t_L g452 ( .A(n_331), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_344), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_337), .B(n_341), .Y(n_421) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g484 ( .A(n_338), .Y(n_484) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NOR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g355 ( .A(n_347), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g424 ( .A(n_347), .Y(n_424) );
AND2x2_ASAP7_75t_L g504 ( .A(n_347), .B(n_463), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_347), .B(n_425), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g527 ( .A(n_347), .B(n_353), .C(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g466 ( .A(n_348), .B(n_412), .Y(n_466) );
INVx1_ASAP7_75t_L g374 ( .A(n_349), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B(n_358), .C(n_360), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_353), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g395 ( .A(n_354), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g415 ( .A(n_354), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g438 ( .A(n_356), .B(n_424), .Y(n_438) );
INVx1_ASAP7_75t_L g516 ( .A(n_356), .Y(n_516) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_360), .A2(n_470), .B1(n_499), .B2(n_501), .C(n_505), .Y(n_498) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g365 ( .A(n_361), .B(n_366), .Y(n_365) );
NOR4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_376), .C(n_386), .D(n_398), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B1(n_371), .B2(n_372), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_364), .A2(n_377), .B1(n_380), .B2(n_384), .Y(n_376) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI21xp33_ASAP7_75t_SL g445 ( .A1(n_365), .A2(n_446), .B(n_447), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_366), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
AND2x2_ASAP7_75t_L g483 ( .A(n_366), .B(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g478 ( .A(n_369), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g480 ( .A1(n_372), .A2(n_481), .B(n_482), .C(n_485), .Y(n_480) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_375), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g456 ( .A(n_375), .B(n_429), .Y(n_456) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g496 ( .A(n_382), .B(n_450), .Y(n_496) );
INVx1_ASAP7_75t_L g521 ( .A(n_383), .Y(n_521) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g471 ( .A(n_385), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B1(n_395), .B2(n_397), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_388), .B(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_R g479 ( .A(n_389), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_390), .A2(n_438), .B1(n_439), .B2(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
NOR2xp33_ASAP7_75t_SL g529 ( .A(n_392), .B(n_488), .Y(n_529) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g523 ( .A(n_393), .B(n_410), .Y(n_523) );
AND2x4_ASAP7_75t_L g468 ( .A(n_394), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g513 ( .A(n_395), .Y(n_513) );
INVx2_ASAP7_75t_L g469 ( .A(n_396), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_401), .A2(n_466), .B1(n_467), .B2(n_470), .C(n_472), .Y(n_465) );
AND2x2_ASAP7_75t_L g477 ( .A(n_404), .B(n_432), .Y(n_477) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
INVx1_ASAP7_75t_L g495 ( .A(n_405), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_426), .C(n_437), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_411), .B2(n_414), .C(n_417), .Y(n_407) );
INVx1_ASAP7_75t_L g512 ( .A(n_408), .Y(n_512) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_412), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_416), .B(n_431), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_423), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_434), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g446 ( .A(n_438), .Y(n_446) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g457 ( .A(n_440), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g464 ( .A(n_440), .B(n_453), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_497), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_465), .C(n_480), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_455), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .C(n_454), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_449), .A2(n_457), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g524 ( .A(n_450), .B(n_479), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_459), .B2(n_464), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_468), .A2(n_516), .B1(n_517), .B2(n_520), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_474), .B1(n_477), .B2(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g481 ( .A(n_473), .Y(n_481) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_490), .B(n_496), .Y(n_485) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_492), .B(n_494), .Y(n_519) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_514), .Y(n_497) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .C(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_539), .A2(n_545), .B(n_918), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_904), .B1(n_905), .B2(n_911), .C(n_914), .Y(n_545) );
OAI22x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_553), .B2(n_898), .Y(n_546) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx8_ASAP7_75t_L g913 ( .A(n_551), .Y(n_913) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
NOR2x1p5_ASAP7_75t_L g555 ( .A(n_556), .B(n_790), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_758), .Y(n_556) );
NOR4xp25_ASAP7_75t_L g557 ( .A(n_558), .B(n_699), .C(n_725), .D(n_744), .Y(n_557) );
OAI211xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_606), .B(n_642), .C(n_687), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_560), .A2(n_681), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_588), .Y(n_560) );
AND2x2_ASAP7_75t_L g802 ( .A(n_561), .B(n_707), .Y(n_802) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_577), .Y(n_561) );
AND2x2_ASAP7_75t_L g666 ( .A(n_562), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g683 ( .A(n_562), .Y(n_683) );
INVx1_ASAP7_75t_L g734 ( .A(n_562), .Y(n_734) );
INVx2_ASAP7_75t_L g762 ( .A(n_562), .Y(n_762) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_562), .Y(n_893) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_569), .B(n_575), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B(n_572), .Y(n_569) );
INVx2_ASAP7_75t_L g664 ( .A(n_577), .Y(n_664) );
INVx1_ASAP7_75t_L g720 ( .A(n_577), .Y(n_720) );
AND2x2_ASAP7_75t_L g761 ( .A(n_577), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g843 ( .A(n_577), .Y(n_843) );
NAND2x1p5_ASAP7_75t_L g577 ( .A(n_578), .B(n_584), .Y(n_577) );
AND2x2_ASAP7_75t_SL g684 ( .A(n_578), .B(n_584), .Y(n_684) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B(n_583), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_582), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g763 ( .A(n_588), .Y(n_763) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g665 ( .A(n_589), .Y(n_665) );
OR2x2_ASAP7_75t_L g686 ( .A(n_589), .B(n_668), .Y(n_686) );
AND2x2_ASAP7_75t_L g889 ( .A(n_589), .B(n_729), .Y(n_889) );
AO21x2_ASAP7_75t_L g697 ( .A1(n_590), .A2(n_603), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_598), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g694 ( .A(n_605), .Y(n_694) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_619), .Y(n_607) );
INVx4_ASAP7_75t_L g661 ( .A(n_608), .Y(n_661) );
INVx2_ASAP7_75t_L g704 ( .A(n_608), .Y(n_704) );
AND2x2_ASAP7_75t_L g721 ( .A(n_608), .B(n_722), .Y(n_721) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g692 ( .A(n_609), .Y(n_692) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g680 ( .A(n_610), .Y(n_680) );
INVx1_ASAP7_75t_L g717 ( .A(n_610), .Y(n_717) );
AOI21x1_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B(n_617), .Y(n_610) );
INVx1_ASAP7_75t_L g631 ( .A(n_616), .Y(n_631) );
AND2x4_ASAP7_75t_L g768 ( .A(n_619), .B(n_740), .Y(n_768) );
AND2x4_ASAP7_75t_L g783 ( .A(n_619), .B(n_784), .Y(n_783) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_627), .Y(n_619) );
AND2x2_ASAP7_75t_L g679 ( .A(n_620), .B(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g710 ( .A(n_620), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g743 ( .A(n_620), .Y(n_743) );
INVx1_ASAP7_75t_L g840 ( .A(n_620), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_623), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g716 ( .A(n_627), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g722 ( .A(n_627), .B(n_646), .Y(n_722) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g645 ( .A(n_628), .B(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g702 ( .A(n_628), .B(n_703), .Y(n_702) );
BUFx3_ASAP7_75t_L g711 ( .A(n_628), .Y(n_711) );
INVx1_ASAP7_75t_L g742 ( .A(n_628), .Y(n_742) );
AND2x4_ASAP7_75t_L g816 ( .A(n_628), .B(n_817), .Y(n_816) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AO31x2_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .A3(n_638), .B(n_639), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NOR2xp33_ASAP7_75t_SL g677 ( .A(n_641), .B(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_662), .B1(n_679), .B2(n_681), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_645), .B(n_661), .Y(n_644) );
AND2x2_ASAP7_75t_L g754 ( .A(n_645), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g884 ( .A(n_645), .B(n_840), .Y(n_884) );
INVx2_ASAP7_75t_L g690 ( .A(n_646), .Y(n_690) );
OR2x2_ASAP7_75t_L g785 ( .A(n_646), .B(n_680), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_646), .B(n_680), .Y(n_788) );
INVx1_ASAP7_75t_L g817 ( .A(n_646), .Y(n_817) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
AND2x2_ASAP7_75t_L g696 ( .A(n_664), .B(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g708 ( .A(n_664), .Y(n_708) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_664), .Y(n_896) );
OR2x2_ASAP7_75t_L g733 ( .A(n_665), .B(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g751 ( .A(n_665), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g695 ( .A(n_666), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g738 ( .A(n_666), .B(n_720), .Y(n_738) );
INVx1_ASAP7_75t_L g752 ( .A(n_667), .Y(n_752) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g707 ( .A(n_668), .B(n_697), .Y(n_707) );
INVx2_ASAP7_75t_L g729 ( .A(n_668), .Y(n_729) );
INVx1_ASAP7_75t_L g747 ( .A(n_668), .Y(n_747) );
INVx1_ASAP7_75t_L g845 ( .A(n_668), .Y(n_845) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_668), .Y(n_849) );
AO31x2_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .A3(n_674), .B(n_677), .Y(n_668) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_680), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_681), .A2(n_768), .B1(n_770), .B2(n_771), .Y(n_769) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
AND2x2_ASAP7_75t_L g778 ( .A(n_682), .B(n_751), .Y(n_778) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_L g714 ( .A(n_683), .B(n_684), .Y(n_714) );
INVx1_ASAP7_75t_L g837 ( .A(n_683), .Y(n_837) );
AOI32xp33_ASAP7_75t_L g726 ( .A1(n_684), .A2(n_710), .A3(n_727), .B1(n_731), .B2(n_732), .Y(n_726) );
INVx2_ASAP7_75t_L g877 ( .A(n_684), .Y(n_877) );
INVx1_ASAP7_75t_L g724 ( .A(n_685), .Y(n_724) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_686), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_695), .Y(n_687) );
AND2x4_ASAP7_75t_SL g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx3_ASAP7_75t_L g740 ( .A(n_690), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_690), .B(n_703), .Y(n_776) );
AND2x2_ASAP7_75t_L g796 ( .A(n_690), .B(n_717), .Y(n_796) );
INVx2_ASAP7_75t_SL g808 ( .A(n_690), .Y(n_808) );
INVx1_ASAP7_75t_L g814 ( .A(n_691), .Y(n_814) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_692), .B(n_703), .Y(n_862) );
INVx2_ASAP7_75t_L g703 ( .A(n_693), .Y(n_703) );
BUFx8_ASAP7_75t_L g755 ( .A(n_693), .Y(n_755) );
INVxp67_ASAP7_75t_L g698 ( .A(n_694), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_695), .B(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_696), .B(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g773 ( .A(n_697), .B(n_762), .Y(n_773) );
AND2x2_ASAP7_75t_L g846 ( .A(n_697), .B(n_734), .Y(n_846) );
AND2x2_ASAP7_75t_L g876 ( .A(n_697), .B(n_877), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_705), .B1(n_709), .B2(n_713), .C(n_715), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx2_ASAP7_75t_L g806 ( .A(n_702), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_703), .B(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g804 ( .A(n_704), .B(n_710), .Y(n_804) );
NOR2x1_ASAP7_75t_L g805 ( .A(n_704), .B(n_806), .Y(n_805) );
OAI21xp33_ASAP7_75t_SL g766 ( .A1(n_705), .A2(n_767), .B(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g718 ( .A(n_707), .B(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g811 ( .A(n_708), .Y(n_811) );
AND2x2_ASAP7_75t_L g829 ( .A(n_708), .B(n_751), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx2_ASAP7_75t_SL g799 ( .A(n_711), .Y(n_799) );
OR2x2_ASAP7_75t_L g775 ( .A(n_712), .B(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_713), .B(n_763), .Y(n_789) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_714), .B(n_881), .Y(n_880) );
AOI22x1_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B1(n_721), .B2(n_723), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_716), .B(n_740), .Y(n_823) );
AND2x2_ASAP7_75t_L g831 ( .A(n_716), .B(n_740), .Y(n_831) );
INVx2_ASAP7_75t_L g730 ( .A(n_717), .Y(n_730) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_717), .Y(n_888) );
OAI21xp33_ASAP7_75t_L g735 ( .A1(n_718), .A2(n_736), .B(n_739), .Y(n_735) );
AND2x4_ASAP7_75t_L g771 ( .A(n_719), .B(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g848 ( .A(n_719), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g867 ( .A(n_719), .Y(n_867) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g731 ( .A(n_722), .B(n_730), .Y(n_731) );
AND2x2_ASAP7_75t_L g765 ( .A(n_722), .B(n_755), .Y(n_765) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_722), .Y(n_770) );
AND2x2_ASAP7_75t_L g872 ( .A(n_722), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_735), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_727), .B(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVxp67_ASAP7_75t_SL g854 ( .A(n_729), .Y(n_854) );
AND2x2_ASAP7_75t_L g757 ( .A(n_730), .B(n_741), .Y(n_757) );
INVx1_ASAP7_75t_L g781 ( .A(n_730), .Y(n_781) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g746 ( .A(n_734), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g750 ( .A(n_734), .Y(n_750) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
NAND4xp25_ASAP7_75t_L g841 ( .A(n_740), .B(n_755), .C(n_842), .D(n_846), .Y(n_841) );
AND2x2_ASAP7_75t_L g780 ( .A(n_741), .B(n_781), .Y(n_780) );
AND2x4_ASAP7_75t_SL g741 ( .A(n_742), .B(n_743), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_753), .C(n_756), .Y(n_744) );
OAI221xp5_ASAP7_75t_L g774 ( .A1(n_745), .A2(n_775), .B1(n_777), .B2(n_779), .C(n_782), .Y(n_774) );
AND2x4_ASAP7_75t_L g875 ( .A(n_746), .B(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
AND2x2_ASAP7_75t_L g809 ( .A(n_751), .B(n_761), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_751), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g786 ( .A(n_755), .B(n_787), .Y(n_786) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_755), .Y(n_857) );
AND2x2_ASAP7_75t_SL g871 ( .A(n_755), .B(n_816), .Y(n_871) );
INVx2_ASAP7_75t_L g873 ( .A(n_755), .Y(n_873) );
NOR3xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_766), .C(n_774), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_764), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
BUFx3_ASAP7_75t_L g850 ( .A(n_761), .Y(n_850) );
AND2x2_ASAP7_75t_L g882 ( .A(n_761), .B(n_763), .Y(n_882) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_L g824 ( .A(n_771), .Y(n_824) );
INVxp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OR2x6_ASAP7_75t_L g853 ( .A(n_773), .B(n_854), .Y(n_853) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_773), .Y(n_897) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_776), .Y(n_801) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_780), .A2(n_811), .B(n_812), .C(n_818), .Y(n_810) );
OAI21xp33_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_786), .B(n_789), .Y(n_782) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI21xp5_ASAP7_75t_SL g822 ( .A1(n_785), .A2(n_806), .B(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g827 ( .A(n_785), .Y(n_827) );
INVx2_ASAP7_75t_L g863 ( .A(n_786), .Y(n_863) );
AND2x4_ASAP7_75t_L g839 ( .A(n_787), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_858), .Y(n_790) );
NOR3xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_820), .C(n_832), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_803), .C(n_810), .Y(n_792) );
OAI21xp33_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_797), .B(n_802), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_796), .B(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_800), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g826 ( .A(n_799), .B(n_827), .Y(n_826) );
OAI32xp33_ASAP7_75t_L g885 ( .A1(n_799), .A2(n_883), .A3(n_886), .B1(n_890), .B2(n_894), .Y(n_885) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OAI31xp33_ASAP7_75t_SL g803 ( .A1(n_804), .A2(n_805), .A3(n_807), .B(n_809), .Y(n_803) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVxp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_824), .B1(n_825), .B2(n_828), .C(n_830), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_847), .C(n_851), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_838), .B(n_841), .Y(n_834) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
OAI21xp33_ASAP7_75t_L g847 ( .A1(n_839), .A2(n_848), .B(n_850), .Y(n_847) );
AND2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_844), .Y(n_881) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_855), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g868 ( .A(n_853), .Y(n_868) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_869), .C(n_885), .Y(n_858) );
AOI21x1_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_863), .B(n_864), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AND2x4_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .Y(n_865) );
INVxp67_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_874), .B1(n_878), .B2(n_883), .Y(n_869) );
NOR2xp33_ASAP7_75t_SL g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NOR2xp33_ASAP7_75t_SL g878 ( .A(n_879), .B(n_882), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
AND2x4_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
BUFx3_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
BUFx12f_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
CKINVDCx11_ASAP7_75t_R g900 ( .A(n_901), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_SL g912 ( .A(n_913), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
BUFx3_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
CKINVDCx6p67_ASAP7_75t_R g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_SL g921 ( .A(n_922), .Y(n_921) );
BUFx2_ASAP7_75t_SL g929 ( .A(n_922), .Y(n_929) );
BUFx5_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
AND2x6_ASAP7_75t_L g923 ( .A(n_924), .B(n_926), .Y(n_923) );
INVx5_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
endmodule