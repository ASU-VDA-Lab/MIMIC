module fake_jpeg_14491_n_601 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_601);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_59),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_6),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_64),
.Y(n_126)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_23),
.B(n_6),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_79),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_78),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_23),
.B(n_6),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_80),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_81),
.B(n_86),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_32),
.B(n_6),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g149 ( 
.A(n_87),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_93),
.B(n_101),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_32),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_38),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_102),
.B(n_103),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_39),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_39),
.B(n_14),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_24),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_44),
.Y(n_113)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_42),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_123),
.B(n_183),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_62),
.B(n_50),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_138),
.B(n_139),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_66),
.B(n_50),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_78),
.A2(n_28),
.B1(n_49),
.B2(n_16),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_181),
.B1(n_89),
.B2(n_24),
.Y(n_201)
);

AO22x2_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_43),
.B1(n_42),
.B2(n_35),
.Y(n_153)
);

AOI22x1_ASAP7_75t_L g214 ( 
.A1(n_153),
.A2(n_56),
.B1(n_114),
.B2(n_116),
.Y(n_214)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_176),
.Y(n_220)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_87),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_57),
.Y(n_180)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_71),
.A2(n_43),
.B1(n_48),
.B2(n_27),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_60),
.B(n_52),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_192),
.Y(n_234)
);

BUFx4f_ASAP7_75t_SL g189 ( 
.A(n_68),
.Y(n_189)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_90),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_72),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_201),
.A2(n_211),
.B1(n_214),
.B2(n_216),
.Y(n_307)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_204),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_128),
.B(n_56),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_166),
.C(n_165),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_141),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_222),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_52),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_210),
.B(n_231),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_153),
.A2(n_98),
.B1(n_94),
.B2(n_112),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_212),
.Y(n_290)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_213),
.Y(n_328)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_153),
.A2(n_96),
.B1(n_84),
.B2(n_99),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_218),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_159),
.A2(n_28),
.B1(n_65),
.B2(n_21),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_223),
.A2(n_254),
.B1(n_259),
.B2(n_168),
.Y(n_300)
);

CKINVDCx9p33_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_224),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_125),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_232),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_133),
.B(n_36),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_227),
.B(n_229),
.Y(n_316)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_122),
.B(n_36),
.Y(n_229)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_129),
.Y(n_230)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_230),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_35),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_170),
.A2(n_48),
.B(n_30),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_146),
.A2(n_97),
.B1(n_100),
.B2(n_80),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_257),
.B1(n_4),
.B2(n_11),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_170),
.B(n_29),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_245),
.Y(n_284)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_125),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_240),
.Y(n_279)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_130),
.A2(n_91),
.B1(n_83),
.B2(n_27),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_239),
.A2(n_160),
.B1(n_148),
.B2(n_132),
.Y(n_280)
);

OR2x4_ASAP7_75t_L g240 ( 
.A(n_126),
.B(n_40),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_150),
.Y(n_241)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_127),
.A2(n_43),
.B1(n_88),
.B2(n_82),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_242),
.A2(n_143),
.B1(n_135),
.B2(n_137),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_127),
.B(n_29),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_155),
.B(n_109),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_246),
.B(n_250),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_142),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_255),
.Y(n_296)
);

CKINVDCx12_ASAP7_75t_R g249 ( 
.A(n_154),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_249),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_126),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx11_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_134),
.B(n_25),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_265),
.Y(n_285)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_164),
.A2(n_25),
.B1(n_66),
.B2(n_70),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_172),
.A2(n_30),
.B1(n_21),
.B2(n_82),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_256),
.A2(n_196),
.B1(n_186),
.B2(n_137),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_136),
.A2(n_109),
.B1(n_88),
.B2(n_9),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_131),
.A2(n_5),
.B1(n_10),
.B2(n_9),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_162),
.Y(n_260)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_157),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_269),
.Y(n_310)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_167),
.Y(n_263)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_173),
.A2(n_158),
.B(n_182),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_0),
.B(n_2),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_185),
.B(n_0),
.Y(n_265)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_167),
.Y(n_266)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_162),
.Y(n_267)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_124),
.Y(n_269)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

CKINVDCx12_ASAP7_75t_R g271 ( 
.A(n_191),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_271),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_278),
.A2(n_280),
.B1(n_287),
.B2(n_308),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_205),
.B(n_145),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_286),
.A2(n_292),
.B(n_299),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_214),
.A2(n_129),
.B1(n_135),
.B2(n_190),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_304),
.C(n_255),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_214),
.A2(n_151),
.B1(n_144),
.B2(n_166),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_165),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_327),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_205),
.B(n_124),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_254),
.B1(n_233),
.B2(n_212),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_194),
.C(n_5),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_265),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_254),
.A2(n_212),
.B1(n_258),
.B2(n_206),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_320),
.A2(n_256),
.B1(n_264),
.B2(n_236),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_252),
.A2(n_4),
.B1(n_9),
.B2(n_11),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_322),
.A2(n_324),
.B1(n_269),
.B2(n_217),
.Y(n_345)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_206),
.Y(n_325)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_229),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_218),
.B1(n_227),
.B2(n_224),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_231),
.B(n_210),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_329),
.A2(n_290),
.B1(n_328),
.B2(n_294),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_226),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_330),
.B(n_335),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_240),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_331),
.B(n_355),
.Y(n_387)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_332),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_235),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_245),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_337),
.B(n_341),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_285),
.B(n_225),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_234),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_348),
.Y(n_381)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_272),
.B(n_209),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_346),
.B(n_349),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_307),
.A2(n_254),
.B1(n_228),
.B2(n_204),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_361),
.B1(n_302),
.B2(n_293),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_282),
.B(n_327),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_310),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_282),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_350),
.B(n_359),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_284),
.B(n_219),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_356),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_318),
.Y(n_390)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_354),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_284),
.B(n_247),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_243),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_304),
.B(n_220),
.CI(n_247),
.CON(n_358),
.SN(n_358)
);

FAx1_ASAP7_75t_SL g393 ( 
.A(n_358),
.B(n_283),
.CI(n_325),
.CON(n_393),
.SN(n_393)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_203),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_244),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_360),
.B(n_363),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_307),
.A2(n_244),
.B1(n_221),
.B2(n_270),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_287),
.B(n_281),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_365),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_221),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_293),
.B(n_203),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_290),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_281),
.B(n_268),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_298),
.B(n_267),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_312),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_313),
.A2(n_215),
.B1(n_213),
.B2(n_260),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_367),
.A2(n_302),
.B1(n_283),
.B2(n_297),
.Y(n_382)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

INVx13_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_311),
.B(n_297),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_384),
.B(n_396),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_371),
.A2(n_278),
.B1(n_309),
.B2(n_317),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_375),
.A2(n_376),
.B1(n_382),
.B2(n_403),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_306),
.B1(n_309),
.B2(n_317),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_363),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_368),
.A2(n_298),
.B(n_312),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_385),
.A2(n_399),
.B1(n_405),
.B2(n_340),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_364),
.Y(n_423)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_400),
.Y(n_415)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_395),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_339),
.B(n_350),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_306),
.B1(n_328),
.B2(n_294),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_314),
.C(n_305),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_334),
.B(n_314),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_407),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_334),
.A2(n_202),
.B1(n_266),
.B2(n_238),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_342),
.A2(n_315),
.B1(n_301),
.B2(n_323),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_348),
.B(n_305),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_400),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_409),
.B(n_420),
.C(n_401),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_396),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_410),
.B(n_416),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_388),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_411),
.A2(n_419),
.B(n_430),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_414),
.B(n_403),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_346),
.Y(n_416)
);

INVx13_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_418),
.Y(n_467)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_329),
.B(n_362),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_343),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_356),
.Y(n_421)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_377),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_431),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_423),
.A2(n_433),
.B1(n_375),
.B2(n_399),
.Y(n_471)
);

AOI22x1_ASAP7_75t_L g424 ( 
.A1(n_394),
.A2(n_355),
.B1(n_366),
.B2(n_332),
.Y(n_424)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

INVx13_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_425),
.Y(n_462)
);

INVx8_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_428),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_392),
.B(n_330),
.Y(n_428)
);

NAND2x1_ASAP7_75t_SL g429 ( 
.A(n_372),
.B(n_332),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_429),
.A2(n_379),
.B(n_383),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_408),
.A2(n_353),
.B(n_365),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_381),
.B(n_341),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_340),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_432),
.A2(n_383),
.B(n_344),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_404),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_436),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_377),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_397),
.B(n_335),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_437),
.B(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_402),
.B(n_337),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_441),
.C(n_331),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_351),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_376),
.A2(n_360),
.B1(n_358),
.B2(n_369),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_442),
.A2(n_358),
.B1(n_391),
.B2(n_389),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_452),
.C(n_454),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_444),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_397),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_453),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_432),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_446),
.B(n_470),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_429),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_448),
.B(n_460),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_386),
.B1(n_408),
.B2(n_406),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_449),
.A2(n_457),
.B1(n_472),
.B2(n_419),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_429),
.A2(n_393),
.B(n_406),
.Y(n_451)
);

AOI21xp33_ASAP7_75t_L g489 ( 
.A1(n_451),
.A2(n_424),
.B(n_411),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_380),
.C(n_393),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_359),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_378),
.C(n_374),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_378),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_427),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_414),
.C(n_410),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_438),
.C(n_434),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_423),
.Y(n_460)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_432),
.A2(n_442),
.B(n_424),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_465),
.B(n_423),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_412),
.A2(n_405),
.B(n_373),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_430),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_419),
.B1(n_421),
.B2(n_434),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_440),
.A2(n_398),
.B1(n_336),
.B2(n_274),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_466),
.A2(n_413),
.B1(n_436),
.B2(n_422),
.Y(n_474)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_474),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_476),
.B(n_452),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_445),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_477),
.B(n_485),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_480),
.A2(n_499),
.B1(n_471),
.B2(n_460),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_456),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_482),
.B(n_493),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_439),
.C(n_431),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_463),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_412),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_444),
.B(n_467),
.Y(n_523)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_489),
.A2(n_468),
.B(n_451),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_490),
.B(n_491),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_427),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_500),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_426),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_455),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_495),
.B(n_501),
.Y(n_514)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_469),
.Y(n_496)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_496),
.Y(n_522)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_497),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_449),
.A2(n_433),
.B1(n_398),
.B2(n_336),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_454),
.B(n_354),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_457),
.B(n_354),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_447),
.Y(n_502)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_484),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_447),
.Y(n_504)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_494),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_511),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_510),
.B(n_520),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_458),
.C(n_450),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_516),
.A2(n_472),
.B1(n_462),
.B2(n_490),
.Y(n_535)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_517),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_478),
.A2(n_464),
.B1(n_473),
.B2(n_467),
.Y(n_519)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_519),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_450),
.C(n_465),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_521),
.Y(n_539)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_523),
.A2(n_464),
.B(n_476),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_481),
.B(n_473),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_524),
.B(n_475),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_480),
.B(n_494),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_529),
.Y(n_550)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_523),
.A2(n_448),
.B(n_481),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_527),
.A2(n_534),
.B(n_507),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_491),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_528),
.B(n_538),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_530),
.B(n_487),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_487),
.C(n_484),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_537),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_505),
.A2(n_485),
.B(n_499),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_516),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_509),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_513),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_515),
.B(n_500),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_540),
.B(n_508),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_542),
.B(n_512),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_544),
.B(n_545),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_518),
.C(n_508),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_546),
.B(n_549),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_547),
.A2(n_555),
.B(n_537),
.Y(n_568)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_511),
.Y(n_548)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_548),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_543),
.A2(n_520),
.B(n_509),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_526),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_558),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_527),
.A2(n_507),
.B(n_522),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_536),
.Y(n_557)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_557),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_518),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_503),
.C(n_502),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_559),
.B(n_512),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_541),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_562),
.B(n_567),
.Y(n_577)
);

AO21x1_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_532),
.B(n_537),
.Y(n_563)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_563),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_572),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_517),
.Y(n_567)
);

AO21x1_ASAP7_75t_L g574 ( 
.A1(n_568),
.A2(n_555),
.B(n_558),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_552),
.A2(n_525),
.B1(n_531),
.B2(n_556),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_569),
.B(n_571),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_550),
.A2(n_525),
.B1(n_529),
.B2(n_425),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_570),
.A2(n_547),
.B(n_546),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_573),
.B(n_576),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_574),
.A2(n_561),
.B1(n_565),
.B2(n_276),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_560),
.B(n_559),
.C(n_553),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_563),
.A2(n_418),
.B(n_301),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_578),
.A2(n_370),
.B(n_276),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_315),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_580),
.B(n_581),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_323),
.C(n_289),
.Y(n_581)
);

AO21x1_ASAP7_75t_L g584 ( 
.A1(n_575),
.A2(n_568),
.B(n_572),
.Y(n_584)
);

OAI211xp5_ASAP7_75t_L g590 ( 
.A1(n_584),
.A2(n_574),
.B(n_582),
.C(n_581),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_565),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_585),
.B(n_587),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_579),
.B(n_370),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_SL g592 ( 
.A(n_588),
.B(n_582),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_589),
.B(n_587),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_590),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_592),
.A2(n_593),
.B(n_586),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_591),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_596),
.B(n_597),
.C(n_289),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_594),
.B(n_583),
.Y(n_597)
);

OAI21xp33_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_273),
.B(n_230),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_207),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_241),
.B1(n_263),
.B2(n_273),
.Y(n_601)
);


endmodule