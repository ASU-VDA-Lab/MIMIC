module fake_netlist_1_2487_n_813 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_813);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_813;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_177;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g165 ( .A(n_17), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_17), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_47), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_152), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_93), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_114), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_10), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_124), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g175 ( .A(n_79), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_158), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_87), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_32), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_104), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_55), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_6), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_64), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_119), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_70), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_65), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_140), .Y(n_189) );
INVxp33_ASAP7_75t_SL g190 ( .A(n_41), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_105), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_19), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_96), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_53), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_128), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_85), .B(n_40), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_74), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_71), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_139), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_41), .Y(n_206) );
INVxp33_ASAP7_75t_SL g207 ( .A(n_20), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_12), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_130), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_160), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_16), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_103), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_49), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_31), .Y(n_218) );
NOR2xp67_ASAP7_75t_L g219 ( .A(n_102), .B(n_127), .Y(n_219) );
INVxp33_ASAP7_75t_SL g220 ( .A(n_26), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_16), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_36), .Y(n_222) );
CKINVDCx14_ASAP7_75t_R g223 ( .A(n_115), .Y(n_223) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_151), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_20), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_11), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_27), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_60), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_49), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_71), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_18), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_44), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_11), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_90), .Y(n_235) );
BUFx2_ASAP7_75t_SL g236 ( .A(n_9), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_56), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_66), .Y(n_238) );
INVxp33_ASAP7_75t_L g239 ( .A(n_154), .Y(n_239) );
CKINVDCx14_ASAP7_75t_R g240 ( .A(n_112), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_116), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_29), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_25), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_129), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_113), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_134), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_100), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_107), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_156), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_121), .Y(n_250) );
INVxp67_ASAP7_75t_SL g251 ( .A(n_125), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_25), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_89), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_30), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_8), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_92), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_88), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_21), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_81), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_29), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_44), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_91), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_37), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_170), .Y(n_264) );
AND2x6_ASAP7_75t_L g265 ( .A(n_170), .B(n_72), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_191), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_172), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_191), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_172), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_173), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_191), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_228), .B(n_0), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_173), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_191), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_174), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_174), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_171), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_171), .Y(n_278) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_176), .A2(n_75), .B(n_73), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_196), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_176), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_195), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_195), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_196), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_177), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_239), .B(n_1), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_228), .B(n_169), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_222), .B(n_1), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_179), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_179), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_180), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_193), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_195), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_195), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_184), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_218), .B(n_2), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_187), .A2(n_77), .B(n_76), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_295), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_274), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_288), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_264), .A2(n_183), .B1(n_188), .B2(n_182), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_277), .B(n_257), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_292), .B(n_201), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_274), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_264), .A2(n_183), .B1(n_188), .B2(n_182), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_277), .B(n_222), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_278), .B(n_230), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
AO22x2_ASAP7_75t_L g313 ( .A1(n_297), .A2(n_199), .B1(n_192), .B2(n_197), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_265), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
AND2x6_ASAP7_75t_L g318 ( .A(n_288), .B(n_187), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_278), .B(n_184), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_267), .B(n_269), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_274), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_280), .B(n_230), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_280), .B(n_175), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_265), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_280), .B(n_223), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_267), .B(n_186), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_269), .B(n_186), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_288), .B(n_284), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_265), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_284), .B(n_240), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
INVx4_ASAP7_75t_L g337 ( .A(n_265), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_270), .B(n_212), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_271), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_273), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_273), .B(n_212), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_305), .B(n_287), .Y(n_343) );
BUFx4f_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_313), .B(n_297), .Y(n_345) );
BUFx8_ASAP7_75t_L g346 ( .A(n_307), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_305), .B(n_275), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_302), .A2(n_275), .B(n_281), .C(n_276), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
XNOR2xp5_ASAP7_75t_SL g354 ( .A(n_304), .B(n_178), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_302), .Y(n_355) );
OR2x6_ASAP7_75t_L g356 ( .A(n_313), .B(n_236), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
INVx4_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_300), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_329), .B(n_286), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_313), .A2(n_265), .B1(n_281), .B2(n_276), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_329), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_304), .B(n_285), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_318), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_318), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_316), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_335), .B(n_285), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_325), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_313), .A2(n_207), .B1(n_220), .B2(n_190), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_333), .B(n_272), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_335), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_325), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
INVx4_ASAP7_75t_L g381 ( .A(n_318), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_334), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_333), .B(n_289), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_302), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_318), .A2(n_265), .B1(n_290), .B2(n_289), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_319), .B(n_291), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_302), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_318), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_309), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_320), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_315), .B(n_337), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_320), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_320), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_309), .B(n_291), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_309), .B(n_296), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_309), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_319), .B(n_296), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_311), .B(n_194), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_311), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_311), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_311), .B(n_168), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_393), .A2(n_337), .B(n_315), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_348), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_350), .A2(n_321), .B(n_340), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_346), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_343), .B(n_340), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_376), .B(n_324), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_345), .A2(n_227), .B1(n_238), .B2(n_181), .Y(n_410) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_370), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_352), .B(n_353), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_373), .B(n_324), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_376), .B(n_324), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_373), .B(n_324), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_350), .A2(n_338), .B(n_331), .Y(n_417) );
INVx6_ASAP7_75t_SL g418 ( .A(n_345), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_401), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
INVx5_ASAP7_75t_L g421 ( .A(n_359), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_384), .Y(n_423) );
NOR2x1_ASAP7_75t_SL g424 ( .A(n_356), .B(n_315), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_349), .B(n_321), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_371), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_365), .B(n_308), .C(n_303), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_355), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_357), .B(n_227), .Y(n_429) );
BUFx6f_ASAP7_75t_SL g430 ( .A(n_400), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_360), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_L g432 ( .A1(n_388), .A2(n_341), .B(n_332), .C(n_308), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_360), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_355), .Y(n_434) );
BUFx5_ASAP7_75t_L g435 ( .A(n_371), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_391), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_344), .Y(n_437) );
INVx8_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_375), .B(n_185), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_372), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_344), .Y(n_441) );
BUFx4_ASAP7_75t_SL g442 ( .A(n_377), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_403), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g444 ( .A(n_359), .B(n_265), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_372), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_344), .Y(n_446) );
INVx4_ASAP7_75t_L g447 ( .A(n_359), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_399), .A2(n_167), .B1(n_208), .B2(n_166), .C(n_165), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_392), .A2(n_298), .B(n_279), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_374), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_367), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_385), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_378), .Y(n_454) );
INVx3_ASAP7_75t_SL g455 ( .A(n_377), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_369), .B(n_265), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_354), .Y(n_457) );
OR2x6_ASAP7_75t_L g458 ( .A(n_379), .B(n_255), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_342), .A2(n_203), .B1(n_217), .B2(n_215), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_358), .A2(n_198), .B(n_200), .C(n_192), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_392), .A2(n_298), .B(n_279), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_379), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_351), .A2(n_221), .B1(n_226), .B2(n_217), .Y(n_463) );
BUFx12f_ASAP7_75t_L g464 ( .A(n_362), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_397), .Y(n_465) );
BUFx12f_ASAP7_75t_L g466 ( .A(n_362), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_397), .B(n_229), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_363), .B(n_237), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_381), .B(n_258), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_381), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_389), .B(n_231), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_390), .A2(n_261), .B1(n_260), .B2(n_232), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_380), .Y(n_473) );
AOI33xp33_ASAP7_75t_L g474 ( .A1(n_386), .A2(n_233), .A3(n_263), .B1(n_234), .B2(n_254), .B3(n_252), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_368), .B(n_242), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_410), .A2(n_395), .B1(n_394), .B2(n_382), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_433), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_405), .B(n_206), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_395), .B1(n_382), .B2(n_387), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_427), .A2(n_387), .B1(n_380), .B2(n_243), .Y(n_480) );
OAI21x1_ASAP7_75t_L g481 ( .A1(n_449), .A2(n_298), .B(n_279), .Y(n_481) );
AOI21x1_ASAP7_75t_L g482 ( .A1(n_449), .A2(n_298), .B(n_279), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_450), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_408), .A2(n_361), .B(n_347), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_405), .B(n_368), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_473), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_414), .A2(n_202), .B1(n_204), .B2(n_200), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_421), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_416), .A2(n_204), .B1(n_205), .B2(n_202), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_467), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_467), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_407), .B(n_347), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g493 ( .A1(n_457), .A2(n_256), .B1(n_262), .B2(n_250), .C1(n_224), .C2(n_251), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_429), .B(n_455), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_458), .B(n_347), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_408), .A2(n_209), .B1(n_211), .B2(n_210), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_471), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_448), .A2(n_219), .B(n_214), .C(n_216), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
INVx4_ASAP7_75t_SL g500 ( .A(n_430), .Y(n_500) );
OR2x6_ASAP7_75t_L g501 ( .A(n_438), .B(n_347), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_430), .A2(n_298), .B1(n_279), .B2(n_213), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_412), .B(n_3), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_468), .Y(n_504) );
AO21x1_ASAP7_75t_L g505 ( .A1(n_444), .A2(n_294), .B(n_271), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_442), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_468), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_418), .Y(n_508) );
OAI21x1_ASAP7_75t_SL g509 ( .A1(n_424), .A2(n_235), .B(n_225), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_404), .A2(n_366), .B(n_364), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_464), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_452), .A2(n_244), .B1(n_246), .B2(n_241), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_404), .A2(n_366), .B(n_364), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_409), .A2(n_248), .B1(n_249), .B2(n_247), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_409), .A2(n_366), .B1(n_383), .B2(n_364), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_422), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_415), .A2(n_245), .B1(n_259), .B2(n_253), .Y(n_518) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_421), .B(n_189), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_465), .B(n_4), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_431), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_440), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_443), .A2(n_268), .B1(n_282), .B2(n_266), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_423), .B(n_5), .Y(n_524) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_461), .A2(n_294), .B(n_283), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_445), .Y(n_526) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_460), .A2(n_306), .A3(n_317), .B(n_312), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_436), .A2(n_293), .B1(n_14), .B2(n_7), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_417), .A2(n_312), .B1(n_317), .B2(n_306), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_447), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_469), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_417), .A2(n_312), .B1(n_317), .B2(n_306), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_425), .A2(n_322), .B1(n_323), .B2(n_317), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_454), .Y(n_535) );
AO31x2_ASAP7_75t_L g536 ( .A1(n_456), .A2(n_323), .A3(n_326), .B(n_322), .Y(n_536) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_456), .A2(n_326), .A3(n_330), .B(n_323), .Y(n_537) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_406), .A2(n_330), .B(n_326), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_466), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_474), .Y(n_540) );
AOI21xp33_ASAP7_75t_L g541 ( .A1(n_432), .A2(n_13), .B(n_15), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_425), .A2(n_336), .B1(n_310), .B2(n_301), .C(n_299), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_413), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_475), .A2(n_80), .B(n_78), .Y(n_545) );
INVx4_ASAP7_75t_L g546 ( .A(n_411), .Y(n_546) );
OAI211xp5_ASAP7_75t_SL g547 ( .A1(n_493), .A2(n_459), .B(n_463), .C(n_472), .Y(n_547) );
BUFx10_ASAP7_75t_L g548 ( .A(n_511), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_488), .Y(n_549) );
BUFx3_ASAP7_75t_L g550 ( .A(n_539), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_488), .Y(n_551) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_505), .A2(n_434), .A3(n_453), .B(n_428), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_503), .B(n_512), .Y(n_553) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_481), .A2(n_470), .B(n_462), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_504), .A2(n_437), .B1(n_446), .B2(n_441), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_507), .A2(n_437), .B1(n_435), .B2(n_420), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_520), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_484), .A2(n_513), .B(n_510), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_540), .A2(n_435), .B1(n_426), .B2(n_301), .Y(n_559) );
CKINVDCx8_ASAP7_75t_R g560 ( .A(n_506), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_531), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
INVxp33_ASAP7_75t_L g563 ( .A(n_478), .Y(n_563) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_482), .A2(n_301), .B(n_299), .Y(n_564) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_525), .A2(n_541), .B(n_509), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_516), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_521), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_531), .B(n_22), .Y(n_569) );
AOI21xp33_ASAP7_75t_L g570 ( .A1(n_498), .A2(n_23), .B(n_24), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_494), .B(n_28), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_522), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_544), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_497), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_574) );
OA21x2_ASAP7_75t_L g575 ( .A1(n_529), .A2(n_83), .B(n_82), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_499), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_496), .A2(n_38), .B1(n_42), .B2(n_43), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_528), .A2(n_45), .B1(n_46), .B2(n_48), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_519), .A2(n_46), .B1(n_50), .B2(n_51), .Y(n_580) );
AO21x2_ASAP7_75t_L g581 ( .A1(n_525), .A2(n_86), .B(n_84), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_490), .B(n_52), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_491), .B(n_54), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_487), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_584) );
INVx6_ASAP7_75t_L g585 ( .A(n_500), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_487), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_535), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_536), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_495), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_536), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_489), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_591) );
HB1xp67_ASAP7_75t_SL g592 ( .A(n_495), .Y(n_592) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_529), .A2(n_94), .B(n_95), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_508), .B(n_97), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_476), .A2(n_98), .B1(n_99), .B2(n_101), .Y(n_595) );
OAI211xp5_ASAP7_75t_SL g596 ( .A1(n_479), .A2(n_106), .B(n_108), .C(n_109), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_480), .A2(n_110), .B(n_111), .Y(n_597) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_538), .A2(n_117), .B(n_118), .Y(n_598) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_532), .A2(n_120), .B(n_122), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_536), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_483), .Y(n_601) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_532), .A2(n_123), .B(n_126), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_485), .Y(n_603) );
BUFx3_ASAP7_75t_L g604 ( .A(n_492), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_514), .A2(n_131), .B1(n_135), .B2(n_136), .C(n_138), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_488), .Y(n_606) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_547), .A2(n_477), .B1(n_486), .B2(n_492), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_547), .A2(n_477), .B1(n_486), .B2(n_518), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_580), .B(n_523), .C(n_502), .Y(n_610) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_592), .Y(n_611) );
OA21x2_ASAP7_75t_L g612 ( .A1(n_558), .A2(n_543), .B(n_545), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_567), .B(n_527), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_553), .A2(n_542), .B1(n_530), .B2(n_534), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_572), .B(n_527), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_561), .B(n_527), .Y(n_618) );
INVx5_ASAP7_75t_L g619 ( .A(n_549), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_590), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_589), .B(n_501), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_563), .B(n_546), .Y(n_623) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_564), .A2(n_533), .B(n_515), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_600), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_554), .Y(n_626) );
AO21x2_ASAP7_75t_L g627 ( .A1(n_565), .A2(n_537), .B(n_536), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_551), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_551), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_577), .B(n_537), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_587), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_551), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_568), .B(n_143), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_606), .B(n_145), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_573), .B(n_148), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_606), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_601), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_603), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_552), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_603), .B(n_159), .Y(n_640) );
NAND2xp33_ASAP7_75t_R g641 ( .A(n_575), .B(n_162), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_552), .Y(n_642) );
NOR2xp33_ASAP7_75t_SL g643 ( .A(n_560), .B(n_548), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_552), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_557), .B(n_562), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_583), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_569), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_579), .A2(n_571), .B1(n_570), .B2(n_574), .C(n_576), .Y(n_648) );
BUFx2_ASAP7_75t_L g649 ( .A(n_604), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_582), .Y(n_650) );
INVx3_ASAP7_75t_L g651 ( .A(n_585), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_594), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_575), .Y(n_653) );
OAI31xp33_ASAP7_75t_L g654 ( .A1(n_578), .A2(n_591), .A3(n_586), .B(n_584), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_552), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_581), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_598), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_594), .Y(n_658) );
OA21x2_ASAP7_75t_L g659 ( .A1(n_599), .A2(n_602), .B(n_597), .Y(n_659) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_595), .A2(n_605), .A3(n_596), .B(n_550), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_598), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_613), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_630), .B(n_593), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_619), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_630), .B(n_555), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_613), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_616), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_617), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_616), .B(n_555), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_638), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_617), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_618), .B(n_556), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_620), .Y(n_673) );
INVx4_ASAP7_75t_L g674 ( .A(n_619), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_620), .Y(n_675) );
INVx3_ASAP7_75t_L g676 ( .A(n_619), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_618), .B(n_559), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_639), .B(n_642), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_625), .B(n_631), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_625), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_615), .A2(n_648), .B1(n_609), .B2(n_647), .C(n_660), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_639), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_621), .B(n_645), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_645), .B(n_627), .Y(n_684) );
AOI33xp33_ASAP7_75t_L g685 ( .A1(n_646), .A2(n_650), .A3(n_637), .B1(n_608), .B2(n_658), .B3(n_652), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_627), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_642), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_644), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_627), .B(n_655), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_611), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_649), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_632), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_626), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_643), .B(n_654), .C(n_623), .D(n_610), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_622), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_653), .Y(n_697) );
INVx4_ASAP7_75t_L g698 ( .A(n_619), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_633), .B(n_635), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_614), .B(n_629), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_614), .B(n_629), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_607), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_619), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_640), .B(n_651), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_636), .B(n_651), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_653), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_636), .B(n_656), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_607), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_671), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_683), .B(n_636), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_695), .B(n_641), .C(n_634), .D(n_661), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_684), .B(n_657), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_684), .B(n_657), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_662), .B(n_612), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_668), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_666), .B(n_612), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_666), .B(n_612), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_667), .B(n_624), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_668), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_667), .B(n_624), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_671), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_681), .B(n_659), .C(n_624), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_673), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_679), .B(n_628), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_664), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_682), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_672), .B(n_659), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_682), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_670), .B(n_696), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_665), .B(n_669), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_687), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_687), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_672), .B(n_680), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_685), .B(n_692), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_690), .B(n_663), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_688), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_690), .B(n_663), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_688), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_680), .B(n_677), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_675), .B(n_678), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_677), .B(n_692), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_675), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_689), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_689), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_699), .B(n_704), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_678), .B(n_686), .Y(n_746) );
BUFx3_ASAP7_75t_L g747 ( .A(n_676), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_686), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_741), .B(n_697), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_729), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_735), .B(n_706), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_737), .B(n_706), .Y(n_752) );
AND2x2_ASAP7_75t_SL g753 ( .A(n_725), .B(n_691), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_709), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_743), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_737), .B(n_678), .Y(n_756) );
NOR2x1p5_ASAP7_75t_L g757 ( .A(n_711), .B(n_698), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_741), .B(n_707), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g759 ( .A1(n_734), .A2(n_705), .B1(n_674), .B2(n_698), .C(n_703), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_730), .B(n_713), .Y(n_760) );
AND2x2_ASAP7_75t_SL g761 ( .A(n_725), .B(n_674), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_709), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_722), .B(n_701), .C(n_700), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_721), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_721), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_723), .Y(n_766) );
NAND4xp25_ASAP7_75t_L g767 ( .A(n_745), .B(n_707), .C(n_693), .D(n_694), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_724), .Y(n_768) );
NOR2xp33_ASAP7_75t_SL g769 ( .A(n_747), .B(n_708), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_733), .B(n_702), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_760), .B(n_740), .Y(n_771) );
INVx3_ASAP7_75t_SL g772 ( .A(n_761), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_754), .Y(n_773) );
AOI21xp33_ASAP7_75t_SL g774 ( .A1(n_753), .A2(n_739), .B(n_710), .Y(n_774) );
AOI222xp33_ASAP7_75t_L g775 ( .A1(n_750), .A2(n_717), .B1(n_716), .B2(n_714), .C1(n_720), .C2(n_718), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_756), .B(n_740), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_754), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_756), .B(n_727), .Y(n_778) );
NAND2x1p5_ASAP7_75t_L g779 ( .A(n_757), .B(n_726), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_755), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_755), .Y(n_781) );
INVx2_ASAP7_75t_SL g782 ( .A(n_768), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_762), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_751), .B(n_746), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_752), .B(n_712), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_764), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_763), .A2(n_731), .B1(n_744), .B2(n_738), .C1(n_736), .C2(n_732), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_759), .A2(n_728), .B1(n_732), .B2(n_731), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_765), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_766), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_758), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_758), .Y(n_792) );
AND2x2_ASAP7_75t_SL g793 ( .A(n_769), .B(n_715), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_L g794 ( .A1(n_767), .A2(n_748), .B(n_719), .C(n_742), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_749), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_777), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_771), .B(n_778), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_772), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_779), .A2(n_794), .B1(n_788), .B2(n_775), .C(n_787), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g800 ( .A(n_793), .B(n_774), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_773), .Y(n_801) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_798), .A2(n_782), .B(n_793), .C(n_795), .Y(n_802) );
AO22x2_ASAP7_75t_L g803 ( .A1(n_800), .A2(n_792), .B1(n_791), .B2(n_790), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g804 ( .A(n_799), .B(n_783), .C(n_786), .Y(n_804) );
NAND4xp25_ASAP7_75t_L g805 ( .A(n_797), .B(n_770), .C(n_785), .D(n_784), .Y(n_805) );
AOI221x1_ASAP7_75t_L g806 ( .A1(n_804), .A2(n_801), .B1(n_796), .B2(n_789), .C(n_783), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_803), .Y(n_807) );
NOR2x1_ASAP7_75t_L g808 ( .A(n_807), .B(n_802), .Y(n_808) );
OAI22x1_ASAP7_75t_L g809 ( .A1(n_808), .A2(n_806), .B1(n_805), .B2(n_776), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_809), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_810), .Y(n_811) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_811), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g813 ( .A1(n_812), .A2(n_780), .B(n_781), .Y(n_813) );
endmodule