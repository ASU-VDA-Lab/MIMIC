module fake_jpeg_29965_n_373 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_373);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_373;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_55),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_16),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_66),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_22),
.B(n_0),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_29),
.B(n_0),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_17),
.B1(n_41),
.B2(n_39),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_87),
.B1(n_91),
.B2(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_17),
.B1(n_41),
.B2(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_17),
.B1(n_39),
.B2(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_88),
.A2(n_111),
.B1(n_18),
.B2(n_47),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_104),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_99),
.A2(n_107),
.B1(n_115),
.B2(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_35),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_27),
.B1(n_31),
.B2(n_43),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_43),
.B1(n_37),
.B2(n_38),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_43),
.B1(n_37),
.B2(n_38),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_54),
.A2(n_42),
.B1(n_36),
.B2(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_36),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_33),
.Y(n_133)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_34),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_34),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_42),
.B1(n_40),
.B2(n_19),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_133),
.Y(n_172)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_64),
.B(n_19),
.C(n_56),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_131),
.Y(n_192)
);

CKINVDCx11_ASAP7_75t_R g129 ( 
.A(n_94),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_129),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_137),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_14),
.B(n_7),
.C(n_11),
.Y(n_131)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_33),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_8),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_144),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_96),
.B(n_50),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_59),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_87),
.B1(n_81),
.B2(n_103),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_149),
.B(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_23),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_153),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_53),
.B1(n_52),
.B2(n_48),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_166),
.B1(n_78),
.B2(n_18),
.Y(n_185)
);

AND2x4_ASAP7_75t_SL g149 ( 
.A(n_90),
.B(n_107),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_23),
.B1(n_33),
.B2(n_18),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_98),
.Y(n_153)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_69),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_23),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_163),
.Y(n_168)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

FAx1_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_100),
.CI(n_101),
.CON(n_162),
.SN(n_162)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_92),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_94),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_121),
.B1(n_82),
.B2(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_164),
.A2(n_145),
.B1(n_152),
.B2(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_106),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_113),
.B1(n_121),
.B2(n_80),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_175),
.B1(n_199),
.B2(n_155),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_80),
.B1(n_102),
.B2(n_82),
.Y(n_175)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_188),
.B1(n_191),
.B2(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_23),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_92),
.B(n_100),
.C(n_46),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_183),
.A2(n_155),
.B(n_159),
.C(n_150),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_185),
.A2(n_204),
.B1(n_5),
.B2(n_6),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_46),
.B1(n_108),
.B2(n_23),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g190 ( 
.A(n_127),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_140),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_1),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_203),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_130),
.B(n_1),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_149),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_143),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_216),
.C(n_171),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_149),
.B1(n_144),
.B2(n_131),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_211),
.B(n_213),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_212),
.A2(n_236),
.B1(n_237),
.B2(n_171),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_143),
.C(n_128),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_142),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_217),
.B(n_219),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_148),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_139),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_220),
.B(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_135),
.B1(n_154),
.B2(n_161),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_238),
.B1(n_195),
.B2(n_202),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_157),
.B1(n_151),
.B2(n_126),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_193),
.B(n_181),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_134),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_230),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_148),
.B(n_4),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_192),
.B(n_183),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_173),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_SL g231 ( 
.A(n_192),
.B(n_186),
.C(n_184),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_231),
.A2(n_186),
.B(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_2),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_234),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_235),
.A2(n_178),
.B1(n_6),
.B2(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_173),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_176),
.B1(n_196),
.B2(n_184),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_258),
.B1(n_264),
.B2(n_257),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_242),
.B(n_223),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_257),
.B(n_223),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_197),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_259),
.C(n_215),
.Y(n_282)
);

AO22x2_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_183),
.B1(n_171),
.B2(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_227),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_260),
.B1(n_235),
.B2(n_232),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_189),
.B(n_167),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_255),
.B(n_229),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_217),
.B(n_177),
.CI(n_193),
.CON(n_254),
.SN(n_254)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_254),
.B(n_223),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_216),
.A2(n_189),
.B(n_181),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_205),
.A2(n_177),
.B1(n_178),
.B2(n_5),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_177),
.C(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_209),
.C(n_205),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_283),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_269),
.B(n_284),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_278),
.B(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_206),
.Y(n_271)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_214),
.Y(n_273)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_226),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_282),
.C(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_281),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_207),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_210),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_280),
.B(n_285),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_221),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_290),
.B1(n_264),
.B2(n_241),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_236),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_248),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_289),
.B1(n_246),
.B2(n_248),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_233),
.B1(n_225),
.B2(n_222),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_239),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_242),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_288),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_255),
.C(n_266),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_252),
.C(n_246),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_246),
.C(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_306),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_308),
.B1(n_277),
.B2(n_289),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_244),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_248),
.C(n_241),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_250),
.B1(n_260),
.B2(n_243),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_268),
.C(n_284),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_307),
.Y(n_315)
);

NAND5xp2_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_285),
.C(n_280),
.D(n_283),
.E(n_270),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_322),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_294),
.A2(n_288),
.B(n_278),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_316),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_279),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_324),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_296),
.A2(n_281),
.A3(n_290),
.B1(n_273),
.B2(n_271),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_293),
.C(n_306),
.Y(n_334)
);

BUFx12f_ASAP7_75t_SL g324 ( 
.A(n_297),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_325),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_303),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_291),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_337),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_339),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_311),
.C(n_318),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_299),
.C(n_300),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_305),
.C(n_313),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_333),
.A2(n_324),
.B(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_346),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_333),
.A2(n_314),
.B(n_321),
.Y(n_343)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_343),
.Y(n_355)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_322),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_312),
.B(n_340),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_328),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_249),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_347),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_307),
.C(n_327),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_348),
.B(n_350),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_325),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_357),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_344),
.A2(n_330),
.B1(n_340),
.B2(n_338),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_353),
.A2(n_272),
.B1(n_263),
.B2(n_256),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_354),
.A2(n_359),
.B(n_276),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_345),
.B(n_323),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_298),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_341),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_360),
.A2(n_263),
.B(n_261),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_359),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_355),
.A2(n_346),
.B1(n_243),
.B2(n_256),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_353),
.Y(n_365)
);

AOI322xp5_ASAP7_75t_L g367 ( 
.A1(n_365),
.A2(n_354),
.A3(n_356),
.B1(n_358),
.B2(n_274),
.C1(n_352),
.C2(n_251),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_368),
.Y(n_369)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_364),
.A3(n_274),
.B1(n_365),
.B2(n_261),
.C1(n_262),
.C2(n_360),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_370),
.A2(n_262),
.B(n_218),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_369),
.B(n_218),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_372),
.B(n_218),
.Y(n_373)
);


endmodule