module fake_jpeg_6687_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_50),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_7),
.CON(n_50),
.SN(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_7),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_54),
.B(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_1),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_64),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_28),
.B(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_37),
.B1(n_23),
.B2(n_26),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_74),
.B1(n_41),
.B2(n_34),
.Y(n_116)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_37),
.B1(n_23),
.B2(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_37),
.B(n_38),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_90),
.B(n_105),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_77),
.B(n_79),
.Y(n_138)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_31),
.B(n_38),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_12),
.Y(n_143)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_83),
.B(n_93),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_17),
.B1(n_16),
.B2(n_26),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_84),
.A2(n_85),
.B1(n_102),
.B2(n_75),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_16),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_35),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_19),
.B1(n_34),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_112),
.B1(n_14),
.B2(n_13),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_106),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_16),
.B1(n_21),
.B2(n_32),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_44),
.A2(n_13),
.B(n_15),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_109),
.Y(n_150)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_1),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_47),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_127),
.B1(n_146),
.B2(n_113),
.Y(n_184)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_70),
.A2(n_41),
.B1(n_30),
.B2(n_27),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_142),
.B1(n_111),
.B2(n_101),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_71),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_123),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_146),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_126),
.B(n_136),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_30),
.B1(n_6),
.B2(n_11),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_129),
.Y(n_167)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_131),
.A2(n_132),
.B1(n_109),
.B2(n_106),
.Y(n_179)
);

BUFx8_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_98),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_140),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_92),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_90),
.B1(n_105),
.B2(n_101),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_3),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_78),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_155),
.Y(n_203)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g213 ( 
.A(n_158),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_92),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_178),
.Y(n_188)
);

OAI22x1_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_76),
.B1(n_67),
.B2(n_100),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_163),
.B1(n_182),
.B2(n_185),
.Y(n_193)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_165),
.Y(n_209)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_169),
.B1(n_184),
.B2(n_119),
.Y(n_199)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_170),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_68),
.B1(n_67),
.B2(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_103),
.Y(n_216)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_177),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_67),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_123),
.Y(n_189)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_143),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_108),
.B1(n_99),
.B2(n_100),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_135),
.B1(n_126),
.B2(n_120),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_78),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_190),
.B1(n_194),
.B2(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_197),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_120),
.B1(n_121),
.B2(n_149),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_121),
.B1(n_119),
.B2(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_207),
.B1(n_205),
.B2(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_117),
.B(n_136),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_215),
.B(n_158),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_139),
.B1(n_117),
.B2(n_130),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_205),
.A2(n_221),
.B1(n_156),
.B2(n_118),
.Y(n_247)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_216),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_130),
.B1(n_99),
.B2(n_134),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_214),
.B1(n_186),
.B2(n_162),
.Y(n_233)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_151),
.A2(n_134),
.B1(n_82),
.B2(n_103),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_3),
.B(n_4),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_4),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_82),
.B1(n_5),
.B2(n_118),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_160),
.C(n_152),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_245),
.C(n_204),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_200),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_230),
.B(n_244),
.Y(n_255)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_229),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_168),
.B(n_170),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_218),
.B1(n_208),
.B2(n_197),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_175),
.B1(n_172),
.B2(n_182),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_246),
.B1(n_193),
.B2(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_247),
.B1(n_214),
.B2(n_189),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_191),
.B(n_216),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_189),
.C(n_172),
.Y(n_240)
);

BUFx12f_ASAP7_75t_SL g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_206),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_178),
.B(n_154),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_165),
.C(n_157),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_174),
.B1(n_155),
.B2(n_156),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_265),
.B1(n_247),
.B2(n_270),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_259),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_262),
.C(n_264),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_260),
.B(n_266),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_199),
.C(n_194),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_192),
.B(n_202),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_231),
.B1(n_242),
.B2(n_226),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_215),
.B(n_208),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_227),
.B1(n_235),
.B2(n_246),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_281),
.B1(n_264),
.B2(n_257),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_280),
.C(n_283),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

AOI31xp67_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_255),
.A3(n_263),
.B(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_228),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_267),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_282),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_255),
.A2(n_227),
.B1(n_231),
.B2(n_248),
.Y(n_281)
);

HB1xp67_ASAP7_75t_SL g283 ( 
.A(n_258),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_248),
.B1(n_190),
.B2(n_211),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_262),
.B1(n_268),
.B2(n_266),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_244),
.C(n_196),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_228),
.C(n_236),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_296),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_294),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_261),
.B1(n_269),
.B2(n_250),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_261),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_229),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_287),
.C(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_284),
.B1(n_276),
.B2(n_282),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_311),
.C(n_312),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_274),
.C(n_279),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_281),
.C(n_272),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_280),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_254),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_301),
.B1(n_300),
.B2(n_289),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_271),
.B1(n_288),
.B2(n_292),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_305),
.B1(n_304),
.B2(n_303),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_297),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_285),
.B1(n_292),
.B2(n_250),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_321),
.B1(n_252),
.B2(n_118),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_241),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_325),
.B1(n_318),
.B2(n_316),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_254),
.C(n_223),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_320),
.B(n_317),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_330),
.B(n_331),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_313),
.Y(n_331)
);

OAI321xp33_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_326),
.A3(n_324),
.B1(n_323),
.B2(n_314),
.C(n_133),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_330),
.C(n_328),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_333),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_133),
.Y(n_337)
);


endmodule