module fake_jpeg_13435_n_180 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_0),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_74),
.Y(n_96)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_2),
.Y(n_91)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_3),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_75),
.B1(n_64),
.B2(n_59),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_60),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_51),
.B1(n_65),
.B2(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_4),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_65),
.B1(n_51),
.B2(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_71),
.B1(n_62),
.B2(n_57),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_52),
.B1(n_56),
.B2(n_63),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_99),
.B(n_60),
.C(n_54),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_49),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_50),
.C(n_55),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_6),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_119),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_4),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_9),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_34),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_77),
.Y(n_119)
);

NOR2x1_ASAP7_75t_R g128 ( 
.A(n_121),
.B(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_54),
.B1(n_7),
.B2(n_9),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_127),
.B(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_120),
.B1(n_108),
.B2(n_118),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_131),
.Y(n_157)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_38),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_11),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_13),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_19),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_39),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_145),
.B1(n_151),
.B2(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_36),
.C(n_37),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_149),
.B(n_153),
.C(n_147),
.D(n_45),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_130),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_156),
.C(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_137),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_161),
.B(n_166),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_129),
.B1(n_134),
.B2(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_154),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_170),
.B1(n_136),
.B2(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_168),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_173),
.B(n_165),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_167),
.B1(n_171),
.B2(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_157),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_144),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);


endmodule