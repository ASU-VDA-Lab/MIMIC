module fake_jpeg_23015_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_44;
wire n_28;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_13),
.A2(n_15),
.B1(n_14),
.B2(n_18),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_12),
.Y(n_32)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_16),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_11),
.B(n_16),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_46),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_20),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_29),
.C(n_9),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_34),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_31),
.C(n_41),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_46),
.B(n_40),
.Y(n_56)
);

AO22x1_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_42),
.B1(n_31),
.B2(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

OAI221xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_52),
.B1(n_47),
.B2(n_48),
.C(n_21),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_60),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_51),
.B(n_21),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_58),
.C(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_20),
.C(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_3),
.B1(n_4),
.B2(n_20),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_3),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_72),
.B(n_73),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_71),
.Y(n_76)
);


endmodule