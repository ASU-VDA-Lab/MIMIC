module fake_jpeg_6294_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_24),
.Y(n_40)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_32),
.B1(n_35),
.B2(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_45),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_46),
.B1(n_48),
.B2(n_14),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_27),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_47),
.C(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_20),
.B2(n_17),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_22),
.B(n_17),
.C(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_60)
);

AOI31xp67_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_38),
.A3(n_10),
.B(n_3),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_43),
.B1(n_31),
.B2(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_29),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_53),
.B1(n_58),
.B2(n_32),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_43),
.C(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_32),
.B1(n_28),
.B2(n_14),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_49),
.B1(n_53),
.B2(n_55),
.C(n_5),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_77),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_52),
.B(n_49),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_77),
.B1(n_71),
.B2(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_60),
.B(n_67),
.C(n_64),
.D(n_61),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_75),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_38),
.C(n_2),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_74),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_1),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_93),
.B1(n_79),
.B2(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_91),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_38),
.B(n_2),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_69),
.B1(n_32),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_86),
.B1(n_84),
.B2(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_96),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_98),
.B(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_89),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_1),
.C(n_4),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_90),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_101),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_107),
.C(n_4),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_4),
.B(n_7),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_8),
.C(n_9),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_8),
.B(n_9),
.Y(n_110)
);


endmodule