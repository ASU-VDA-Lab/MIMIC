module fake_jpeg_8117_n_291 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_16),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_18),
.B(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g38 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_21),
.B(n_35),
.C(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_34),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_20),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_51),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_55),
.B1(n_65),
.B2(n_19),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_21),
.B(n_22),
.C(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_62),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_19),
.B1(n_30),
.B2(n_34),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_31),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_29),
.B1(n_34),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_70),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_83),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_20),
.B(n_24),
.C(n_27),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_88),
.B1(n_19),
.B2(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_87),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_18),
.B(n_26),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_90),
.B(n_91),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_17),
.C(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_94),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_24),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_109),
.B1(n_86),
.B2(n_70),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_106),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_60),
.B1(n_47),
.B2(n_54),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_101),
.B1(n_78),
.B2(n_75),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_100),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_18),
.B(n_32),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_19),
.B1(n_56),
.B2(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_112),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_115),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_116),
.B1(n_120),
.B2(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_64),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_95),
.B1(n_109),
.B2(n_102),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_125),
.B1(n_142),
.B2(n_98),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_86),
.B1(n_78),
.B2(n_90),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_83),
.C(n_77),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_128),
.C(n_137),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_73),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_138),
.B(n_150),
.C(n_99),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_81),
.C(n_74),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_101),
.C(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_149),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_81),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_74),
.B(n_87),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_45),
.B(n_74),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_141),
.B(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_84),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_1),
.Y(n_141)
);

OAI22x1_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_72),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_72),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_67),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_67),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_45),
.B(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_151),
.B(n_153),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_112),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_167),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_124),
.B1(n_135),
.B2(n_142),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_163),
.B(n_26),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_119),
.C(n_107),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_168),
.C(n_176),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_98),
.B1(n_115),
.B2(n_107),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_165),
.B1(n_178),
.B2(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_103),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_175),
.Y(n_187)
);

NOR4xp25_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_103),
.C(n_100),
.D(n_108),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_108),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_82),
.C(n_45),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_53),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_139),
.C(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_24),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_191),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_189),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_135),
.B(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_123),
.B1(n_133),
.B2(n_138),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_133),
.B1(n_138),
.B2(n_134),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_196),
.C(n_199),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_131),
.B1(n_141),
.B2(n_147),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_197),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_79),
.B1(n_71),
.B2(n_32),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_203),
.B1(n_204),
.B2(n_2),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_53),
.C(n_79),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_79),
.C(n_71),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_203),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_161),
.C(n_168),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_213),
.C(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_215),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_151),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_172),
.C(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_162),
.B1(n_166),
.B2(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_192),
.B1(n_5),
.B2(n_6),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_218),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_17),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_17),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_10),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_191),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_241),
.B(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_196),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_238),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_199),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_182),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_219),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_205),
.B(n_206),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_249),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_227),
.A2(n_222),
.B1(n_192),
.B2(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_241),
.B1(n_233),
.B2(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_229),
.A2(n_223),
.B1(n_222),
.B2(n_221),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_250),
.B1(n_232),
.B2(n_236),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_248),
.B(n_237),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_225),
.B(n_5),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_10),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_3),
.C(n_6),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_259),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_7),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_250),
.C(n_253),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_230),
.C(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_246),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_240),
.C(n_239),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_262),
.C(n_245),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_12),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_270),
.C(n_273),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_249),
.C(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_3),
.C(n_9),
.Y(n_273)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_254),
.B1(n_257),
.B2(n_255),
.C(n_262),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_273),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_12),
.B(n_13),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_13),
.C(n_15),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_16),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_269),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_278),
.C(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_287),
.C(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_285),
.C(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_270),
.Y(n_291)
);


endmodule