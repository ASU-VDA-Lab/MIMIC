module fake_jpeg_13255_n_83 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_3),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_5),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_30),
.Y(n_51)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_43),
.A3(n_29),
.B1(n_25),
.B2(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_56),
.B(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_58),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_28),
.CON(n_56),
.SN(n_56)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_36),
.B(n_42),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_62),
.B1(n_8),
.B2(n_10),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_4),
.B(n_5),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_6),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_15),
.C(n_18),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_71),
.C(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_21),
.B(n_22),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_64),
.B(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_69),
.C(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_72),
.B(n_75),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_71),
.B(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_57),
.Y(n_83)
);


endmodule