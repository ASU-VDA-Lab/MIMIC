module fake_jpeg_6447_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

AND2x2_ASAP7_75t_L g5 ( 
.A(n_2),
.B(n_3),
.Y(n_5)
);

INVx6_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

AOI322xp5_ASAP7_75t_L g10 ( 
.A1(n_9),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_0),
.C1(n_1),
.C2(n_2),
.Y(n_10)
);

OA21x2_ASAP7_75t_SL g11 ( 
.A1(n_10),
.A2(n_0),
.B(n_6),
.Y(n_11)
);


endmodule