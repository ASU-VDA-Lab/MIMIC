module fake_jpeg_19319_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_20),
.B(n_19),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_37),
.B(n_38),
.C(n_36),
.Y(n_80)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_21),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_31),
.B1(n_32),
.B2(n_30),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_62),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_63),
.B(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_48),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_0),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_25),
.B1(n_29),
.B2(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_20),
.B1(n_33),
.B2(n_24),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_88),
.B1(n_52),
.B2(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_23),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_30),
.B1(n_16),
.B2(n_2),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_77),
.B1(n_82),
.B2(n_91),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_30),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_117),
.Y(n_132)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_0),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_86),
.Y(n_128)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_7),
.C(n_14),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_63),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_1),
.B(n_2),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_60),
.B(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_147),
.B(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_84),
.B1(n_73),
.B2(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_128),
.Y(n_157)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_112),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_92),
.B1(n_65),
.B2(n_67),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_142),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_72),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_143),
.B(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_98),
.A2(n_93),
.B1(n_94),
.B2(n_74),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_150),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_151),
.B1(n_103),
.B2(n_114),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_64),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_65),
.B1(n_64),
.B2(n_75),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_120),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_88),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_89),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_115),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_155),
.B(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_114),
.B1(n_96),
.B2(n_118),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_123),
.B(n_98),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_165),
.B(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_160),
.B(n_186),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_105),
.B1(n_99),
.B2(n_107),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_168),
.B1(n_141),
.B2(n_117),
.Y(n_192)
);

XOR2x2_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_132),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_147),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_103),
.B(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_133),
.A2(n_107),
.B1(n_119),
.B2(n_101),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_107),
.B(n_111),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_173),
.A2(n_1),
.B(n_3),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_174),
.B(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_109),
.Y(n_177)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_117),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_152),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_121),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_168),
.Y(n_224)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_171),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_161),
.B1(n_169),
.B2(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_106),
.B1(n_136),
.B2(n_114),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_213),
.B1(n_216),
.B2(n_187),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_145),
.B(n_108),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_202),
.B(n_215),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_200),
.B(n_214),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_108),
.B(n_131),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_174),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_176),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_145),
.C(n_102),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_210),
.C(n_171),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_96),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_10),
.C(n_14),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_187),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_15),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_10),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_160),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_178),
.B1(n_201),
.B2(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_232),
.B1(n_238),
.B2(n_199),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_164),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_164),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_162),
.B1(n_163),
.B2(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_234),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_166),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_237),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_155),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_179),
.C(n_172),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_206),
.C(n_208),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_189),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_210),
.C(n_192),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_247),
.C(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_195),
.C(n_202),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_185),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_239),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_194),
.C(n_198),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_261),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_203),
.C(n_179),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_233),
.C(n_232),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_223),
.B(n_228),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_241),
.C(n_233),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_273),
.C(n_246),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_223),
.B(n_231),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_220),
.B1(n_221),
.B2(n_205),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_275),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_220),
.B(n_215),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_238),
.C(n_190),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_244),
.A2(n_205),
.B(n_212),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_159),
.B1(n_209),
.B2(n_180),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_185),
.B1(n_5),
.B2(n_6),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_256),
.C(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_290),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_253),
.C(n_249),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_263),
.B(n_269),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_255),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_255),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_265),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_299),
.C(n_281),
.Y(n_310)
);

AOI31xp33_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_300),
.A3(n_285),
.B(n_280),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_276),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_301),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_262),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_270),
.B(n_271),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_11),
.B(n_5),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_277),
.B(n_270),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_288),
.B(n_262),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_306),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_287),
.B1(n_286),
.B2(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_312),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_301),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_278),
.B(n_275),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_311),
.B(n_4),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_298),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_296),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_293),
.B(n_306),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_5),
.C(n_6),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.C(n_320),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_5),
.B(n_6),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_317),
.B(n_316),
.C(n_6),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_317),
.Y(n_324)
);


endmodule