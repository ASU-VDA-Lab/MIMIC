module real_jpeg_29499_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_244;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_10),
.B(n_61),
.C(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_67),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_4),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_5),
.A2(n_25),
.B1(n_29),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_48),
.B1(n_57),
.B2(n_58),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_7),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_97),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_97),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_7),
.A2(n_25),
.B1(n_29),
.B2(n_97),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_25),
.B1(n_29),
.B2(n_40),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_9),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_10),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_55),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_38),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_10),
.A2(n_38),
.B(n_42),
.C(n_202),
.D(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_71),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_10),
.A2(n_24),
.B(n_215),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_10),
.A2(n_58),
.B(n_70),
.C(n_152),
.D(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_10),
.B(n_58),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_38),
.B(n_43),
.C(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_25),
.B1(n_29),
.B2(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_12),
.A2(n_25),
.B1(n_29),
.B2(n_64),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_64),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_13),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_77),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_77),
.Y(n_190)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_74),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_88),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_21),
.B(n_81),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_51),
.B2(n_80),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_23),
.B(n_36),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_28),
.B1(n_33),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_24),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_24),
.A2(n_31),
.B1(n_146),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_24),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_24),
.B(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_25),
.B(n_44),
.Y(n_203)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_29),
.A2(n_39),
.A3(n_45),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_29),
.B(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_31),
.A2(n_222),
.B(n_230),
.Y(n_229)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_32),
.A2(n_92),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_32),
.B(n_216),
.Y(n_215)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_33),
.B(n_141),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_39),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g251 ( 
.A1(n_38),
.A2(n_57),
.A3(n_244),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g253 ( 
.A(n_39),
.B(n_73),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_41),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_46),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_46),
.B1(n_85),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_42),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_42),
.A2(n_46),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_49),
.A2(n_94),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_49),
.B(n_168),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_49),
.A2(n_166),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_49),
.B(n_141),
.Y(n_228)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_68),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_52),
.B(n_68),
.C(n_80),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B(n_65),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_54),
.B(n_66),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_54),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_56),
.A2(n_58),
.B(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_SL g58 ( 
.A(n_57),
.Y(n_58)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_65),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_69),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_70),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_71),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_70),
.A2(n_71),
.B1(n_150),
.B2(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_73),
.Y(n_252)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_78),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_78),
.B(n_102),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_78),
.A2(n_100),
.B(n_174),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_87),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_87),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.C(n_98),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_93),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_123),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_112),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_120),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_155),
.B(n_274),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_153),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_128),
.B(n_153),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_132),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_134),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_147),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_147),
.B2(n_148),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_144),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_194),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_193),
.Y(n_157)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_159),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_172),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_165),
.B1(n_172),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_179),
.B(n_181),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_185),
.B(n_187),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_188),
.B(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_190),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_272),
.C(n_273),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_267),
.B(n_271),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_255),
.B(n_266),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_239),
.B(n_254),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_218),
.B(n_238),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_206),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_204),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_205),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B(n_237),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_225),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_231),
.B(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_232),
.B(n_236),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_241),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);


endmodule