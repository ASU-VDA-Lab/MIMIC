module fake_jpeg_12143_n_628 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_628);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_628;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_2),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_62),
.B(n_95),
.Y(n_153)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_76),
.B(n_91),
.Y(n_146)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_79),
.Y(n_207)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_81),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g178 ( 
.A(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_36),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_101),
.Y(n_132)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_86),
.Y(n_127)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_87),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_36),
.B(n_10),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_14),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_53),
.B(n_15),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_103),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_14),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_109),
.B(n_111),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_14),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_114),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_119),
.Y(n_203)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g206 ( 
.A(n_121),
.Y(n_206)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_38),
.Y(n_125)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_125),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_31),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_51),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_60),
.A2(n_29),
.B1(n_24),
.B2(n_41),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_138),
.A2(n_143),
.B1(n_144),
.B2(n_160),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_51),
.B1(n_53),
.B2(n_34),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_64),
.A2(n_51),
.B1(n_56),
.B2(n_28),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_37),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_42),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_156),
.B(n_186),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_24),
.B1(n_41),
.B2(n_30),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_157),
.A2(n_197),
.B1(n_209),
.B2(n_194),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_65),
.A2(n_21),
.B1(n_56),
.B2(n_44),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_35),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_191),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_105),
.A2(n_40),
.B1(n_35),
.B2(n_43),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_177),
.B1(n_126),
.B2(n_123),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_69),
.A2(n_28),
.B1(n_44),
.B2(n_21),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_93),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_179),
.A2(n_52),
.B(n_38),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_111),
.B(n_33),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_59),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_188),
.B(n_189),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_59),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_82),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_190),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_86),
.B(n_59),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_59),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_192),
.B(n_195),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_97),
.B(n_18),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_110),
.A2(n_41),
.B1(n_37),
.B2(n_30),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_99),
.B(n_37),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_204),
.B(n_13),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_72),
.B(n_33),
.C(n_18),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_103),
.C(n_115),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_211),
.A2(n_229),
.B1(n_247),
.B2(n_257),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_217),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_131),
.B(n_37),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_214),
.B(n_222),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_144),
.A2(n_94),
.B1(n_107),
.B2(n_102),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_215),
.A2(n_221),
.B1(n_226),
.B2(n_268),
.Y(n_320)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_147),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_160),
.A2(n_92),
.B1(n_81),
.B2(n_100),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_134),
.B(n_0),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_0),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_223),
.B(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_85),
.B1(n_73),
.B2(n_98),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_227),
.A2(n_240),
.B(n_238),
.Y(n_326)
);

AOI32xp33_ASAP7_75t_L g228 ( 
.A1(n_146),
.A2(n_99),
.A3(n_113),
.B1(n_116),
.B2(n_88),
.Y(n_228)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_228),
.A2(n_237),
.A3(n_241),
.B1(n_247),
.B2(n_212),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_138),
.A2(n_52),
.B1(n_38),
.B2(n_3),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_158),
.A2(n_153),
.B1(n_157),
.B2(n_127),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_230),
.A2(n_243),
.B1(n_265),
.B2(n_281),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_147),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_152),
.Y(n_235)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_168),
.A2(n_190),
.B(n_128),
.Y(n_236)
);

BUFx24_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_170),
.A2(n_38),
.B(n_52),
.C(n_11),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_169),
.Y(n_239)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_182),
.A2(n_52),
.B1(n_15),
.B2(n_13),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_129),
.B(n_0),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_241),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_136),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_242),
.B(n_259),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_127),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_245),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_176),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_SL g248 ( 
.A1(n_136),
.A2(n_11),
.B(n_12),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_254),
.C(n_274),
.Y(n_298)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_154),
.Y(n_249)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_184),
.B(n_4),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_167),
.A2(n_5),
.B1(n_6),
.B2(n_15),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_132),
.B(n_166),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_142),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_267),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_178),
.Y(n_301)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_133),
.B(n_6),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_164),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_264),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_142),
.A2(n_6),
.B1(n_12),
.B2(n_145),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_196),
.A2(n_208),
.B1(n_167),
.B2(n_165),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_266),
.A2(n_209),
.B1(n_148),
.B2(n_198),
.Y(n_308)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_145),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_133),
.A2(n_185),
.B1(n_159),
.B2(n_166),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_155),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_178),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_272),
.Y(n_321)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_140),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_273),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_174),
.B(n_193),
.Y(n_274)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_275),
.Y(n_323)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_279),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_150),
.B(n_137),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_207),
.Y(n_313)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_139),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_163),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_213),
.Y(n_339)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_163),
.Y(n_281)
);

OA22x2_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_194),
.B1(n_185),
.B2(n_159),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_301),
.B(n_338),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_282),
.A2(n_148),
.B1(n_165),
.B2(n_198),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_318),
.B1(n_327),
.B2(n_281),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_229),
.A2(n_152),
.B1(n_139),
.B2(n_187),
.Y(n_303)
);

OAI22x1_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_309),
.B1(n_333),
.B2(n_308),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_332),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_308),
.A2(n_317),
.B1(n_335),
.B2(n_296),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_238),
.A2(n_152),
.B1(n_187),
.B2(n_207),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_203),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_316),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_223),
.B(n_207),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_210),
.A2(n_206),
.B1(n_274),
.B2(n_257),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_214),
.A2(n_263),
.B1(n_217),
.B2(n_278),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g319 ( 
.A1(n_237),
.A2(n_227),
.B1(n_241),
.B2(n_236),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_319),
.B(n_334),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_296),
.B(n_313),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_250),
.A2(n_216),
.B1(n_258),
.B2(n_240),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_254),
.A2(n_274),
.B(n_275),
.C(n_277),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_264),
.A2(n_273),
.B1(n_262),
.B2(n_251),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_241),
.B(n_254),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_334),
.B(n_289),
.Y(n_359)
);

AO22x1_ASAP7_75t_SL g336 ( 
.A1(n_212),
.A2(n_220),
.B1(n_218),
.B2(n_239),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_336),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_277),
.Y(n_338)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_339),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_343),
.B(n_376),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_296),
.A2(n_234),
.B1(n_235),
.B2(n_269),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

OAI32xp33_ASAP7_75t_L g346 ( 
.A1(n_292),
.A2(n_225),
.A3(n_256),
.B1(n_245),
.B2(n_255),
.Y(n_346)
);

AOI32xp33_ASAP7_75t_L g418 ( 
.A1(n_346),
.A2(n_369),
.A3(n_373),
.B1(n_343),
.B2(n_379),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_299),
.A2(n_249),
.B1(n_260),
.B2(n_280),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_363),
.B1(n_365),
.B2(n_370),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_285),
.B(n_272),
.C(n_233),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_358),
.C(n_380),
.Y(n_388)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_353),
.Y(n_395)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_296),
.A2(n_232),
.B1(n_246),
.B2(n_298),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_355),
.A2(n_377),
.B(n_379),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_301),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_300),
.B(n_318),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_285),
.B(n_322),
.C(n_289),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_359),
.B(n_340),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_302),
.A2(n_335),
.B1(n_320),
.B2(n_299),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_360),
.A2(n_364),
.B1(n_382),
.B2(n_369),
.Y(n_421)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_361),
.B(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_366),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_285),
.A2(n_293),
.B1(n_292),
.B2(n_312),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_293),
.A2(n_326),
.B1(n_319),
.B2(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_294),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_295),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_371),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_374),
.C(n_286),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_307),
.A2(n_319),
.B1(n_298),
.B2(n_336),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_295),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_372),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_305),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_385),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_323),
.A2(n_314),
.B1(n_307),
.B2(n_306),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_378),
.B(n_383),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_316),
.A2(n_307),
.B1(n_336),
.B2(n_323),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_329),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_314),
.A2(n_311),
.B1(n_325),
.B2(n_304),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_310),
.B1(n_287),
.B2(n_297),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_325),
.A2(n_306),
.B1(n_337),
.B2(n_304),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_371),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_328),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_283),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_396),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_399),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_286),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_414),
.C(n_417),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_283),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_401),
.B(n_409),
.Y(n_456)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_382),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_411),
.Y(n_450)
);

AO21x1_ASAP7_75t_L g428 ( 
.A1(n_406),
.A2(n_418),
.B(n_353),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_380),
.B(n_287),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_408),
.B(n_401),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_342),
.B(n_330),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_416),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_381),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_340),
.B(n_310),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_413),
.A2(n_361),
.B(n_352),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_358),
.B(n_297),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_342),
.A2(n_310),
.B1(n_315),
.B2(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_415),
.A2(n_350),
.B1(n_351),
.B2(n_366),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_341),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_315),
.C(n_374),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_353),
.B(n_349),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_414),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_421),
.A2(n_352),
.B1(n_368),
.B2(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_425),
.A2(n_427),
.B(n_442),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_393),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_426),
.B(n_441),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_406),
.A2(n_420),
.B(n_417),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_428),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_398),
.A2(n_360),
.B1(n_415),
.B2(n_418),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_430),
.A2(n_432),
.B1(n_436),
.B2(n_437),
.Y(n_475)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_431),
.Y(n_466)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

XOR2x1_ASAP7_75t_SL g434 ( 
.A(n_410),
.B(n_368),
.Y(n_434)
);

XNOR2x2_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_395),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_352),
.B1(n_368),
.B2(n_344),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_411),
.A2(n_344),
.B1(n_355),
.B2(n_348),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_438),
.A2(n_403),
.B1(n_387),
.B2(n_407),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_346),
.B(n_383),
.Y(n_440)
);

AO22x2_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_395),
.B1(n_410),
.B2(n_389),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_362),
.B1(n_376),
.B2(n_378),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_399),
.A2(n_354),
.B1(n_384),
.B2(n_416),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_409),
.A2(n_404),
.B1(n_400),
.B2(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_444),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_396),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_386),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_445),
.B(n_446),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g446 ( 
.A(n_397),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_447),
.B(n_405),
.Y(n_471)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_452),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_399),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_399),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_402),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_454),
.B(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_388),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_388),
.C(n_454),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_459),
.B(n_465),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_470),
.C(n_473),
.Y(n_496)
);

O2A1O1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_462),
.A2(n_483),
.B(n_450),
.C(n_448),
.Y(n_509)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_457),
.B(n_419),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_469),
.Y(n_506)
);

MAJx2_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_395),
.C(n_408),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_392),
.C(n_398),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_448),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_472),
.A2(n_442),
.B1(n_440),
.B2(n_437),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_429),
.B(n_389),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_413),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_476),
.B(n_482),
.C(n_484),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_436),
.B(n_422),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_489),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_403),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_407),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_427),
.B(n_397),
.C(n_452),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_487),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_424),
.B(n_431),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_426),
.B(n_444),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_488),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_428),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_486),
.A2(n_425),
.B(n_453),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_490),
.A2(n_509),
.B(n_511),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_492),
.A2(n_516),
.B1(n_518),
.B2(n_462),
.Y(n_541)
);

INVx13_ASAP7_75t_L g493 ( 
.A(n_478),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_493),
.Y(n_524)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_481),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_503),
.Y(n_521)
);

INVx13_ASAP7_75t_L g497 ( 
.A(n_479),
.Y(n_497)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_497),
.Y(n_530)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_463),
.A2(n_428),
.B1(n_432),
.B2(n_423),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_500),
.Y(n_534)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_477),
.Y(n_502)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_502),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_464),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_515),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_474),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_510),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_485),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_468),
.A2(n_435),
.B(n_450),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_512),
.A2(n_435),
.B(n_456),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_472),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_513),
.B(n_514),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_475),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_484),
.B(n_456),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_460),
.B(n_447),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_519),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_520),
.B(n_541),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_461),
.C(n_465),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_526),
.B(n_529),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_496),
.B(n_470),
.C(n_459),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_469),
.C(n_480),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_531),
.B(n_538),
.C(n_542),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_510),
.A2(n_462),
.B1(n_423),
.B2(n_468),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_535),
.A2(n_508),
.B1(n_516),
.B2(n_501),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_517),
.B(n_476),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_536),
.B(n_537),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_506),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_505),
.B(n_489),
.C(n_467),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_505),
.B(n_449),
.C(n_455),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_462),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_507),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_438),
.C(n_441),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_518),
.C(n_512),
.Y(n_559)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_521),
.Y(n_545)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_545),
.Y(n_565)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_521),
.Y(n_546)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_546),
.Y(n_576)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_533),
.Y(n_547)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_547),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_491),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_549),
.A2(n_556),
.B(n_562),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_539),
.A2(n_510),
.B1(n_503),
.B2(n_491),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_551),
.A2(n_554),
.B1(n_557),
.B2(n_564),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_552),
.B(n_535),
.Y(n_574)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_527),
.B(n_495),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_540),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_522),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_558),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_559),
.B(n_561),
.Y(n_578)
);

XNOR2x1_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_536),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_528),
.B(n_498),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_494),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_500),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_563),
.B(n_523),
.Y(n_570)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_534),
.Y(n_564)
);

FAx1_ASAP7_75t_SL g567 ( 
.A(n_559),
.B(n_531),
.CI(n_523),
.CON(n_567),
.SN(n_567)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_581),
.Y(n_585)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_570),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_529),
.C(n_526),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_571),
.B(n_577),
.Y(n_593)
);

MAJx2_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_538),
.C(n_507),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_574),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_579),
.C(n_580),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_550),
.B(n_560),
.C(n_548),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_548),
.B(n_541),
.C(n_539),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_555),
.B(n_543),
.C(n_537),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_525),
.C(n_515),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_525),
.C(n_520),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_582),
.B(n_508),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_579),
.A2(n_545),
.B1(n_549),
.B2(n_508),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_592),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_573),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_584),
.A2(n_595),
.B1(n_596),
.B2(n_587),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_581),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_586),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_588),
.Y(n_600)
);

NOR2xp67_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_502),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_591),
.A2(n_564),
.B(n_530),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_578),
.B(n_524),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_556),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_582),
.Y(n_602)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_568),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_585),
.A2(n_569),
.B(n_576),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_597),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_593),
.B(n_572),
.C(n_574),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_602),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_586),
.A2(n_565),
.B(n_567),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_603),
.B(n_604),
.Y(n_613)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_589),
.B(n_580),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_575),
.C(n_554),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_605),
.B(n_606),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_607),
.B(n_530),
.Y(n_610)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_610),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_590),
.C(n_589),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_611),
.B(n_614),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_604),
.B(n_583),
.C(n_501),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_601),
.B(n_584),
.Y(n_615)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_615),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_598),
.C(n_613),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_618),
.B(n_620),
.Y(n_621)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_609),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_618),
.A2(n_612),
.B(n_598),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_622),
.B(n_616),
.C(n_617),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_623),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_624),
.A2(n_621),
.B(n_612),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_625),
.B(n_619),
.C(n_490),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_626),
.B(n_493),
.C(n_497),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_627),
.B(n_509),
.Y(n_628)
);


endmodule