module real_aes_1952_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_1066;
wire n_684;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_503;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_577;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1053;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_1025;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_725;
wire n_960;
wire n_504;
wire n_455;
wire n_671;
wire n_973;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_936;
wire n_581;
wire n_610;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_449;
wire n_1006;
wire n_607;
wire n_417;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_1031;
wire n_432;
wire n_880;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_756;
wire n_598;
wire n_404;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_727;
wire n_1014;
wire n_1056;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_765;
wire n_498;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_703;
wire n_652;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_0), .A2(n_334), .B1(n_516), .B2(n_518), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_1), .A2(n_209), .B1(n_539), .B2(n_540), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_2), .A2(n_11), .B1(n_815), .B2(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_3), .A2(n_114), .B1(n_467), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_4), .A2(n_96), .B1(n_539), .B2(n_540), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_5), .A2(n_241), .B1(n_815), .B2(n_963), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_6), .A2(n_319), .B1(n_489), .B2(n_492), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_7), .A2(n_277), .B1(n_736), .B2(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_8), .A2(n_88), .B1(n_462), .B2(n_627), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_9), .A2(n_166), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_10), .A2(n_337), .B1(n_675), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_12), .A2(n_122), .B1(n_596), .B2(n_635), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_13), .Y(n_588) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_14), .A2(n_163), .B1(n_191), .B2(n_420), .C1(n_444), .C2(n_598), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_15), .A2(n_379), .B1(n_936), .B2(n_937), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_16), .A2(n_175), .B1(n_462), .B2(n_467), .Y(n_986) );
AOI222xp33_ASAP7_75t_L g988 ( .A1(n_17), .A2(n_112), .B1(n_299), .B2(n_708), .C1(n_921), .C2(n_989), .Y(n_988) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_18), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_19), .A2(n_376), .B1(n_474), .B2(n_476), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_20), .A2(n_74), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g920 ( .A1(n_21), .A2(n_361), .B1(n_385), .B2(n_450), .C1(n_596), .C2(n_921), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_22), .A2(n_29), .B1(n_595), .B2(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_23), .B(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_24), .A2(n_244), .B1(n_520), .B2(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_25), .A2(n_149), .B1(n_490), .B2(n_787), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_26), .A2(n_243), .B1(n_543), .B2(n_573), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_27), .A2(n_245), .B1(n_677), .B2(n_946), .Y(n_945) );
INVx1_ASAP7_75t_SL g427 ( .A(n_28), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_28), .B(n_38), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_30), .A2(n_56), .B1(n_552), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_31), .A2(n_212), .B1(n_526), .B2(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_32), .A2(n_380), .B1(n_501), .B2(n_913), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_33), .A2(n_308), .B1(n_626), .B2(n_627), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_34), .A2(n_84), .B1(n_500), .B2(n_609), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_35), .A2(n_77), .B1(n_461), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_36), .A2(n_57), .B1(n_494), .B2(n_737), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_37), .A2(n_276), .B1(n_789), .B2(n_805), .Y(n_967) );
AO22x2_ASAP7_75t_L g429 ( .A1(n_38), .A2(n_377), .B1(n_426), .B2(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_39), .B(n_533), .Y(n_847) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_40), .A2(n_100), .B1(n_120), .B2(n_596), .C1(n_634), .C2(n_635), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_41), .A2(n_265), .B1(n_494), .B2(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_42), .A2(n_297), .B1(n_596), .B2(n_635), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_43), .A2(n_217), .B1(n_478), .B2(n_512), .Y(n_828) );
OA22x2_ASAP7_75t_L g414 ( .A1(n_44), .A2(n_415), .B1(n_416), .B2(n_502), .Y(n_414) );
INVx1_ASAP7_75t_L g502 ( .A(n_44), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_45), .A2(n_382), .B1(n_462), .B2(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_46), .A2(n_116), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_47), .A2(n_372), .B1(n_476), .B2(n_606), .Y(n_811) );
INVx1_ASAP7_75t_L g428 ( .A(n_48), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_49), .A2(n_255), .B1(n_501), .B2(n_902), .Y(n_940) );
AO22x1_ASAP7_75t_L g613 ( .A1(n_50), .A2(n_160), .B1(n_614), .B2(n_615), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_51), .A2(n_240), .B1(n_510), .B2(n_512), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_52), .A2(n_260), .B1(n_560), .B2(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_53), .B(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_54), .A2(n_104), .B1(n_542), .B2(n_543), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_55), .A2(n_127), .B1(n_675), .B2(n_902), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_58), .A2(n_59), .B1(n_646), .B2(n_878), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_60), .A2(n_378), .B1(n_520), .B2(n_787), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_61), .A2(n_251), .B1(n_485), .B2(n_672), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_62), .B(n_642), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_63), .A2(n_399), .B1(n_408), .B2(n_1025), .C(n_1026), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_64), .A2(n_140), .B1(n_611), .B2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_65), .A2(n_395), .B1(n_629), .B2(n_1004), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_66), .A2(n_159), .B1(n_529), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_67), .A2(n_271), .B1(n_439), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_68), .A2(n_115), .B1(n_482), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_69), .A2(n_174), .B1(n_667), .B2(n_807), .Y(n_1061) );
AO22x2_ASAP7_75t_L g436 ( .A1(n_70), .A2(n_187), .B1(n_426), .B2(n_437), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_71), .A2(n_390), .B1(n_494), .B2(n_699), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_72), .A2(n_273), .B1(n_439), .B2(n_444), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_73), .A2(n_318), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_75), .A2(n_373), .B1(n_737), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_76), .A2(n_269), .B1(n_492), .B2(n_520), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_78), .A2(n_248), .B1(n_527), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_79), .A2(n_349), .B1(n_476), .B2(n_609), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_80), .A2(n_753), .B(n_1031), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_81), .A2(n_173), .B1(n_554), .B2(n_555), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_82), .B(n_420), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_83), .A2(n_124), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_85), .A2(n_261), .B1(n_557), .B2(n_558), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_86), .A2(n_301), .B1(n_473), .B2(n_476), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_87), .A2(n_295), .B1(n_462), .B2(n_524), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_89), .A2(n_274), .B1(n_626), .B2(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_90), .A2(n_151), .B1(n_627), .B2(n_691), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_91), .A2(n_304), .B1(n_670), .B2(n_673), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_92), .A2(n_208), .B1(n_449), .B2(n_454), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_93), .A2(n_306), .B1(n_529), .B2(n_753), .Y(n_973) );
XOR2x2_ASAP7_75t_L g780 ( .A(n_94), .B(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_95), .A2(n_347), .B1(n_474), .B2(n_478), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_97), .A2(n_263), .B1(n_609), .B2(n_611), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_98), .A2(n_289), .B1(n_545), .B2(n_546), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_99), .A2(n_392), .B1(n_439), .B2(n_601), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_101), .A2(n_176), .B1(n_554), .B2(n_555), .Y(n_587) );
AOI22x1_ASAP7_75t_L g863 ( .A1(n_102), .A2(n_864), .B1(n_882), .B2(n_883), .Y(n_863) );
CKINVDCx14_ASAP7_75t_R g883 ( .A(n_102), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_103), .A2(n_203), .B1(n_450), .B2(n_596), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_105), .A2(n_330), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_106), .A2(n_126), .B1(n_529), .B2(n_596), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_107), .A2(n_224), .B1(n_485), .B2(n_614), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_108), .A2(n_130), .B1(n_462), .B2(n_524), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_109), .A2(n_210), .B1(n_482), .B2(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_110), .A2(n_358), .B1(n_607), .B2(n_853), .Y(n_852) );
AO22x2_ASAP7_75t_L g433 ( .A1(n_111), .A2(n_316), .B1(n_426), .B2(n_434), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_113), .A2(n_388), .B1(n_667), .B2(n_942), .Y(n_941) );
OA22x2_ASAP7_75t_L g976 ( .A1(n_117), .A2(n_977), .B1(n_978), .B2(n_990), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_117), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_118), .A2(n_270), .B1(n_520), .B2(n_521), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_119), .A2(n_288), .B1(n_481), .B2(n_485), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_121), .A2(n_283), .B1(n_500), .B2(n_672), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_123), .A2(n_282), .B1(n_545), .B2(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_125), .A2(n_131), .B1(n_527), .B2(n_598), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_128), .A2(n_315), .B1(n_695), .B2(n_716), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_129), .A2(n_387), .B1(n_485), .B2(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_132), .A2(n_272), .B1(n_450), .B2(n_596), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_133), .A2(n_386), .B1(n_601), .B2(n_960), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_134), .A2(n_194), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_135), .A2(n_234), .B1(n_518), .B2(n_670), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_136), .A2(n_172), .B1(n_474), .B2(n_1013), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1038 ( .A1(n_137), .A2(n_305), .B1(n_677), .B2(n_946), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_138), .A2(n_216), .B1(n_539), .B2(n_540), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_139), .A2(n_257), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_141), .A2(n_294), .B1(n_678), .B2(n_853), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_142), .A2(n_335), .B1(n_489), .B2(n_944), .Y(n_1039) );
BUFx2_ASAP7_75t_R g680 ( .A(n_143), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_144), .A2(n_314), .B1(n_805), .B2(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_145), .A2(n_259), .B1(n_596), .B2(n_635), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_146), .A2(n_302), .B1(n_807), .B2(n_808), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_147), .A2(n_352), .B1(n_551), .B2(n_552), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_148), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_150), .A2(n_351), .B1(n_808), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_152), .A2(n_285), .B1(n_560), .B2(n_673), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_153), .A2(n_211), .B1(n_807), .B2(n_969), .Y(n_968) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_154), .A2(n_252), .B1(n_665), .B2(n_667), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_155), .A2(n_222), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_156), .A2(n_357), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_157), .A2(n_250), .B1(n_494), .B2(n_520), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_158), .A2(n_375), .B1(n_543), .B2(n_573), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_161), .A2(n_307), .B1(n_598), .B2(n_897), .Y(n_896) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_162), .A2(n_267), .B1(n_659), .B2(n_663), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_164), .A2(n_221), .B1(n_545), .B2(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_165), .B(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_167), .A2(n_170), .B1(n_467), .B2(n_626), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_168), .A2(n_199), .B1(n_475), .B2(n_510), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_169), .B(n_753), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_171), .A2(n_345), .B1(n_482), .B2(n_611), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_177), .A2(n_327), .B1(n_672), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_178), .A2(n_179), .B1(n_738), .B2(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g751 ( .A(n_180), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_181), .A2(n_346), .B1(n_462), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_182), .A2(n_233), .B1(n_646), .B2(n_1050), .Y(n_1049) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_183), .A2(n_354), .B1(n_542), .B2(n_543), .Y(n_779) );
OA22x2_ASAP7_75t_L g701 ( .A1(n_184), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_184), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_185), .A2(n_350), .B1(n_497), .B2(n_697), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_186), .A2(n_200), .B1(n_716), .B2(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g1023 ( .A(n_187), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_188), .A2(n_312), .B1(n_497), .B2(n_499), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_189), .A2(n_348), .B1(n_561), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_190), .A2(n_342), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g686 ( .A(n_192), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_193), .A2(n_397), .B1(n_699), .B2(n_944), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_195), .A2(n_311), .B1(n_461), .B2(n_466), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g1010 ( .A1(n_196), .A2(n_249), .B1(n_667), .B2(n_942), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_197), .A2(n_329), .B1(n_649), .B2(n_937), .Y(n_1052) );
OA22x2_ASAP7_75t_L g505 ( .A1(n_198), .A2(n_506), .B1(n_507), .B2(n_534), .Y(n_505) );
INVx1_ASAP7_75t_L g534 ( .A(n_198), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_201), .A2(n_300), .B1(n_485), .B2(n_741), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_202), .A2(n_231), .B1(n_902), .B2(n_946), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_204), .A2(n_281), .B1(n_527), .B2(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_205), .A2(n_266), .B1(n_607), .B2(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_206), .A2(n_284), .B1(n_497), .B2(n_697), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_207), .A2(n_1028), .B1(n_1029), .B2(n_1040), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_207), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_213), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_214), .A2(n_225), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_215), .A2(n_328), .B1(n_449), .B2(n_454), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_218), .A2(n_227), .B1(n_527), .B2(n_654), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_219), .B(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_220), .A2(n_303), .B1(n_482), .B2(n_510), .Y(n_509) );
AO22x2_ASAP7_75t_L g925 ( .A1(n_223), .A2(n_926), .B1(n_927), .B2(n_947), .Y(n_925) );
INVx1_ASAP7_75t_L g947 ( .A(n_223), .Y(n_947) );
INVx1_ASAP7_75t_L g591 ( .A(n_226), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_228), .A2(n_268), .B1(n_494), .B2(n_659), .Y(n_1011) );
INVx2_ASAP7_75t_L g404 ( .A(n_229), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_230), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_232), .A2(n_331), .B1(n_598), .B2(n_824), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_235), .A2(n_296), .B1(n_557), .B2(n_558), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_236), .A2(n_394), .B1(n_626), .B2(n_627), .Y(n_825) );
OA22x2_ASAP7_75t_L g729 ( .A1(n_237), .A2(n_730), .B1(n_731), .B2(n_756), .Y(n_729) );
INVx1_ASAP7_75t_L g756 ( .A(n_237), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_238), .A2(n_247), .B1(n_646), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g643 ( .A(n_239), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_242), .A2(n_383), .B1(n_450), .B2(n_596), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_246), .A2(n_356), .B1(n_444), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_253), .A2(n_256), .B1(n_510), .B2(n_716), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_254), .A2(n_369), .B1(n_474), .B2(n_510), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_258), .A2(n_309), .B1(n_596), .B2(n_635), .Y(n_793) );
XNOR2x1_ASAP7_75t_L g820 ( .A(n_262), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g1044 ( .A(n_264), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_275), .B(n_420), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_278), .A2(n_321), .B1(n_462), .B2(n_524), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_279), .A2(n_956), .B1(n_957), .B2(n_974), .Y(n_955) );
INVx1_ASAP7_75t_L g974 ( .A(n_279), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_280), .B(n_634), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_286), .A2(n_362), .B1(n_439), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_287), .A2(n_393), .B1(n_520), .B2(n_521), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_290), .A2(n_292), .B1(n_765), .B2(n_1058), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_291), .Y(n_775) );
INVx1_ASAP7_75t_L g750 ( .A(n_293), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_298), .B(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_310), .A2(n_365), .B1(n_551), .B2(n_552), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_313), .A2(n_343), .B1(n_482), .B2(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_316), .B(n_1022), .Y(n_1021) );
OA22x2_ASAP7_75t_L g892 ( .A1(n_317), .A2(n_893), .B1(n_906), .B2(n_907), .Y(n_892) );
INVx1_ASAP7_75t_L g906 ( .A(n_317), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_320), .A2(n_370), .B1(n_512), .B2(n_611), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_322), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_323), .A2(n_363), .B1(n_601), .B2(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_324), .B(n_420), .Y(n_599) );
XOR2x2_ASAP7_75t_L g619 ( .A(n_325), .B(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_326), .A2(n_368), .B1(n_675), .B2(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_332), .A2(n_355), .B1(n_598), .B2(n_746), .Y(n_792) );
INVx3_ASAP7_75t_L g426 ( .A(n_333), .Y(n_426) );
XNOR2x2_ASAP7_75t_L g535 ( .A(n_336), .B(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_338), .A2(n_360), .B1(n_551), .B2(n_552), .Y(n_586) );
INVx1_ASAP7_75t_L g755 ( .A(n_339), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_340), .A2(n_366), .B1(n_665), .B2(n_1013), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_341), .B(n_753), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_344), .A2(n_364), .B1(n_736), .B2(n_738), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_353), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_359), .B(n_642), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_367), .A2(n_396), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g838 ( .A(n_371), .Y(n_838) );
XNOR2x1_ASAP7_75t_L g801 ( .A(n_374), .B(n_802), .Y(n_801) );
AND2x4_ASAP7_75t_L g406 ( .A(n_381), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g1019 ( .A(n_381), .Y(n_1019) );
AO21x1_ASAP7_75t_L g1065 ( .A1(n_381), .A2(n_402), .B(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g407 ( .A(n_384), .Y(n_407) );
AND2x2_ASAP7_75t_R g1042 ( .A(n_384), .B(n_1019), .Y(n_1042) );
INVxp67_ASAP7_75t_L g403 ( .A(n_389), .Y(n_403) );
NAND2xp33_ASAP7_75t_SL g1007 ( .A(n_391), .B(n_1008), .Y(n_1007) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_405), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_407), .B(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1066 ( .A(n_407), .Y(n_1066) );
AOI31xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_887), .A3(n_888), .B(n_1016), .Y(n_408) );
AO21x1_ASAP7_75t_L g1025 ( .A1(n_409), .A2(n_887), .B(n_888), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_725), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_411), .B(n_726), .Y(n_887) );
XNOR2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_563), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AO22x2_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_503), .B1(n_504), .B2(n_562), .Y(n_413) );
INVx2_ASAP7_75t_L g562 ( .A(n_414), .Y(n_562) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_471), .Y(n_416) );
NAND4xp25_ASAP7_75t_SL g417 ( .A(n_418), .B(n_438), .C(n_448), .D(n_460), .Y(n_417) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx4_ASAP7_75t_SL g533 ( .A(n_421), .Y(n_533) );
INVx4_ASAP7_75t_SL g548 ( .A(n_421), .Y(n_548) );
INVx3_ASAP7_75t_L g634 ( .A(n_421), .Y(n_634) );
INVx3_ASAP7_75t_SL g642 ( .A(n_421), .Y(n_642) );
BUFx2_ASAP7_75t_L g875 ( .A(n_421), .Y(n_875) );
INVx6_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_431), .Y(n_422) );
AND2x4_ASAP7_75t_L g446 ( .A(n_423), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g468 ( .A(n_423), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g540 ( .A(n_423), .B(n_469), .Y(n_540) );
AND2x2_ASAP7_75t_L g543 ( .A(n_423), .B(n_447), .Y(n_543) );
AND2x2_ASAP7_75t_L g574 ( .A(n_423), .B(n_447), .Y(n_574) );
AND2x4_ASAP7_75t_L g578 ( .A(n_423), .B(n_431), .Y(n_578) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_429), .Y(n_423) );
INVx2_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
AND2x2_ASAP7_75t_L g452 ( .A(n_424), .B(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
OAI22x1_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_426), .Y(n_430) );
INVx2_ASAP7_75t_L g434 ( .A(n_426), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_426), .Y(n_437) );
AND2x2_ASAP7_75t_L g442 ( .A(n_429), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g453 ( .A(n_429), .Y(n_453) );
BUFx2_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
AND2x4_ASAP7_75t_L g475 ( .A(n_431), .B(n_452), .Y(n_475) );
AND2x4_ASAP7_75t_L g484 ( .A(n_431), .B(n_479), .Y(n_484) );
AND2x2_ASAP7_75t_L g498 ( .A(n_431), .B(n_442), .Y(n_498) );
AND2x6_ASAP7_75t_L g551 ( .A(n_431), .B(n_442), .Y(n_551) );
AND2x2_ASAP7_75t_L g554 ( .A(n_431), .B(n_452), .Y(n_554) );
AND2x2_ASAP7_75t_L g584 ( .A(n_431), .B(n_479), .Y(n_584) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g441 ( .A(n_433), .B(n_435), .Y(n_441) );
AND2x2_ASAP7_75t_L g458 ( .A(n_433), .B(n_436), .Y(n_458) );
INVx1_ASAP7_75t_L g465 ( .A(n_433), .Y(n_465) );
INVxp67_ASAP7_75t_L g447 ( .A(n_435), .Y(n_447) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g464 ( .A(n_436), .B(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g526 ( .A(n_440), .Y(n_526) );
BUFx3_ASAP7_75t_L g598 ( .A(n_440), .Y(n_598) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_440), .Y(n_655) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x2_ASAP7_75t_L g451 ( .A(n_441), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g501 ( .A(n_441), .B(n_479), .Y(n_501) );
AND2x2_ASAP7_75t_L g542 ( .A(n_441), .B(n_442), .Y(n_542) );
AND2x4_ASAP7_75t_L g545 ( .A(n_441), .B(n_452), .Y(n_545) );
AND2x2_ASAP7_75t_L g561 ( .A(n_441), .B(n_479), .Y(n_561) );
AND2x2_ASAP7_75t_L g573 ( .A(n_441), .B(n_442), .Y(n_573) );
AND2x2_ASAP7_75t_L g491 ( .A(n_442), .B(n_464), .Y(n_491) );
AND2x2_ASAP7_75t_L g557 ( .A(n_442), .B(n_464), .Y(n_557) );
AND2x4_ASAP7_75t_L g479 ( .A(n_443), .B(n_453), .Y(n_479) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g527 ( .A(n_445), .Y(n_527) );
INVx2_ASAP7_75t_L g629 ( .A(n_445), .Y(n_629) );
INVx1_ASAP7_75t_L g746 ( .A(n_445), .Y(n_746) );
INVx2_ASAP7_75t_SL g815 ( .A(n_445), .Y(n_815) );
INVx2_ASAP7_75t_L g824 ( .A(n_445), .Y(n_824) );
INVx2_ASAP7_75t_L g897 ( .A(n_445), .Y(n_897) );
INVx6_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g749 ( .A(n_449), .Y(n_749) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
BUFx5_ASAP7_75t_L g635 ( .A(n_451), .Y(n_635) );
BUFx3_ASAP7_75t_L g878 ( .A(n_451), .Y(n_878) );
AND2x2_ASAP7_75t_L g463 ( .A(n_452), .B(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g539 ( .A(n_452), .B(n_464), .Y(n_539) );
INVx1_ASAP7_75t_L g972 ( .A(n_454), .Y(n_972) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g531 ( .A(n_456), .Y(n_531) );
INVx3_ASAP7_75t_L g646 ( .A(n_456), .Y(n_646) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx12f_ASAP7_75t_L g596 ( .A(n_457), .Y(n_596) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AND2x4_ASAP7_75t_L g478 ( .A(n_458), .B(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g494 ( .A(n_458), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_458), .B(n_459), .Y(n_546) );
AND2x4_ASAP7_75t_L g555 ( .A(n_458), .B(n_479), .Y(n_555) );
AND2x4_ASAP7_75t_L g558 ( .A(n_458), .B(n_495), .Y(n_558) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_458), .B(n_459), .Y(n_708) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_463), .Y(n_626) );
INVx3_ASAP7_75t_L g652 ( .A(n_463), .Y(n_652) );
AND2x4_ASAP7_75t_L g487 ( .A(n_464), .B(n_479), .Y(n_487) );
AND2x6_ASAP7_75t_L g552 ( .A(n_464), .B(n_479), .Y(n_552) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_465), .Y(n_470) );
BUFx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g524 ( .A(n_468), .Y(n_524) );
INVx2_ASAP7_75t_L g602 ( .A(n_468), .Y(n_602) );
BUFx4f_ASAP7_75t_L g627 ( .A(n_468), .Y(n_627) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .C(n_488), .D(n_496), .Y(n_471) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
INVx6_ASAP7_75t_L g610 ( .A(n_475), .Y(n_610) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_SL g607 ( .A(n_477), .Y(n_607) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g510 ( .A(n_478), .Y(n_510) );
BUFx2_ASAP7_75t_SL g678 ( .A(n_478), .Y(n_678) );
BUFx3_ASAP7_75t_L g871 ( .A(n_478), .Y(n_871) );
BUFx2_ASAP7_75t_SL g1056 ( .A(n_478), .Y(n_1056) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g560 ( .A(n_483), .Y(n_560) );
INVx2_ASAP7_75t_SL g606 ( .A(n_483), .Y(n_606) );
INVx3_ASAP7_75t_L g716 ( .A(n_483), .Y(n_716) );
INVx2_ASAP7_75t_L g902 ( .A(n_483), .Y(n_902) );
INVx3_ASAP7_75t_SL g913 ( .A(n_483), .Y(n_913) );
INVx8_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g518 ( .A(n_486), .Y(n_518) );
INVx2_ASAP7_75t_SL g615 ( .A(n_486), .Y(n_615) );
INVx2_ASAP7_75t_L g667 ( .A(n_486), .Y(n_667) );
INVx2_ASAP7_75t_L g697 ( .A(n_486), .Y(n_697) );
INVx1_ASAP7_75t_SL g808 ( .A(n_486), .Y(n_808) );
INVx2_ASAP7_75t_L g834 ( .A(n_486), .Y(n_834) );
INVx2_ASAP7_75t_L g969 ( .A(n_486), .Y(n_969) );
INVx8_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_491), .Y(n_520) );
INVx2_ASAP7_75t_L g662 ( .A(n_491), .Y(n_662) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g521 ( .A(n_493), .Y(n_521) );
INVx2_ASAP7_75t_L g663 ( .A(n_493), .Y(n_663) );
INVx2_ASAP7_75t_L g944 ( .A(n_493), .Y(n_944) );
INVx5_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g738 ( .A(n_494), .Y(n_738) );
BUFx2_ASAP7_75t_L g765 ( .A(n_494), .Y(n_765) );
BUFx3_ASAP7_75t_L g787 ( .A(n_494), .Y(n_787) );
BUFx3_ASAP7_75t_L g942 ( .A(n_497), .Y(n_942) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g517 ( .A(n_498), .Y(n_517) );
BUFx2_ASAP7_75t_L g672 ( .A(n_498), .Y(n_672) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g843 ( .A(n_500), .Y(n_843) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g514 ( .A(n_501), .Y(n_514) );
BUFx3_ASAP7_75t_L g611 ( .A(n_501), .Y(n_611) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_501), .Y(n_675) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
XNOR2x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_535), .Y(n_504) );
INVx1_ASAP7_75t_L g721 ( .A(n_505), .Y(n_721) );
BUFx2_ASAP7_75t_L g723 ( .A(n_505), .Y(n_723) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_522), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .C(n_515), .D(n_519), .Y(n_508) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_510), .Y(n_946) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g695 ( .A(n_514), .Y(n_695) );
INVx1_ASAP7_75t_L g789 ( .A(n_514), .Y(n_789) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g614 ( .A(n_517), .Y(n_614) );
INVx3_ASAP7_75t_L g741 ( .A(n_517), .Y(n_741) );
INVx2_ASAP7_75t_SL g807 ( .A(n_517), .Y(n_807) );
INVx2_ASAP7_75t_SL g855 ( .A(n_517), .Y(n_855) );
NAND4xp25_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .C(n_528), .D(n_532), .Y(n_522) );
BUFx6f_ASAP7_75t_SL g1008 ( .A(n_524), .Y(n_1008) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_549), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .C(n_544), .D(n_547), .Y(n_537) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_545), .Y(n_989) );
BUFx2_ASAP7_75t_L g930 ( .A(n_548), .Y(n_930) );
NAND4xp25_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .C(n_556), .D(n_559), .Y(n_549) );
INVx1_ASAP7_75t_L g768 ( .A(n_551), .Y(n_768) );
INVx2_ASAP7_75t_L g666 ( .A(n_560), .Y(n_666) );
BUFx6f_ASAP7_75t_L g853 ( .A(n_560), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_681), .B1(n_682), .B2(n_724), .Y(n_563) );
INVx1_ASAP7_75t_L g724 ( .A(n_564), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_617), .B2(n_618), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AO22x2_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_589), .B1(n_590), .B2(n_616), .Y(n_566) );
OA22x2_ASAP7_75t_L g861 ( .A1(n_567), .A2(n_616), .B1(n_862), .B2(n_863), .Y(n_861) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_588), .Y(n_568) );
XOR2x2_ASAP7_75t_L g616 ( .A(n_569), .B(n_588), .Y(n_616) );
NAND2x1_ASAP7_75t_SL g569 ( .A(n_570), .B(n_580), .Y(n_569) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_576), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx2_ASAP7_75t_SL g774 ( .A(n_578), .Y(n_774) );
BUFx2_ASAP7_75t_L g921 ( .A(n_578), .Y(n_921) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_585), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_593), .B(n_603), .Y(n_592) );
AND4x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .C(n_599), .D(n_600), .Y(n_593) );
INVx2_ASAP7_75t_L g754 ( .A(n_596), .Y(n_754) );
INVx1_ASAP7_75t_L g933 ( .A(n_598), .Y(n_933) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g938 ( .A(n_602), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_613), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .C(n_612), .Y(n_604) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g677 ( .A(n_610), .Y(n_677) );
INVx2_ASAP7_75t_L g785 ( .A(n_610), .Y(n_785) );
INVx2_ASAP7_75t_L g805 ( .A(n_610), .Y(n_805) );
INVx2_ASAP7_75t_L g1055 ( .A(n_610), .Y(n_1055) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_636), .Y(n_618) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .C(n_630), .D(n_633), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .Y(n_624) );
BUFx6f_ASAP7_75t_SL g936 ( .A(n_626), .Y(n_936) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AOI22x1_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_679), .B2(n_680), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_656), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_647), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_643), .B(n_644), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_642), .Y(n_753) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_653), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx4_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g691 ( .A(n_652), .Y(n_691) );
INVx1_ASAP7_75t_L g961 ( .A(n_652), .Y(n_961) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx4f_ASAP7_75t_SL g963 ( .A(n_655), .Y(n_963) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_655), .Y(n_1004) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_668), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_664), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_661), .Y(n_810) );
INVx1_ASAP7_75t_L g1059 ( .A(n_661), .Y(n_1059) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g699 ( .A(n_662), .Y(n_699) );
INVx1_ASAP7_75t_L g737 ( .A(n_662), .Y(n_737) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_676), .Y(n_668) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx6f_ASAP7_75t_L g1013 ( .A(n_675), .Y(n_1013) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx4_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_720), .B2(n_722), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI22x1_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_701), .B1(n_718), .B2(n_719), .Y(n_684) );
INVx1_ASAP7_75t_SL g719 ( .A(n_685), .Y(n_719) );
XNOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_693), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .C(n_692), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .C(n_698), .D(n_700), .Y(n_693) );
INVx3_ASAP7_75t_L g718 ( .A(n_701), .Y(n_718) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_705), .B(n_711), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .C(n_709), .D(n_710), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .C(n_717), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
XNOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_797), .Y(n_726) );
AOI22x1_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_757), .B2(n_758), .Y(n_727) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_743), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_739), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
OAI222xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_752), .C1(n_754), .C2(n_755), .Y(n_748) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OA22x2_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_780), .B1(n_795), .B2(n_796), .Y(n_758) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_759), .Y(n_796) );
XNOR2x1_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2x1p5_ASAP7_75t_L g761 ( .A(n_762), .B(n_772), .Y(n_761) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_769), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
NOR2x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_777), .Y(n_772) );
OAI21xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_775), .B(n_776), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g795 ( .A(n_780), .Y(n_795) );
NOR2xp67_ASAP7_75t_L g781 ( .A(n_782), .B(n_790), .Y(n_781) );
NAND4xp25_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .C(n_786), .D(n_788), .Y(n_782) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .C(n_793), .D(n_794), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_859), .B2(n_886), .Y(n_797) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B1(n_818), .B2(n_819), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OR2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_812), .Y(n_802) );
NAND4xp25_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .C(n_809), .D(n_811), .Y(n_803) );
NAND4xp25_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .C(n_816), .D(n_817), .Y(n_812) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_836), .B1(n_857), .B2(n_858), .Y(n_819) );
INVx2_ASAP7_75t_L g858 ( .A(n_820), .Y(n_858) );
INVx1_ASAP7_75t_L g860 ( .A(n_820), .Y(n_860) );
NAND4xp75_ASAP7_75t_L g821 ( .A(n_822), .B(n_826), .C(n_829), .D(n_832), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
AND2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g857 ( .A(n_836), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_845), .B2(n_856), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_840), .B(n_846), .C(n_851), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_844), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OR2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_851), .Y(n_845) );
NAND4xp25_ASAP7_75t_SL g846 ( .A(n_847), .B(n_848), .C(n_849), .D(n_850), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_854), .Y(n_851) );
INVx2_ASAP7_75t_L g886 ( .A(n_859), .Y(n_886) );
AO22x2_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B1(n_884), .B2(n_885), .Y(n_859) );
INVx1_ASAP7_75t_L g884 ( .A(n_860), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_861), .Y(n_885) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g882 ( .A(n_864), .Y(n_882) );
AND2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_873), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_869), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_872), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_879), .Y(n_873) );
OAI21xp5_ASAP7_75t_SL g874 ( .A1(n_875), .A2(n_876), .B(n_877), .Y(n_874) );
BUFx6f_ASAP7_75t_SL g1006 ( .A(n_878), .Y(n_1006) );
INVx1_ASAP7_75t_L g1051 ( .A(n_878), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_950), .B1(n_951), .B2(n_1015), .Y(n_888) );
INVx1_ASAP7_75t_L g1015 ( .A(n_889), .Y(n_1015) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
AOI22x1_ASAP7_75t_SL g890 ( .A1(n_891), .A2(n_925), .B1(n_948), .B2(n_949), .Y(n_890) );
INVx1_ASAP7_75t_L g949 ( .A(n_891), .Y(n_949) );
AO22x1_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_908), .B1(n_923), .B2(n_924), .Y(n_891) );
INVx1_ASAP7_75t_L g923 ( .A(n_892), .Y(n_923) );
INVx1_ASAP7_75t_L g907 ( .A(n_893), .Y(n_907) );
NOR2x1_ASAP7_75t_L g893 ( .A(n_894), .B(n_900), .Y(n_893) );
NAND4xp25_ASAP7_75t_L g894 ( .A(n_895), .B(n_896), .C(n_898), .D(n_899), .Y(n_894) );
NAND4xp25_ASAP7_75t_L g900 ( .A(n_901), .B(n_903), .C(n_904), .D(n_905), .Y(n_900) );
INVx1_ASAP7_75t_SL g924 ( .A(n_908), .Y(n_924) );
XOR2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_922), .Y(n_908) );
NAND4xp75_ASAP7_75t_L g909 ( .A(n_910), .B(n_914), .C(n_917), .D(n_920), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
AND2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
INVx4_ASAP7_75t_L g948 ( .A(n_925), .Y(n_948) );
INVx2_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
OR2x2_ASAP7_75t_L g927 ( .A(n_928), .B(n_939), .Y(n_927) );
NAND4xp25_ASAP7_75t_SL g928 ( .A(n_929), .B(n_931), .C(n_934), .D(n_935), .Y(n_928) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx3_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NAND4xp25_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .C(n_943), .D(n_945), .Y(n_939) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B1(n_992), .B2(n_995), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
AO22x1_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_975), .B2(n_991), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
NOR3xp33_ASAP7_75t_SL g957 ( .A(n_958), .B(n_964), .C(n_970), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_962), .Y(n_958) );
BUFx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVxp33_ASAP7_75t_L g1001 ( .A(n_961), .Y(n_1001) );
NAND4xp25_ASAP7_75t_SL g964 ( .A(n_965), .B(n_966), .C(n_967), .D(n_968), .Y(n_964) );
OAI21xp5_ASAP7_75t_SL g970 ( .A1(n_971), .A2(n_972), .B(n_973), .Y(n_970) );
BUFx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVxp67_ASAP7_75t_L g991 ( .A(n_976), .Y(n_991) );
INVx2_ASAP7_75t_L g990 ( .A(n_978), .Y(n_990) );
NAND4xp75_ASAP7_75t_L g978 ( .A(n_979), .B(n_982), .C(n_985), .D(n_988), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_980), .B(n_981), .Y(n_979) );
AND2x2_ASAP7_75t_L g982 ( .A(n_983), .B(n_984), .Y(n_982) );
AND2x2_ASAP7_75t_L g985 ( .A(n_986), .B(n_987), .Y(n_985) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
XNOR2x1_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
OR2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1009), .Y(n_997) );
NAND4xp25_ASAP7_75t_L g998 ( .A(n_999), .B(n_1003), .C(n_1005), .D(n_1007), .Y(n_998) );
OA21x2_ASAP7_75t_SL g999 ( .A1(n_1000), .A2(n_1001), .B(n_1002), .Y(n_999) );
NAND4xp25_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .C(n_1012), .D(n_1014), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_1017), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1020), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1018), .B(n_1021), .Y(n_1064) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
OAI222xp33_ASAP7_75t_R g1026 ( .A1(n_1027), .A2(n_1041), .B1(n_1043), .B2(n_1044), .C1(n_1062), .C2(n_1065), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_1029), .Y(n_1028) );
AND5x1_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1034), .C(n_1035), .D(n_1038), .E(n_1039), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
INVx1_ASAP7_75t_SL g1041 ( .A(n_1042), .Y(n_1041) );
XNOR2x2_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
NOR2x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1053), .Y(n_1045) );
NAND4xp25_ASAP7_75t_SL g1046 ( .A(n_1047), .B(n_1048), .C(n_1049), .D(n_1052), .Y(n_1046) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
NAND4xp25_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1057), .C(n_1060), .D(n_1061), .Y(n_1053) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_SL g1062 ( .A(n_1063), .Y(n_1062) );
CKINVDCx6p67_ASAP7_75t_R g1063 ( .A(n_1064), .Y(n_1063) );
endmodule