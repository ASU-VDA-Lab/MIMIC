module real_jpeg_14029_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_205, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_205;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_5),
.A2(n_35),
.B1(n_62),
.B2(n_64),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_5),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_5),
.B(n_57),
.C(n_59),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_5),
.A2(n_7),
.B(n_56),
.C(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_89),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_24),
.C(n_40),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_75),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_73),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_46),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_10),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_27),
.B1(n_44),
.B2(n_45),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_119),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_118),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_16),
.B(n_99),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_79),
.C(n_86),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_51),
.B2(n_52),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_53),
.C(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_21),
.A2(n_36),
.B1(n_37),
.B2(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_21),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_28),
.B(n_30),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_22),
.A2(n_28),
.B1(n_32),
.B2(n_82),
.Y(n_81)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_23),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_23),
.B(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_28),
.A2(n_30),
.B(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_28),
.B(n_35),
.Y(n_161)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_29),
.B(n_31),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_34),
.B(n_113),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_35),
.A2(n_45),
.B(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_35),
.B(n_38),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_36),
.A2(n_37),
.B1(n_146),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_36),
.A2(n_37),
.B1(n_107),
.B2(n_109),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_37),
.B(n_109),
.C(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_37),
.B(n_146),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_47),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_38),
.A2(n_47),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_38),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_50),
.Y(n_49)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_84)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_44),
.B(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_48),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_49),
.Y(n_185)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_53),
.A2(n_54),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_53),
.B(n_107),
.C(n_184),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OA21x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_65),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_73),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_67),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_76),
.B(n_77),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_76),
.B1(n_77),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_98),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_79),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_84),
.A2(n_85),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_84),
.A2(n_85),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_84),
.B(n_94),
.C(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_84),
.B(n_130),
.C(n_141),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_86),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.C(n_96),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_87),
.A2(n_96),
.B1(n_97),
.B2(n_110),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_90),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_152),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_94),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_94),
.B(n_163),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_97),
.B1(n_132),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_97),
.B(n_133),
.C(n_136),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_107),
.A2(n_109),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI321xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_188),
.A3(n_198),
.B1(n_201),
.B2(n_202),
.C(n_205),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_174),
.B(n_187),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_142),
.B(n_173),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_123),
.B(n_129),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_124),
.A2(n_125),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_167),
.B(n_172),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_154),
.B(n_166),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B(n_165),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B(n_164),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_175),
.B(n_176),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_194),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_192),
.CI(n_194),
.CON(n_200),
.SN(n_200)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_200),
.Y(n_203)
);


endmodule