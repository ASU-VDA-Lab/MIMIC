module fake_jpeg_2235_n_486 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_486);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_486;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_46),
.Y(n_116)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_51),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_69),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_68),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g121 ( 
.A(n_67),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_33),
.B(n_8),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_79),
.Y(n_123)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_42),
.B(n_18),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_92),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_38),
.Y(n_127)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_49),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_41),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_41),
.B1(n_15),
.B2(n_36),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_145),
.B1(n_50),
.B2(n_92),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_54),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_107),
.B(n_113),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_60),
.B(n_23),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_115),
.A2(n_152),
.B1(n_83),
.B2(n_64),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_128),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_34),
.C(n_15),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_24),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_146),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_47),
.A2(n_30),
.B1(n_31),
.B2(n_24),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_66),
.B(n_31),
.C(n_22),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_43),
.B(n_18),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_49),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_67),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_61),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_155),
.B(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_150),
.B1(n_149),
.B2(n_129),
.Y(n_203)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_48),
.B1(n_88),
.B2(n_87),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_160),
.A2(n_166),
.B1(n_150),
.B2(n_129),
.Y(n_208)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_0),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_188),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_103),
.A2(n_130),
.B1(n_139),
.B2(n_153),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_85),
.B(n_91),
.C(n_30),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_108),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_175),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_176),
.Y(n_217)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_72),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_178),
.Y(n_214)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_180),
.Y(n_219)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_73),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_192),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_120),
.B1(n_135),
.B2(n_143),
.Y(n_209)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_30),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_195),
.Y(n_213)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_0),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_191),
.Y(n_222)
);

CKINVDCx11_ASAP7_75t_R g191 ( 
.A(n_116),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_64),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_90),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_194),
.Y(n_229)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_141),
.B(n_81),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_80),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_143),
.Y(n_221)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_152),
.B1(n_115),
.B2(n_149),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_225),
.B1(n_155),
.B2(n_195),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_208),
.B1(n_186),
.B2(n_166),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_131),
.B(n_135),
.C(n_101),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_157),
.B(n_177),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_228),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_158),
.A2(n_96),
.B1(n_124),
.B2(n_45),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_96),
.B1(n_124),
.B2(n_59),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_191),
.B1(n_111),
.B2(n_134),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_167),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_157),
.B(n_131),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_161),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_234),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_164),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_155),
.B(n_186),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_213),
.B1(n_203),
.B2(n_227),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_157),
.C(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_222),
.C(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_199),
.B(n_183),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_223),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_243),
.Y(n_260)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

BUFx24_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_161),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_251),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_253),
.B1(n_202),
.B2(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_165),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_213),
.B(n_206),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_210),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_255),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_188),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_226),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_211),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_228),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_172),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_219),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_259),
.B(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_206),
.B(n_216),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_247),
.B(n_237),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_275),
.B1(n_276),
.B2(n_244),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_273),
.C(n_272),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_277),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_212),
.Y(n_273)
);

OAI22x1_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_244),
.B1(n_226),
.B2(n_232),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_242),
.B1(n_249),
.B2(n_247),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_208),
.B1(n_203),
.B2(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_212),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_234),
.B(n_222),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_281),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_267),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_287),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_238),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_284),
.B(n_265),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_283),
.B1(n_265),
.B2(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_291),
.B1(n_307),
.B2(n_275),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_233),
.B1(n_246),
.B2(n_232),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_252),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_294),
.C(n_302),
.Y(n_333)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_252),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_261),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_303),
.Y(n_324)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_239),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_196),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_246),
.B1(n_248),
.B2(n_252),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_252),
.C(n_245),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_302),
.C(n_287),
.Y(n_334)
);

HAxp5_ASAP7_75t_SL g309 ( 
.A(n_270),
.B(n_214),
.CON(n_309),
.SN(n_309)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_259),
.B(n_214),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_278),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_312),
.A2(n_315),
.B1(n_250),
.B2(n_254),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_270),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_190),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_316),
.B(n_319),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_290),
.A2(n_276),
.B1(n_274),
.B2(n_284),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_323),
.B1(n_289),
.B2(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_272),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_321),
.A2(n_263),
.B(n_241),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_291),
.B1(n_288),
.B2(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_280),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_326),
.B(n_328),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_224),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_310),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_299),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_293),
.B(n_271),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_331),
.B(n_219),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_336),
.C(n_338),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_292),
.B(n_265),
.C(n_271),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_294),
.B(n_266),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_295),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_235),
.C(n_221),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_349),
.B1(n_352),
.B2(n_356),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_345),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_286),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_286),
.B(n_309),
.C(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_335),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_298),
.B1(n_250),
.B2(n_257),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_329),
.Y(n_350)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_243),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_361),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_324),
.A2(n_209),
.B1(n_254),
.B2(n_263),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_353),
.A2(n_322),
.B1(n_320),
.B2(n_329),
.Y(n_375)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_335),
.B1(n_322),
.B2(n_318),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_357),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_201),
.C(n_215),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_333),
.C(n_337),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_314),
.B(n_241),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_364),
.C(n_338),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_334),
.B(n_156),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_360),
.B(n_175),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_333),
.B(n_210),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_362),
.A2(n_363),
.B(n_330),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g363 ( 
.A1(n_336),
.A2(n_263),
.B(n_205),
.C(n_220),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_365),
.A2(n_383),
.B(n_363),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_347),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_367),
.B(n_379),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_368),
.B(n_364),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_380),
.Y(n_407)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_320),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_374),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_356),
.B1(n_349),
.B2(n_341),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_327),
.C(n_201),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_327),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_263),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_204),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_348),
.A2(n_218),
.B(n_215),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_179),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_215),
.C(n_218),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_388),
.C(n_362),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_218),
.C(n_168),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_231),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_368),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_169),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_391),
.A2(n_198),
.B1(n_180),
.B2(n_51),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_398),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_385),
.A2(n_339),
.B1(n_344),
.B2(n_363),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_393),
.A2(n_400),
.B1(n_403),
.B2(n_408),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_386),
.C(n_369),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_395),
.B(n_397),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_363),
.C(n_353),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_365),
.A2(n_231),
.B(n_204),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_399),
.A2(n_371),
.B(n_366),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_382),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_406),
.Y(n_415)
);

AO221x1_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_205),
.B1(n_185),
.B2(n_189),
.C(n_187),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_402),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_194),
.C(n_178),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_389),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_372),
.A2(n_205),
.B1(n_134),
.B2(n_162),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_370),
.A2(n_75),
.B1(n_56),
.B2(n_53),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_410),
.A2(n_366),
.B1(n_387),
.B2(n_383),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_378),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_416),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_377),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_421),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_375),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_424),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_423),
.A2(n_405),
.B1(n_394),
.B2(n_400),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_374),
.C(n_376),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_426),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_159),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_171),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_427),
.B(n_428),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_409),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_429),
.A2(n_399),
.B1(n_390),
.B2(n_404),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_413),
.A2(n_405),
.B(n_398),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_430),
.A2(n_438),
.B1(n_442),
.B2(n_415),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_397),
.B(n_403),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_432),
.A2(n_414),
.B(n_425),
.Y(n_448)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_434),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_173),
.C(n_143),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_436),
.B(n_412),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_424),
.A2(n_173),
.B(n_106),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_420),
.B(n_109),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_439),
.B(n_8),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_109),
.B1(n_105),
.B2(n_98),
.Y(n_441)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_441),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_421),
.A2(n_109),
.B1(n_105),
.B2(n_98),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_449),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_431),
.A2(n_430),
.B(n_440),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_447),
.A2(n_448),
.B(n_450),
.Y(n_462)
);

O2A1O1Ixp5_ASAP7_75t_L g450 ( 
.A1(n_433),
.A2(n_429),
.B(n_30),
.C(n_2),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_432),
.A2(n_105),
.B1(n_106),
.B2(n_32),
.Y(n_451)
);

AOI211xp5_ASAP7_75t_L g461 ( 
.A1(n_451),
.A2(n_442),
.B(n_32),
.C(n_5),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_1),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_9),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_2),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_437),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_455),
.B(n_444),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_32),
.C(n_0),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_436),
.C(n_438),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_458),
.B(n_10),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_467),
.C(n_466),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_463),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_461),
.Y(n_469)
);

AOI322xp5_ASAP7_75t_L g464 ( 
.A1(n_446),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_464),
.A2(n_456),
.B1(n_465),
.B2(n_467),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_3),
.B(n_6),
.C(n_9),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_465),
.A2(n_462),
.B(n_454),
.Y(n_468)
);

INVx11_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_470),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_471),
.A2(n_472),
.B(n_463),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_460),
.A2(n_457),
.B(n_11),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_11),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_477),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_476),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_473),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_12),
.Y(n_479)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_479),
.B(n_12),
.CI(n_13),
.CON(n_481),
.SN(n_481)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_481),
.A2(n_478),
.B(n_13),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_480),
.B(n_482),
.Y(n_484)
);

AOI31xp33_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_13),
.A3(n_14),
.B(n_477),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_13),
.Y(n_486)
);


endmodule