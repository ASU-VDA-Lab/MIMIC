module real_jpeg_15740_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_SL g89 ( 
.A(n_0),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_2),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_4),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_4),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_5),
.B(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_7),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_7),
.B(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_18),
.Y(n_17)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_10),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_10),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_79),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_95),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_64),
.B(n_94),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_49),
.B(n_63),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_26),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_16),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_22),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_21),
.B(n_88),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_40),
.C(n_44),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_62),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_66),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_82),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_84),
.C(n_85),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_80),
.C(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_80),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_127),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_99),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

XNOR2x1_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);


endmodule