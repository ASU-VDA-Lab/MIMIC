module fake_jpeg_23892_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_26),
.A2(n_28),
.B1(n_14),
.B2(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_31),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_18),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_42),
.B(n_44),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_28),
.B1(n_15),
.B2(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_18),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_15),
.Y(n_44)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_50),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_30),
.B(n_29),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_59),
.B(n_21),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_29),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_7),
.B(n_8),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_26),
.B1(n_44),
.B2(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_34),
.Y(n_63)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_30),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_70),
.C(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_34),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_58),
.C(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_46),
.B1(n_58),
.B2(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_80),
.B1(n_65),
.B2(n_53),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_81),
.C(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_70),
.B(n_49),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_86),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_59),
.C(n_61),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_74),
.B1(n_83),
.B2(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_83),
.B1(n_76),
.B2(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_100),
.B1(n_12),
.B2(n_23),
.Y(n_103)
);

AOI21x1_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_53),
.B(n_21),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_12),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_61),
.B(n_38),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_100),
.C(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_102),
.A3(n_17),
.B1(n_23),
.B2(n_11),
.C1(n_7),
.C2(n_2),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_106),
.C(n_1),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_108),
.C(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_2),
.Y(n_111)
);


endmodule