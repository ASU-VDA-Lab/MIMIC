module fake_jpeg_24925_n_160 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_160);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_26),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_23),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_17),
.B1(n_22),
.B2(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_25),
.B1(n_13),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_17),
.B1(n_22),
.B2(n_15),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_21),
.B1(n_19),
.B2(n_29),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_29),
.B(n_28),
.C(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_61),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_45),
.B(n_23),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_56),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_76),
.B1(n_37),
.B2(n_40),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_52),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_45),
.C(n_44),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_37),
.B1(n_40),
.B2(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_84),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_64),
.C(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_28),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_90),
.B(n_75),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_94),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_88),
.B(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_97),
.B1(n_98),
.B2(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_68),
.B1(n_72),
.B2(n_63),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_101),
.C(n_104),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_65),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_67),
.C(n_28),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_84),
.B1(n_78),
.B2(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_112),
.B1(n_20),
.B2(n_91),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_78),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_115),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_77),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_110),
.C(n_33),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_101),
.B1(n_96),
.B2(n_102),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_82),
.B1(n_67),
.B2(n_14),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_57),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_42),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_119),
.C(n_125),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_123),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_42),
.B1(n_33),
.B2(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_33),
.C(n_31),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_106),
.C(n_113),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_108),
.C(n_107),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_20),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B1(n_118),
.B2(n_120),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_31),
.B1(n_42),
.B2(n_65),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_122),
.C(n_2),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_139),
.C(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_122),
.C(n_2),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_1),
.C(n_3),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_1),
.C(n_4),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_6),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_5),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_8),
.Y(n_152)
);

AOI31xp33_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_145),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_5),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_7),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_148),
.B(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_151),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_8),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_147),
.B(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_9),
.C(n_10),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_156),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_157),
.B(n_153),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_10),
.Y(n_160)
);


endmodule