module fake_jpeg_29257_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_7),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_13),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_22),
.B(n_6),
.Y(n_25)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_9),
.Y(n_20)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_10),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_10),
.B1(n_7),
.B2(n_6),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_28),
.B1(n_15),
.B2(n_20),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_27),
.B(n_24),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_34),
.C(n_25),
.Y(n_37)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_28),
.C(n_23),
.Y(n_38)
);


endmodule