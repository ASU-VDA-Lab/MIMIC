module fake_jpeg_19610_n_42 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_42);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_42;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_19),
.B1(n_22),
.B2(n_21),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_22),
.B1(n_18),
.B2(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_11),
.C(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_1),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_31),
.B(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_25),
.B1(n_26),
.B2(n_6),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_25),
.C(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_36),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_4),
.B(n_7),
.Y(n_41)
);

AOI221xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_4),
.B1(n_9),
.B2(n_13),
.C(n_15),
.Y(n_42)
);


endmodule