module real_jpeg_15489_n_25 (n_17, n_8, n_0, n_157, n_21, n_168, n_2, n_10, n_9, n_12, n_156, n_24, n_165, n_166, n_6, n_159, n_161, n_162, n_169, n_167, n_23, n_11, n_14, n_160, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_25);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_168;
input n_2;
input n_10;
input n_9;
input n_12;
input n_156;
input n_24;
input n_165;
input n_166;
input n_6;
input n_159;
input n_161;
input n_162;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_160;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_1),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_4),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_4),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_5),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_5),
.B(n_68),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_7),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.C(n_120),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_11),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_11),
.B(n_96),
.C(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_12),
.B(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

AOI322xp5_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_74),
.A3(n_86),
.B1(n_89),
.B2(n_127),
.C1(n_129),
.C2(n_167),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_15),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_45),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_17),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_21),
.B(n_64),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g93 ( 
.A1(n_22),
.A2(n_94),
.B(n_106),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_24),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_24),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_30),
.B(n_152),
.Y(n_151)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_31),
.B(n_90),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_149),
.B(n_154),
.Y(n_35)
);

OAI31xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_60),
.A3(n_132),
.B(n_135),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.C(n_55),
.Y(n_37)
);

AOI321xp33_ASAP7_75t_L g135 ( 
.A1(n_38),
.A2(n_48),
.A3(n_136),
.B1(n_137),
.B2(n_140),
.C(n_168),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_44),
.Y(n_38)
);

OAI322xp33_ASAP7_75t_L g140 ( 
.A1(n_39),
.A2(n_49),
.A3(n_141),
.B1(n_146),
.B2(n_147),
.C1(n_148),
.C2(n_169),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_44),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_55),
.B(n_142),
.C(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_56),
.B(n_59),
.Y(n_136)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI31xp67_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.A3(n_91),
.B(n_123),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_73),
.C(n_79),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_81),
.C(n_128),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_79),
.A3(n_124),
.B1(n_125),
.B2(n_126),
.C(n_166),
.Y(n_123)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_113),
.C(n_114),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.C(n_102),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_153),
.Y(n_154)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_156),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_157),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_158),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_159),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_160),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_161),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_162),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_163),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_164),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_165),
.Y(n_121)
);


endmodule