module fake_jpeg_6258_n_77 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_0),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_57),
.B1(n_41),
.B2(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_61),
.B1(n_42),
.B2(n_38),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_50),
.B1(n_46),
.B2(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_58),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.C(n_68),
.Y(n_69)
);

A2O1A1O1Ixp25_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_10),
.B(n_12),
.C(n_15),
.D(n_18),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_19),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_21),
.B(n_23),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_24),
.C(n_25),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_26),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_29),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_30),
.B(n_31),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_35),
.Y(n_77)
);


endmodule