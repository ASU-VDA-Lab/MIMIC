module fake_jpeg_18801_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_24),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_13),
.Y(n_49)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_34),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_19),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_12),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_48),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_27),
.B1(n_25),
.B2(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_55),
.B1(n_62),
.B2(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_30),
.B1(n_17),
.B2(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_7),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_30),
.B(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_47),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_30),
.B1(n_11),
.B2(n_13),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_11),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_35),
.B1(n_41),
.B2(n_30),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_56),
.B1(n_54),
.B2(n_53),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_35),
.B1(n_47),
.B2(n_10),
.Y(n_74)
);

OAI22x1_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_52),
.B1(n_55),
.B2(n_62),
.Y(n_81)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_65),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_70),
.C(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_58),
.B(n_50),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_82),
.B1(n_67),
.B2(n_57),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_80),
.B(n_79),
.C(n_75),
.D(n_76),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.C(n_81),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_76),
.C(n_75),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_85),
.C(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.C(n_94),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_61),
.C(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_93),
.B1(n_63),
.B2(n_9),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_8),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_99),
.C(n_63),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_101),
.Y(n_104)
);


endmodule