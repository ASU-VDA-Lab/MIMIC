module fake_jpeg_2666_n_532 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_532);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_514;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

AND2x4_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_18),
.Y(n_59)
);

OR2x4_ASAP7_75t_L g137 ( 
.A(n_59),
.B(n_35),
.Y(n_137)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_97),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_67),
.B(n_81),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_29),
.A2(n_52),
.B1(n_44),
.B2(n_27),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_35),
.B1(n_48),
.B2(n_33),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_22),
.B(n_8),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_90),
.A2(n_99),
.B(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_47),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_102),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_100),
.Y(n_145)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_31),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_31),
.B1(n_30),
.B2(n_46),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_106),
.A2(n_119),
.B1(n_135),
.B2(n_140),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_50),
.B(n_49),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_113),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_69),
.A2(n_31),
.B1(n_28),
.B2(n_33),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_84),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_50),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_150),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_79),
.A2(n_98),
.B1(n_96),
.B2(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_137),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_48),
.B1(n_45),
.B2(n_36),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_54),
.A2(n_46),
.B(n_43),
.C(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_54),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_76),
.B(n_37),
.C(n_43),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_31),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_49),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_56),
.A2(n_19),
.B1(n_42),
.B2(n_21),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_39),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_72),
.A2(n_45),
.B1(n_36),
.B2(n_37),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_74),
.A2(n_19),
.B1(n_42),
.B2(n_21),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_87),
.B(n_39),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_116),
.Y(n_203)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_165),
.B(n_166),
.Y(n_240)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_167),
.Y(n_249)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_169),
.Y(n_242)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_171),
.B(n_172),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_137),
.B1(n_88),
.B2(n_80),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_175),
.A2(n_193),
.B1(n_198),
.B2(n_204),
.Y(n_257)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_101),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_199),
.Y(n_245)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_75),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_187),
.Y(n_230)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_90),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_129),
.A2(n_95),
.B1(n_115),
.B2(n_94),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_197),
.B1(n_213),
.B2(n_215),
.Y(n_224)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_63),
.B1(n_61),
.B2(n_70),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_148),
.B1(n_106),
.B2(n_116),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_194),
.A2(n_6),
.B1(n_16),
.B2(n_13),
.Y(n_263)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_124),
.A2(n_103),
.B1(n_99),
.B2(n_93),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_31),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_201),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_126),
.B(n_10),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_203),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_127),
.A2(n_47),
.B1(n_41),
.B2(n_26),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_207),
.Y(n_260)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_120),
.B(n_9),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_7),
.C(n_16),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_119),
.B1(n_124),
.B2(n_147),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_238),
.B1(n_239),
.B2(n_214),
.Y(n_277)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_173),
.A2(n_136),
.A3(n_111),
.B1(n_117),
.B2(n_108),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_169),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_197),
.B1(n_173),
.B2(n_165),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_237),
.B1(n_248),
.B2(n_191),
.Y(n_267)
);

AO22x1_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_109),
.B1(n_107),
.B2(n_147),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_234),
.A2(n_4),
.B(n_5),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_161),
.B1(n_149),
.B2(n_142),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_181),
.A2(n_161),
.B1(n_149),
.B2(n_141),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_47),
.B(n_41),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_183),
.B(n_208),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_187),
.A2(n_41),
.B1(n_9),
.B2(n_10),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_10),
.Y(n_286)
);

MAJx3_ASAP7_75t_L g261 ( 
.A(n_163),
.B(n_176),
.C(n_180),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_261),
.B(n_0),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_11),
.B(n_17),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_162),
.C(n_167),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_294),
.C(n_299),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_275),
.B1(n_282),
.B2(n_300),
.Y(n_313)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_270),
.A2(n_249),
.B1(n_250),
.B2(n_254),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_255),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_283),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_277),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_164),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_278),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_195),
.B1(n_184),
.B2(n_190),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_245),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_170),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_284),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_280),
.A2(n_281),
.B(n_296),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_219),
.A2(n_178),
.B1(n_182),
.B2(n_196),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_240),
.A2(n_192),
.B1(n_186),
.B2(n_199),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_240),
.B(n_212),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_209),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_288),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_0),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_243),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_6),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_297),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_261),
.B(n_213),
.Y(n_291)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_292),
.B(n_295),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_258),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_1),
.C(n_2),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_234),
.A2(n_11),
.B1(n_16),
.B2(n_3),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_222),
.B(n_1),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_257),
.A2(n_11),
.B1(n_16),
.B2(n_3),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_248),
.B1(n_262),
.B2(n_233),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_1),
.C(n_2),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_237),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_3),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_308),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_302),
.A2(n_225),
.B(n_252),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_4),
.Y(n_303)
);

OAI211xp5_ASAP7_75t_SL g341 ( 
.A1(n_303),
.A2(n_305),
.B(n_308),
.C(n_285),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_224),
.A2(n_5),
.B(n_11),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_304),
.A2(n_302),
.B(n_294),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_12),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_243),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_307),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_243),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_260),
.B(n_12),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_260),
.B(n_12),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_252),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_312),
.A2(n_324),
.B1(n_313),
.B2(n_322),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_314),
.B(n_325),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_316),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_323),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_305),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_267),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_335),
.B1(n_342),
.B2(n_348),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_218),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_347),
.C(n_266),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_272),
.A2(n_218),
.B1(n_226),
.B2(n_253),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_269),
.B1(n_276),
.B2(n_292),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_225),
.B(n_226),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_309),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_333),
.B(n_344),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_277),
.B1(n_275),
.B2(n_299),
.Y(n_335)
);

AO22x1_ASAP7_75t_L g336 ( 
.A1(n_291),
.A2(n_233),
.B1(n_235),
.B2(n_262),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_336),
.A2(n_294),
.B(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_246),
.B1(n_253),
.B2(n_221),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_345),
.A2(n_346),
.B(n_283),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_288),
.A2(n_284),
.B(n_279),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_266),
.B(n_235),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_282),
.A2(n_246),
.B1(n_250),
.B2(n_249),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_314),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_356),
.A2(n_358),
.B1(n_362),
.B2(n_371),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_291),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_363),
.C(n_378),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_331),
.A2(n_271),
.B1(n_291),
.B2(n_304),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_330),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_376),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_360),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_301),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_373),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_293),
.B1(n_300),
.B2(n_287),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_293),
.C(n_301),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_315),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_317),
.Y(n_370)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_316),
.A2(n_306),
.B1(n_289),
.B2(n_307),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_310),
.B(n_290),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_335),
.A2(n_298),
.B1(n_296),
.B2(n_281),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_325),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_268),
.B1(n_286),
.B2(n_274),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_384),
.B1(n_342),
.B2(n_332),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_333),
.B(n_232),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_377),
.B(n_379),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_310),
.B(n_264),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_228),
.C(n_254),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_381),
.C(n_326),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_228),
.C(n_264),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_345),
.Y(n_408)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_373),
.B(n_319),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_406),
.C(n_372),
.Y(n_417)
);

AO22x2_ASAP7_75t_L g388 ( 
.A1(n_354),
.A2(n_328),
.B1(n_339),
.B2(n_336),
.Y(n_388)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_366),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_397),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_367),
.A2(n_336),
.B(n_311),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_415),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_352),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_337),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_405),
.C(n_389),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_384),
.A2(n_313),
.B1(n_323),
.B2(n_340),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_402),
.A2(n_404),
.B1(n_414),
.B2(n_374),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_353),
.B(n_351),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_412),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_413),
.B1(n_358),
.B2(n_367),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_368),
.Y(n_410)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_410),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_411),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_380),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_364),
.A2(n_340),
.B1(n_321),
.B2(n_338),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_362),
.A2(n_338),
.B1(n_346),
.B2(n_337),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_375),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_431),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_378),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_398),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_419),
.A2(n_438),
.B1(n_388),
.B2(n_392),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_387),
.A2(n_382),
.B1(n_360),
.B2(n_368),
.Y(n_420)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

OAI21xp33_ASAP7_75t_L g421 ( 
.A1(n_387),
.A2(n_360),
.B(n_354),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_421),
.B(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_424),
.A2(n_407),
.B1(n_395),
.B2(n_392),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_425),
.A2(n_436),
.B1(n_393),
.B2(n_400),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_433),
.C(n_434),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_399),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_410),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_403),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_439),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_357),
.C(n_363),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_389),
.B(n_361),
.C(n_318),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_391),
.A2(n_312),
.B1(n_370),
.B2(n_369),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_398),
.B(n_318),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_433),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_397),
.A2(n_350),
.B1(n_383),
.B2(n_311),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_441),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_385),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_442),
.B(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_446),
.A2(n_448),
.B1(n_464),
.B2(n_438),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_425),
.A2(n_409),
.B1(n_396),
.B2(n_402),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_411),
.B(n_385),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_460),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_401),
.C(n_435),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_455),
.C(n_458),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_456),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_408),
.C(n_414),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_407),
.C(n_395),
.Y(n_458)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_424),
.B(n_426),
.CI(n_388),
.CON(n_460),
.SN(n_460)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_462),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_416),
.A2(n_388),
.B1(n_350),
.B2(n_341),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_344),
.C(n_388),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_453),
.C(n_458),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_416),
.A2(n_348),
.B1(n_327),
.B2(n_274),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_443),
.B(n_432),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_470),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_457),
.A2(n_422),
.B(n_426),
.Y(n_469)
);

NOR3xp33_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_476),
.C(n_439),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_429),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_447),
.Y(n_484)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_451),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_472),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_429),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_475),
.B(n_481),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_445),
.A2(n_422),
.B(n_423),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_437),
.C(n_440),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_447),
.C(n_445),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_484),
.Y(n_503)
);

AOI221xp5_ASAP7_75t_L g485 ( 
.A1(n_477),
.A2(n_446),
.B1(n_461),
.B2(n_460),
.C(n_454),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_488),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_456),
.C(n_455),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_479),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_474),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_442),
.B1(n_464),
.B2(n_459),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_495),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_463),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_494),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_436),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_492),
.A2(n_476),
.B(n_469),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_462),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_467),
.B(n_327),
.C(n_460),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_468),
.A2(n_251),
.B1(n_270),
.B2(n_264),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_496),
.A2(n_480),
.B(n_474),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_264),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_465),
.Y(n_510)
);

NOR2x1_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_477),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_500),
.A2(n_508),
.B(n_486),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_504),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_510),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_478),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_506),
.B(n_507),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_487),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_493),
.A2(n_465),
.B(n_270),
.Y(n_508)
);

OAI21x1_ASAP7_75t_SL g522 ( 
.A1(n_511),
.A2(n_513),
.B(n_515),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_488),
.C(n_497),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_498),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_509),
.A2(n_485),
.B1(n_251),
.B2(n_242),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_518),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_505),
.A2(n_227),
.B(n_232),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_521),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_500),
.C(n_499),
.Y(n_521)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_516),
.A2(n_509),
.B(n_510),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_516),
.B(n_511),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_526),
.B(n_242),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_520),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_520),
.Y(n_527)
);

OAI21x1_ASAP7_75t_SL g529 ( 
.A1(n_527),
.A2(n_528),
.B(n_227),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g530 ( 
.A(n_529),
.Y(n_530)
);

OAI321xp33_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_13),
.A3(n_17),
.B1(n_229),
.B2(n_241),
.C(n_526),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_229),
.C(n_241),
.Y(n_532)
);


endmodule