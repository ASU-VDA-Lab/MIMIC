module fake_jpeg_2062_n_96 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_24),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_30),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_33),
.B1(n_27),
.B2(n_32),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_39),
.B1(n_36),
.B2(n_40),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_30),
.C(n_27),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_29),
.A3(n_34),
.B1(n_26),
.B2(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_25),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_40),
.B(n_39),
.C(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_56),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_34),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_15),
.B(n_23),
.C(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_26),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_50),
.B1(n_6),
.B2(n_7),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_64),
.B1(n_62),
.B2(n_66),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_77),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_50),
.B(n_6),
.C(n_7),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_5),
.B(n_8),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_75),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_8),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_14),
.C(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_83),
.B1(n_85),
.B2(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_84),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_87),
.C(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_81),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_78),
.B(n_80),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_75),
.Y(n_96)
);


endmodule