module fake_jpeg_23913_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_17),
.Y(n_48)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_23),
.B1(n_29),
.B2(n_32),
.Y(n_57)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_55),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_23),
.B1(n_16),
.B2(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_40),
.B1(n_37),
.B2(n_54),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_18),
.B(n_26),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_19),
.B1(n_26),
.B2(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_19),
.B1(n_39),
.B2(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_17),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_41),
.B1(n_36),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_68),
.B1(n_59),
.B2(n_50),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_73),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_41),
.B1(n_36),
.B2(n_40),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_42),
.B(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_37),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_42),
.B(n_49),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_59),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_74),
.B1(n_82),
.B2(n_79),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_35),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_102),
.C(n_107),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_101),
.B(n_110),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_35),
.B(n_54),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_67),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_112),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_40),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_40),
.C(n_62),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_76),
.C(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_24),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_27),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_78),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_64),
.B1(n_72),
.B2(n_84),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_127),
.B1(n_131),
.B2(n_111),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_137),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_72),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_129),
.C(n_100),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_81),
.B(n_87),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_132),
.B(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_74),
.B1(n_82),
.B2(n_50),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_138),
.B1(n_21),
.B2(n_20),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_37),
.B1(n_49),
.B2(n_73),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_62),
.B(n_37),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_62),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_98),
.B(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_24),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_108),
.B1(n_106),
.B2(n_102),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_113),
.B(n_96),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_111),
.B(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_90),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_38),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_92),
.Y(n_164)
);

XOR2x2_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_17),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_147),
.C(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_157),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_34),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_158),
.B1(n_159),
.B2(n_168),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_34),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_143),
.B(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_47),
.B1(n_100),
.B2(n_69),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_124),
.B1(n_131),
.B2(n_129),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_103),
.CI(n_69),
.CON(n_160),
.SN(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_47),
.B1(n_86),
.B2(n_95),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_172),
.B1(n_142),
.B2(n_21),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_133),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_103),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_103),
.B1(n_27),
.B2(n_21),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_92),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_86),
.B1(n_28),
.B2(n_25),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_141),
.B1(n_119),
.B2(n_136),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_28),
.C(n_25),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_130),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_187),
.Y(n_200)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_139),
.B1(n_132),
.B2(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_176),
.A2(n_182),
.B1(n_183),
.B2(n_197),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_132),
.B(n_123),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_196),
.C(n_147),
.Y(n_203)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_174),
.B1(n_192),
.B2(n_193),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_118),
.B1(n_120),
.B2(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_140),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_193),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_163),
.B1(n_156),
.B2(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_119),
.B(n_122),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_192),
.B(n_152),
.Y(n_217)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_177),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_217),
.B(n_202),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_145),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_213),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_206),
.B1(n_218),
.B2(n_192),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_205),
.C(n_207),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_150),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_208),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_153),
.C(n_148),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_167),
.C(n_159),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_160),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_160),
.C(n_149),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_212),
.C(n_20),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_158),
.C(n_156),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_151),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_184),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_178),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_230),
.B1(n_198),
.B2(n_217),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_190),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_188),
.B1(n_186),
.B2(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_183),
.B(n_178),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_184),
.B1(n_182),
.B2(n_197),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_173),
.B(n_180),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_1),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_187),
.B(n_1),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_28),
.C(n_25),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_0),
.B(n_1),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_203),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_205),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_204),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_200),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_3),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_247),
.C(n_232),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_22),
.C(n_2),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_220),
.B1(n_225),
.B2(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_239),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_226),
.B(n_229),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.C(n_247),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_231),
.C(n_224),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_222),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_257),
.B(n_259),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_241),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_236),
.B(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_9),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_239),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_254),
.B(n_250),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_252),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_9),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_265),
.B1(n_9),
.B2(n_5),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_15),
.B1(n_8),
.B2(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_250),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_8),
.A3(n_13),
.B1(n_5),
.B2(n_6),
.C1(n_15),
.C2(n_10),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_268),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_275),
.A2(n_267),
.B(n_269),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_277),
.A3(n_278),
.B1(n_279),
.B2(n_272),
.C1(n_10),
.C2(n_6),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.C(n_12),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_270),
.A3(n_272),
.B1(n_6),
.B2(n_8),
.C1(n_10),
.C2(n_12),
.Y(n_281)
);

AOI321xp33_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_3),
.A3(n_4),
.B1(n_12),
.B2(n_13),
.C(n_227),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_13),
.Y(n_284)
);


endmodule