module fake_jpeg_1850_n_316 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_51),
.B(n_53),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_1),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_57),
.Y(n_111)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_59),
.Y(n_118)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_19),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_73),
.Y(n_110)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_68),
.B(n_80),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_35),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_89),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_20),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_102),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_45),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_99),
.Y(n_137)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_30),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_17),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_17),
.B1(n_48),
.B2(n_46),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_49),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_32),
.B1(n_48),
.B2(n_46),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_121),
.B1(n_128),
.B2(n_142),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_32),
.B1(n_23),
.B2(n_42),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_145),
.B1(n_86),
.B2(n_100),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_23),
.B1(n_44),
.B2(n_42),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_24),
.B1(n_44),
.B2(n_30),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_93),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_51),
.B(n_50),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_53),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_103),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_88),
.B1(n_64),
.B2(n_84),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_24),
.B1(n_5),
.B2(n_8),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_151),
.B1(n_139),
.B2(n_108),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_3),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_11),
.B1(n_3),
.B2(n_10),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_95),
.B1(n_87),
.B2(n_80),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_85),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_156),
.A2(n_161),
.B1(n_153),
.B2(n_119),
.Y(n_206)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_158),
.Y(n_197)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_179),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_70),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_163),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_82),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_164),
.B(n_166),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_99),
.B1(n_72),
.B2(n_97),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_195),
.B(n_127),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_110),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_121),
.B(n_106),
.C(n_123),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_183),
.B(n_184),
.C(n_153),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_122),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_91),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_170),
.B(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_135),
.A2(n_105),
.B(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_163),
.C(n_162),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_114),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_104),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_107),
.C(n_109),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_152),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_152),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_185),
.Y(n_216)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_128),
.B(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_125),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_124),
.B(n_125),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_191),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_129),
.B(n_151),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_190),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_148),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_122),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_158),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_147),
.Y(n_195)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_208),
.B1(n_179),
.B2(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_217),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_113),
.B1(n_119),
.B2(n_162),
.Y(n_208)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_186),
.A3(n_173),
.B1(n_168),
.B2(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_221),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_215),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_183),
.B1(n_180),
.B2(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_238),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_180),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_244),
.C(n_223),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_241),
.B1(n_246),
.B2(n_244),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_195),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_240),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_180),
.B1(n_184),
.B2(n_167),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_195),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_180),
.B1(n_184),
.B2(n_190),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_157),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_249),
.Y(n_265)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_215),
.B1(n_207),
.B2(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_192),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_188),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_204),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_210),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_218),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_252),
.C(n_259),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_219),
.C(n_199),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_230),
.B(n_241),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_236),
.B(n_243),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_223),
.B1(n_226),
.B2(n_222),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_197),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_211),
.C(n_198),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_247),
.C(n_235),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_248),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_235),
.C(n_239),
.Y(n_267)
);

OAI322xp33_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_271),
.A3(n_265),
.B1(n_264),
.B2(n_257),
.C1(n_262),
.C2(n_252),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_249),
.B(n_228),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_255),
.B1(n_260),
.B2(n_224),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_198),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_251),
.C(n_259),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_238),
.B(n_236),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_275),
.B(n_276),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_197),
.B(n_224),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_255),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_289),
.Y(n_295)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_263),
.C(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_269),
.C(n_278),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_279),
.B1(n_273),
.B2(n_276),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_282),
.B1(n_287),
.B2(n_284),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_279),
.C(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_291),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_285),
.B1(n_284),
.B2(n_275),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_292),
.C(n_289),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_301),
.B(n_294),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_309),
.B(n_222),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_300),
.B1(n_298),
.B2(n_295),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_310),
.B(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_210),
.B(n_196),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_196),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_314),
.Y(n_316)
);


endmodule