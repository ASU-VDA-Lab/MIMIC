module fake_netlist_6_3023_n_1898 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1898);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1898;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_3),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_67),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_54),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_89),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_6),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_118),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_3),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_80),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_37),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_27),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_86),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_25),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_99),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_63),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_69),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_45),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_51),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_117),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_147),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_5),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_54),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_19),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_171),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_76),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_109),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_22),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_37),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_72),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_77),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_161),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_70),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_11),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_44),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_130),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_60),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_39),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_14),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_119),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_18),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_88),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_5),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_51),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_18),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_46),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_94),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_116),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_33),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_61),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_133),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_12),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_114),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_46),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_159),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_87),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_138),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_13),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_91),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_8),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_124),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_8),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_15),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_39),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_156),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_110),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_149),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_170),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_126),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_115),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_68),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_79),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_28),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_71),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_11),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_127),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_17),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_162),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_184),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_58),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_6),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_1),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_25),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_167),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_38),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_135),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_43),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_75),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_36),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_35),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_21),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_29),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_16),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_65),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_90),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_84),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_15),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_181),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_38),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_13),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_139),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_120),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_145),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_112),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_125),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_41),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_140),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_152),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_108),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_175),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_41),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_9),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_123),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_95),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_148),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_57),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_48),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_73),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_30),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_19),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_141),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_23),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_177),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_32),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_59),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_57),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_146),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_85),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_62),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_74),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_0),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_83),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_144),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_43),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_53),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_165),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_180),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_17),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_122),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_100),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_134),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_50),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_45),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_81),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_187),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_240),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_221),
.B(n_0),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_218),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_257),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_223),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_226),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_186),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_186),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_256),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_186),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_227),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_267),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_250),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_234),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_235),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_186),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_186),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_277),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_284),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_221),
.B(n_2),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_236),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_R g392 ( 
.A(n_189),
.B(n_289),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_277),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_238),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_245),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_277),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_193),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_247),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_261),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_290),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_277),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_262),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_307),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_221),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_303),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_303),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_240),
.B(n_4),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_271),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_303),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_336),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_273),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_303),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_209),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_250),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_241),
.B(n_4),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_272),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_272),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_275),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_303),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_343),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_193),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_196),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_195),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_196),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_278),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_213),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_188),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_283),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_219),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_285),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_220),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_266),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_286),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_222),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_291),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_189),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_292),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_294),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_229),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_309),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_296),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_298),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_299),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_204),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_231),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_360),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_300),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_189),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_316),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_232),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_239),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_317),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_242),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_198),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_323),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_324),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_315),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_325),
.Y(n_460)
);

INVx6_ASAP7_75t_L g461 ( 
.A(n_429),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_405),
.B(n_289),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_372),
.B(n_289),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_372),
.B(n_241),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_398),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_383),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_365),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_429),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_383),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_379),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_417),
.B(n_365),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_449),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_418),
.B(n_192),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_456),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_228),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_396),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_396),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_416),
.A2(n_252),
.B(n_228),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_415),
.B(n_252),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_406),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_390),
.B(n_348),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_390),
.B(n_348),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_410),
.A2(n_263),
.B(n_253),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_415),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_408),
.B(n_192),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_420),
.B(n_361),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_361),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_371),
.B(n_194),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_425),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_209),
.Y(n_528)
);

NAND2x1p5_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_258),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

BUFx12f_ASAP7_75t_L g531 ( 
.A(n_369),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_436),
.B(n_190),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_392),
.B(n_190),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_436),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_441),
.B(n_254),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_441),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_457),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_426),
.B(n_446),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_447),
.B(n_254),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_424),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_510),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_510),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_466),
.B(n_190),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_485),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_475),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_512),
.B(n_370),
.Y(n_547)
);

AND3x1_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_274),
.C(n_268),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_512),
.B(n_373),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_485),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_475),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_512),
.B(n_375),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_465),
.B(n_190),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_204),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_519),
.A2(n_428),
.B1(n_442),
.B2(n_434),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_529),
.B(n_428),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_469),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_524),
.A2(n_295),
.B1(n_287),
.B2(n_340),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_510),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_510),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_459),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_527),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_516),
.B(n_382),
.C(n_381),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_463),
.B(n_447),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_529),
.B(n_190),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_529),
.B(n_208),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_537),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_374),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_527),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_531),
.B(n_529),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_376),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_524),
.B(n_384),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_468),
.B(n_385),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_527),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_468),
.B(n_391),
.Y(n_583)
);

BUFx6f_ASAP7_75t_SL g584 ( 
.A(n_466),
.Y(n_584)
);

OAI21xp33_ASAP7_75t_SL g585 ( 
.A1(n_464),
.A2(n_304),
.B(n_293),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_524),
.A2(n_334),
.B1(n_319),
.B2(n_366),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_473),
.B(n_394),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_473),
.B(n_395),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_529),
.B(n_208),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_530),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_536),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_465),
.B(n_208),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_483),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_486),
.A2(n_448),
.B1(n_403),
.B2(n_458),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_469),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_536),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_469),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_465),
.B(n_208),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_483),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_538),
.Y(n_604)
);

BUFx4f_ASAP7_75t_L g605 ( 
.A(n_531),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_469),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_462),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_461),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_465),
.B(n_466),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_461),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_461),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_462),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_484),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_462),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_463),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_484),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_467),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_486),
.A2(n_460),
.B1(n_399),
.B2(n_454),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_468),
.B(n_400),
.Y(n_624)
);

AND3x4_ASAP7_75t_L g625 ( 
.A(n_509),
.B(n_459),
.C(n_401),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_471),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_466),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_494),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_465),
.B(n_208),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_465),
.B(n_409),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_473),
.B(n_412),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_494),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_477),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_477),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_538),
.A2(n_200),
.B1(n_311),
.B2(n_357),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_472),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_472),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_472),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

INVx6_ASAP7_75t_L g640 ( 
.A(n_474),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_509),
.B(n_482),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_500),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_516),
.B(n_419),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_494),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_476),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_478),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_500),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_495),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_466),
.B(n_427),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_533),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_478),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_477),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_470),
.B(n_430),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_533),
.A2(n_367),
.B1(n_314),
.B2(n_452),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_474),
.Y(n_658)
);

AND3x2_ASAP7_75t_L g659 ( 
.A(n_466),
.B(n_202),
.C(n_414),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_477),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_464),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_470),
.B(n_432),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_495),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_464),
.A2(n_440),
.B1(n_451),
.B2(n_445),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_506),
.B(n_435),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_477),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_500),
.Y(n_667)
);

INVxp33_ASAP7_75t_L g668 ( 
.A(n_482),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_478),
.Y(n_669)
);

AND2x2_ASAP7_75t_SL g670 ( 
.A(n_506),
.B(n_507),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_506),
.B(n_389),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_495),
.Y(n_672)
);

BUFx4f_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_495),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_463),
.B(n_437),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_480),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_480),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_497),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_480),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_477),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_506),
.B(n_439),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_489),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_487),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_506),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_497),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_489),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_528),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_533),
.A2(n_455),
.B1(n_453),
.B2(n_452),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_497),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_497),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_481),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_645),
.B(n_533),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_673),
.B(n_474),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_668),
.B(n_443),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_645),
.B(n_644),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_670),
.A2(n_404),
.B1(n_411),
.B2(n_507),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_565),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_656),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_667),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_668),
.B(n_444),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

BUFx2_ASAP7_75t_R g702 ( 
.A(n_551),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_540),
.A2(n_533),
.B1(n_507),
.B2(n_506),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_533),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_541),
.A2(n_533),
.B1(n_463),
.B2(n_492),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_673),
.B(n_474),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_662),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_546),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_546),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_662),
.B(n_533),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_541),
.B(n_492),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_542),
.A2(n_533),
.B1(n_507),
.B2(n_498),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_578),
.B(n_580),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_670),
.A2(n_533),
.B1(n_492),
.B2(n_461),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_661),
.A2(n_687),
.B1(n_610),
.B2(n_630),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_566),
.Y(n_717)
);

AND2x4_ASAP7_75t_SL g718 ( 
.A(n_577),
.B(n_315),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_588),
.B(n_492),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_571),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_652),
.B(n_474),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_570),
.B(n_518),
.C(n_493),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_652),
.B(n_474),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_649),
.B(n_518),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_652),
.B(n_490),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_544),
.B(n_507),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_571),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_576),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_684),
.B(n_490),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_544),
.B(n_507),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_590),
.B(n_518),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_684),
.B(n_490),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_597),
.B(n_487),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_631),
.B(n_490),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_582),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_581),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_684),
.B(n_490),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_587),
.B(n_490),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_589),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_584),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_592),
.Y(n_742)
);

AO22x1_ASAP7_75t_L g743 ( 
.A1(n_583),
.A2(n_205),
.B1(n_362),
.B2(n_359),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_610),
.A2(n_318),
.B1(n_341),
.B2(n_288),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_627),
.B(n_487),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_552),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_493),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_596),
.B(n_599),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_543),
.A2(n_498),
.B1(n_535),
.B2(n_539),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_567),
.Y(n_750)
);

NOR2x1p5_ASAP7_75t_L g751 ( 
.A(n_547),
.B(n_205),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_617),
.B(n_493),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_608),
.Y(n_753)
);

BUFx5_ASAP7_75t_L g754 ( 
.A(n_556),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_671),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_641),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_613),
.B(n_461),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_675),
.B(n_528),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_615),
.B(n_461),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_630),
.B(n_528),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_688),
.B(n_256),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_616),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_641),
.B(n_194),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_604),
.B(n_535),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_567),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_641),
.B(n_583),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_659),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_624),
.B(n_535),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_624),
.B(n_539),
.C(n_224),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_627),
.B(n_487),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_621),
.B(n_461),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_627),
.B(n_487),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_664),
.B(n_197),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_568),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_626),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_665),
.A2(n_335),
.B1(n_338),
.B2(n_346),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_568),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_609),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_637),
.B(n_525),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_665),
.B(n_681),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_609),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_638),
.B(n_525),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_550),
.A2(n_487),
.B(n_498),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_620),
.B(n_539),
.Y(n_785)
);

BUFx12f_ASAP7_75t_L g786 ( 
.A(n_557),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_569),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_554),
.B(n_453),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_688),
.B(n_487),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_564),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_639),
.B(n_525),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_642),
.B(n_525),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_647),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_651),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_648),
.B(n_525),
.Y(n_795)
);

OAI221xp5_ASAP7_75t_L g796 ( 
.A1(n_561),
.A2(n_414),
.B1(n_201),
.B2(n_320),
.C(n_203),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_657),
.B(n_487),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_654),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_545),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_657),
.B(n_487),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_669),
.B(n_525),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_681),
.B(n_197),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_676),
.B(n_525),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_677),
.B(n_525),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_577),
.B(n_455),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_679),
.B(n_517),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_569),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_682),
.B(n_517),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_686),
.B(n_517),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_562),
.B(n_517),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_577),
.B(n_214),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_555),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_611),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_315),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_563),
.A2(n_517),
.B1(n_251),
.B2(n_244),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_572),
.B(n_256),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_572),
.B(n_517),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_594),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_594),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_658),
.B(n_256),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_559),
.B(n_237),
.C(n_216),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_573),
.B(n_256),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_601),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_573),
.B(n_591),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_601),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_629),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_591),
.B(n_532),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_548),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_560),
.B(n_532),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_629),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_595),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_651),
.B(n_256),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_559),
.A2(n_329),
.B1(n_331),
.B2(n_206),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_558),
.B(n_522),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_564),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_595),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_SL g837 ( 
.A(n_605),
.B(n_191),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_585),
.B(n_256),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_602),
.Y(n_839)
);

INVxp33_ASAP7_75t_SL g840 ( 
.A(n_575),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_658),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_560),
.B(n_653),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_602),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_653),
.B(n_532),
.Y(n_844)
);

INVxp33_ASAP7_75t_L g845 ( 
.A(n_625),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_655),
.B(n_532),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_655),
.B(n_532),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_549),
.B(n_579),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_549),
.B(n_532),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_606),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_549),
.B(n_489),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_549),
.B(n_256),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_561),
.B(n_199),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_545),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_579),
.B(n_491),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_586),
.A2(n_199),
.B1(n_206),
.B2(n_210),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_605),
.B(n_522),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_635),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_606),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_611),
.Y(n_860)
);

O2A1O1Ixp5_ASAP7_75t_L g861 ( 
.A1(n_553),
.A2(n_511),
.B(n_479),
.C(n_488),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_764),
.B(n_574),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_860),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_713),
.B(n_586),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_835),
.B(n_522),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_698),
.B(n_625),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_703),
.A2(n_598),
.B(n_553),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_713),
.B(n_579),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_831),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_699),
.B(n_635),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_707),
.B(n_579),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_831),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_784),
.A2(n_618),
.B(n_614),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_703),
.Y(n_874)
);

AOI21xp33_ASAP7_75t_L g875 ( 
.A1(n_773),
.A2(n_635),
.B(n_246),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_752),
.A2(n_598),
.B(n_553),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_732),
.B(n_603),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_704),
.A2(n_600),
.B(n_598),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_848),
.A2(n_623),
.B(n_600),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_860),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_695),
.B(n_248),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_699),
.B(n_354),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_732),
.B(n_603),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_761),
.A2(n_526),
.B(n_534),
.C(n_356),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_782),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_720),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_782),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_711),
.B(n_768),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_727),
.A2(n_623),
.B(n_600),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_737),
.B(n_794),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_727),
.A2(n_634),
.B(n_623),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_781),
.A2(n_353),
.B(n_344),
.C(n_330),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_727),
.A2(n_680),
.B(n_634),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_711),
.B(n_603),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_799),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_710),
.A2(n_680),
.B(n_634),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_719),
.B(n_603),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_781),
.A2(n_640),
.B1(n_612),
.B2(n_217),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_782),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_724),
.B(n_612),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_728),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_838),
.A2(n_796),
.B(n_726),
.C(n_731),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_727),
.A2(n_849),
.B(n_824),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_719),
.B(n_607),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_692),
.A2(n_680),
.B(n_633),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_694),
.B(n_607),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_754),
.B(n_555),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_785),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_758),
.B(n_788),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_782),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_694),
.B(n_607),
.Y(n_911)
);

NOR2x2_ASAP7_75t_L g912 ( 
.A(n_811),
.B(n_207),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_700),
.B(n_210),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_810),
.A2(n_633),
.B(n_607),
.Y(n_914)
);

NAND2x1_ASAP7_75t_L g915 ( 
.A(n_779),
.B(n_640),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_779),
.A2(n_660),
.B(n_633),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_827),
.A2(n_660),
.B(n_633),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_817),
.A2(n_666),
.B(n_660),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_841),
.B(n_523),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_754),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_829),
.A2(n_666),
.B(n_660),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_844),
.A2(n_666),
.B(n_683),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_861),
.A2(n_618),
.B(n_614),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_712),
.A2(n_628),
.B(n_619),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_700),
.B(n_666),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_758),
.B(n_691),
.Y(n_926)
);

OAI21xp33_ASAP7_75t_L g927 ( 
.A1(n_853),
.A2(n_215),
.B(n_207),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_788),
.B(n_715),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_813),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_802),
.B(n_249),
.C(n_243),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_802),
.A2(n_363),
.B(n_368),
.C(n_327),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_712),
.A2(n_628),
.B(n_619),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_754),
.B(n_691),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_846),
.A2(n_683),
.B(n_691),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_749),
.A2(n_643),
.B(n_632),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_756),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_717),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_697),
.B(n_260),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_749),
.A2(n_643),
.B(n_632),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_847),
.A2(n_683),
.B(n_689),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_854),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_813),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_717),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_842),
.A2(n_690),
.B(n_689),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_754),
.B(n_555),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_702),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_745),
.A2(n_690),
.B(n_685),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_813),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_754),
.B(n_736),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_754),
.B(n_555),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_714),
.A2(n_685),
.B(n_678),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_813),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_740),
.B(n_555),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_742),
.B(n_646),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_766),
.B(n_858),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_751),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_729),
.Y(n_957)
);

BUFx12f_ASAP7_75t_L g958 ( 
.A(n_786),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_753),
.B(n_646),
.Y(n_959)
);

OR2x6_ASAP7_75t_SL g960 ( 
.A(n_696),
.B(n_215),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_745),
.A2(n_678),
.B(n_674),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_770),
.A2(n_674),
.B(n_672),
.Y(n_962)
);

AO21x1_ASAP7_75t_L g963 ( 
.A1(n_832),
.A2(n_270),
.B(n_326),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_793),
.B(n_650),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_828),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_705),
.A2(n_672),
.B(n_663),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_770),
.A2(n_663),
.B(n_650),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_798),
.B(n_640),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_818),
.A2(n_305),
.B(n_225),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_773),
.B(n_211),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_762),
.B(n_230),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_772),
.A2(n_534),
.B(n_526),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_775),
.B(n_233),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_772),
.A2(n_534),
.B(n_526),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_853),
.A2(n_265),
.B(n_264),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_L g976 ( 
.A(n_743),
.B(n_211),
.C(n_212),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_819),
.A2(n_259),
.B(n_255),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_760),
.B(n_837),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_701),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_760),
.A2(n_212),
.B1(n_350),
.B2(n_351),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_790),
.B(n_534),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_757),
.A2(n_501),
.B(n_502),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_857),
.B(n_350),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_776),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_812),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_776),
.B(n_491),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_759),
.A2(n_501),
.B(n_502),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_823),
.A2(n_351),
.B1(n_352),
.B2(n_355),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_814),
.B(n_352),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_834),
.B(n_347),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_838),
.A2(n_496),
.B(n_491),
.C(n_504),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_747),
.B(n_496),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_748),
.B(n_496),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_771),
.A2(n_508),
.B(n_501),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_693),
.A2(n_508),
.B(n_501),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_744),
.B(n_504),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_825),
.B(n_504),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_826),
.A2(n_505),
.B(n_513),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_830),
.A2(n_355),
.B1(n_358),
.B2(n_364),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_769),
.B(n_358),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_701),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_812),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_805),
.B(n_364),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_722),
.B(n_505),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_832),
.B(n_505),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_693),
.A2(n_508),
.B(n_502),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_L g1008 ( 
.A(n_815),
.B(n_763),
.C(n_833),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_706),
.A2(n_508),
.B(n_502),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_787),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_706),
.A2(n_515),
.B(n_479),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_805),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_836),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_767),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_763),
.B(n_269),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_806),
.A2(n_515),
.B(n_479),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_816),
.A2(n_513),
.B(n_479),
.C(n_488),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_815),
.B(n_513),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_790),
.B(n_523),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_807),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_808),
.A2(n_515),
.B(n_479),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_859),
.B(n_488),
.Y(n_1022)
);

NOR2xp67_ASAP7_75t_L g1023 ( 
.A(n_755),
.B(n_523),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_809),
.A2(n_488),
.B(n_503),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_839),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_843),
.B(n_488),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_735),
.A2(n_333),
.B1(n_279),
.B2(n_280),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_701),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_840),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_850),
.B(n_503),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_721),
.A2(n_515),
.B(n_511),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_780),
.A2(n_503),
.B(n_511),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_721),
.A2(n_511),
.B(n_503),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_845),
.B(n_777),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_734),
.B(n_520),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_723),
.A2(n_520),
.B(n_514),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_708),
.B(n_520),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_783),
.A2(n_520),
.B(n_276),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_723),
.A2(n_514),
.B(n_499),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_741),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_816),
.A2(n_332),
.B(n_521),
.C(n_499),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_725),
.A2(n_739),
.B(n_855),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_725),
.A2(n_514),
.B(n_499),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_851),
.A2(n_514),
.B(n_499),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_811),
.B(n_821),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_791),
.A2(n_514),
.B(n_499),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_718),
.B(n_347),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_709),
.B(n_521),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_718),
.B(n_349),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_920),
.A2(n_730),
.B(n_733),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_970),
.A2(n_822),
.B(n_820),
.C(n_811),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_880),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_869),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_862),
.B(n_741),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_881),
.B(n_856),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_908),
.B(n_741),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_875),
.A2(n_822),
.B(n_852),
.C(n_730),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_SL g1058 ( 
.A(n_866),
.B(n_349),
.C(n_359),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_975),
.A2(n_852),
.B(n_733),
.C(n_738),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_888),
.B(n_716),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_957),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_908),
.B(n_738),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_864),
.B(n_746),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_874),
.B(n_750),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_881),
.B(n_792),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_874),
.A2(n_1008),
.B1(n_920),
.B2(n_928),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_941),
.B(n_795),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_882),
.B(n_801),
.Y(n_1068)
);

AO22x1_ASAP7_75t_L g1069 ( 
.A1(n_990),
.A2(n_362),
.B1(n_281),
.B2(n_313),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_868),
.A2(n_909),
.B1(n_960),
.B2(n_949),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1034),
.A2(n_804),
.B1(n_803),
.B2(n_765),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_907),
.A2(n_789),
.B(n_800),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_900),
.B(n_1002),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_1002),
.B(n_980),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1015),
.A2(n_778),
.B(n_774),
.C(n_800),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_882),
.B(n_321),
.C(n_297),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_867),
.A2(n_789),
.B(n_797),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_900),
.B(n_797),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_936),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_913),
.A2(n_282),
.B(n_301),
.C(n_302),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1023),
.B(n_337),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_872),
.Y(n_1082)
);

AO21x1_ASAP7_75t_L g1083 ( 
.A1(n_906),
.A2(n_332),
.B(n_9),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_991),
.B(n_328),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_937),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_936),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_899),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_943),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_1028),
.B(n_521),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_1012),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_969),
.A2(n_342),
.B1(n_308),
.B2(n_310),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_976),
.B(n_927),
.C(n_1001),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_870),
.B(n_345),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_1040),
.B(n_306),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1012),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_958),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_965),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_978),
.A2(n_339),
.B1(n_312),
.B2(n_521),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_985),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1034),
.B(n_332),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_919),
.B(n_521),
.Y(n_1101)
);

INVx5_ASAP7_75t_L g1102 ( 
.A(n_977),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_925),
.B(n_521),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_906),
.B(n_521),
.Y(n_1104)
);

AO21x1_ASAP7_75t_L g1105 ( 
.A1(n_911),
.A2(n_332),
.B(n_10),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_1014),
.B(n_521),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_954),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_897),
.A2(n_514),
.B(n_499),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_886),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_911),
.B(n_332),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_866),
.B(n_7),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_L g1112 ( 
.A1(n_1042),
.A2(n_332),
.B(n_78),
.C(n_183),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_955),
.A2(n_514),
.B1(n_499),
.B2(n_481),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_977),
.B(n_514),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_959),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_880),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_956),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_890),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_977),
.B(n_499),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_877),
.B(n_332),
.Y(n_1120)
);

INVx6_ASAP7_75t_L g1121 ( 
.A(n_880),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_904),
.A2(n_481),
.B(n_129),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1029),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_955),
.A2(n_481),
.B1(n_10),
.B2(n_14),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_880),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_883),
.B(n_332),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_976),
.A2(n_481),
.B1(n_21),
.B2(n_22),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_993),
.B(n_994),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_979),
.A2(n_481),
.B1(n_64),
.B2(n_82),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_895),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_894),
.B(n_481),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_902),
.A2(n_481),
.B(n_23),
.C(n_24),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_871),
.B(n_926),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_938),
.B(n_7),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_878),
.A2(n_93),
.B(n_173),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_902),
.A2(n_174),
.B(n_169),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1045),
.B(n_930),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_901),
.B(n_26),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1020),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_863),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_931),
.A2(n_26),
.B(n_27),
.C(n_31),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1020),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_977),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_938),
.B(n_31),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_986),
.B(n_96),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_984),
.B(n_1004),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1010),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1047),
.B(n_32),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_863),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_1027),
.B(n_33),
.C(n_34),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_873),
.A2(n_1035),
.B(n_903),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1013),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_896),
.A2(n_97),
.B(n_164),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1045),
.B(n_166),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1025),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_892),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_899),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_899),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_964),
.Y(n_1159)
);

CKINVDCx11_ASAP7_75t_R g1160 ( 
.A(n_946),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1049),
.B(n_40),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1019),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1162)
);

INVx3_ASAP7_75t_SL g1163 ( 
.A(n_912),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_876),
.A2(n_104),
.B(n_155),
.Y(n_1164)
);

AOI22x1_ASAP7_75t_L g1165 ( 
.A1(n_1033),
.A2(n_1011),
.B1(n_947),
.B2(n_962),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_933),
.A2(n_103),
.B(n_151),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_989),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_987),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_998),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_971),
.B(n_973),
.C(n_997),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_981),
.B(n_47),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_L g1172 ( 
.A(n_986),
.B(n_102),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_865),
.B(n_107),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1018),
.B(n_50),
.C(n_52),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1000),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1005),
.A2(n_55),
.B1(n_56),
.B2(n_113),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1037),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_885),
.B(n_128),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_910),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_905),
.A2(n_137),
.B(n_158),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_910),
.Y(n_1181)
);

OR2x6_ASAP7_75t_SL g1182 ( 
.A(n_968),
.B(n_953),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1006),
.A2(n_884),
.B(n_1038),
.C(n_999),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_986),
.B(n_1003),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_885),
.B(n_887),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_945),
.A2(n_950),
.B(n_879),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_887),
.B(n_952),
.Y(n_1187)
);

INVx8_ASAP7_75t_L g1188 ( 
.A(n_986),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1022),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_910),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_923),
.A2(n_944),
.B(n_914),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_910),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_982),
.B(n_963),
.C(n_884),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1026),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1030),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_889),
.A2(n_891),
.B(n_893),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_917),
.A2(n_918),
.B(n_932),
.Y(n_1197)
);

NOR2x1_ASAP7_75t_L g1198 ( 
.A(n_942),
.B(n_952),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_924),
.A2(n_939),
.B(n_935),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_SL g1200 ( 
.A(n_982),
.B(n_898),
.C(n_1024),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_929),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_SL g1202 ( 
.A1(n_951),
.A2(n_966),
.B(n_1032),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_929),
.B(n_948),
.Y(n_1203)
);

AOI22x1_ASAP7_75t_L g1204 ( 
.A1(n_961),
.A2(n_967),
.B1(n_972),
.B2(n_974),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_929),
.A2(n_948),
.B1(n_1003),
.B2(n_942),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_929),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_948),
.B(n_921),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_948),
.B(n_1003),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1199),
.A2(n_915),
.B(n_916),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_SL g1210 ( 
.A1(n_1132),
.A2(n_1048),
.B(n_992),
.C(n_1031),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1079),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1092),
.A2(n_1021),
.B1(n_1016),
.B2(n_1009),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1134),
.A2(n_1007),
.B1(n_996),
.B2(n_940),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1196),
.A2(n_922),
.B(n_934),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1169),
.B(n_1044),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1136),
.A2(n_1105),
.B(n_1083),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_1136),
.A2(n_992),
.B(n_1036),
.C(n_1043),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1183),
.A2(n_1039),
.B(n_1046),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1197),
.A2(n_983),
.A3(n_988),
.B(n_995),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1202),
.A2(n_1017),
.B(n_1041),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1116),
.Y(n_1221)
);

AO21x1_ASAP7_75t_L g1222 ( 
.A1(n_1144),
.A2(n_1041),
.B(n_1017),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1097),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1128),
.A2(n_1050),
.B(n_1103),
.Y(n_1224)
);

NAND3x1_ASAP7_75t_L g1225 ( 
.A(n_1171),
.B(n_1111),
.C(n_1076),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1128),
.A2(n_1059),
.B(n_1104),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1077),
.A2(n_1066),
.B(n_1135),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1061),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1200),
.A2(n_1051),
.B(n_1170),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1170),
.A2(n_1186),
.B(n_1207),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1068),
.B(n_1065),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_L g1232 ( 
.A(n_1150),
.B(n_1127),
.C(n_1091),
.Y(n_1232)
);

AO32x2_ASAP7_75t_L g1233 ( 
.A1(n_1066),
.A2(n_1124),
.A3(n_1070),
.B1(n_1091),
.B2(n_1113),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1152),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1153),
.A2(n_1075),
.B(n_1072),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1090),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1148),
.A2(n_1161),
.B1(n_1078),
.B2(n_1174),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1167),
.A2(n_1115),
.B1(n_1107),
.B2(n_1168),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1110),
.A2(n_1126),
.A3(n_1120),
.B(n_1070),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1130),
.A2(n_1123),
.B1(n_1118),
.B2(n_1138),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1057),
.A2(n_1060),
.B(n_1131),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1060),
.A2(n_1131),
.B(n_1063),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1154),
.A2(n_1062),
.B(n_1173),
.C(n_1100),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1086),
.B(n_1146),
.Y(n_1244)
);

AOI221x1_ASAP7_75t_L g1245 ( 
.A1(n_1124),
.A2(n_1122),
.B1(n_1193),
.B2(n_1164),
.C(n_1180),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1151),
.A2(n_1191),
.B(n_1165),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1184),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1204),
.A2(n_1108),
.B(n_1178),
.Y(n_1248)
);

OA22x2_ASAP7_75t_L g1249 ( 
.A1(n_1095),
.A2(n_1163),
.B1(n_1093),
.B2(n_1054),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1084),
.B(n_1109),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1137),
.B(n_1081),
.Y(n_1251)
);

NAND3x1_ASAP7_75t_L g1252 ( 
.A(n_1129),
.B(n_1198),
.C(n_1160),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_SL g1253 ( 
.A(n_1102),
.B(n_1143),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1133),
.A2(n_1120),
.B(n_1126),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1117),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1098),
.A2(n_1166),
.B1(n_1133),
.B2(n_1064),
.C(n_1113),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1155),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1064),
.A2(n_1119),
.B(n_1114),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1112),
.A2(n_1071),
.B(n_1189),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1074),
.Y(n_1260)
);

BUFx4f_ASAP7_75t_SL g1261 ( 
.A(n_1056),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1114),
.A2(n_1119),
.B(n_1203),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1080),
.A2(n_1175),
.B(n_1156),
.C(n_1141),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1184),
.A2(n_1205),
.B(n_1143),
.Y(n_1264)
);

BUFx8_ASAP7_75t_L g1265 ( 
.A(n_1116),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1194),
.A2(n_1195),
.B(n_1177),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_SL g1267 ( 
.A(n_1102),
.B(n_1052),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1098),
.A2(n_1185),
.A3(n_1187),
.B(n_1159),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1172),
.A2(n_1208),
.B(n_1102),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1102),
.A2(n_1078),
.B(n_1101),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1067),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1087),
.A2(n_1157),
.B(n_1145),
.Y(n_1272)
);

AOI221x1_ASAP7_75t_L g1273 ( 
.A1(n_1087),
.A2(n_1157),
.B1(n_1181),
.B2(n_1182),
.C(n_1085),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1088),
.B(n_1099),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1073),
.A2(n_1145),
.B(n_1201),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1053),
.B(n_1082),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1162),
.A2(n_1176),
.B(n_1147),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1140),
.B(n_1149),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1106),
.A2(n_1089),
.B1(n_1142),
.B2(n_1139),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1073),
.B(n_1069),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1116),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1206),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1101),
.A2(n_1106),
.B(n_1188),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1125),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1192),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1058),
.A2(n_1188),
.B(n_1125),
.C(n_1190),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1179),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1190),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1052),
.A2(n_1121),
.B1(n_1089),
.B2(n_1094),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1089),
.A2(n_1074),
.B(n_1179),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1188),
.A2(n_1158),
.B(n_1190),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1121),
.B(n_1158),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1074),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1079),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1084),
.B(n_862),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1097),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1079),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1300)
);

NOR2xp67_ASAP7_75t_L g1301 ( 
.A(n_1123),
.B(n_737),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1055),
.A2(n_970),
.B1(n_1008),
.B2(n_1092),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1061),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1128),
.B(n_888),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1151),
.A2(n_873),
.B(n_1196),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1151),
.A2(n_873),
.B(n_1196),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1151),
.A2(n_873),
.B(n_1196),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1083),
.A2(n_1105),
.A3(n_1197),
.B(n_1066),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1079),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1055),
.B(n_698),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1136),
.A2(n_1105),
.B(n_1083),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1151),
.A2(n_873),
.B(n_1196),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1184),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1090),
.B(n_604),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1055),
.B(n_695),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1152),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1134),
.A2(n_970),
.B(n_707),
.C(n_698),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1055),
.A2(n_970),
.B(n_707),
.Y(n_1322)
);

AO32x2_ASAP7_75t_L g1323 ( 
.A1(n_1066),
.A2(n_1124),
.A3(n_1070),
.B1(n_1091),
.B2(n_1027),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1202),
.A2(n_1199),
.B(n_1136),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1097),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1090),
.B(n_604),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_SL g1327 ( 
.A(n_1055),
.B(n_970),
.C(n_537),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1116),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1202),
.A2(n_1199),
.B(n_1136),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1090),
.B(n_604),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1134),
.A2(n_970),
.B(n_707),
.C(n_698),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1061),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1128),
.B(n_888),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1079),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1055),
.A2(n_970),
.B(n_781),
.C(n_707),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1151),
.A2(n_873),
.B(n_1196),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1134),
.A2(n_970),
.B(n_707),
.C(n_698),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_1191),
.B(n_1199),
.Y(n_1339)
);

NAND2x1_ASAP7_75t_L g1340 ( 
.A(n_1184),
.B(n_1143),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1128),
.A2(n_864),
.B1(n_874),
.B2(n_698),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1055),
.A2(n_970),
.B(n_781),
.C(n_707),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1079),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1083),
.A2(n_1105),
.A3(n_1197),
.B(n_1066),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1055),
.A2(n_970),
.B1(n_881),
.B2(n_389),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1128),
.A2(n_864),
.B1(n_874),
.B2(n_698),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1136),
.A2(n_1191),
.B(n_1199),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1050),
.A2(n_1062),
.B(n_1151),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_1123),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1055),
.B(n_698),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1055),
.A2(n_970),
.B(n_781),
.C(n_707),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1199),
.A2(n_673),
.B(n_703),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1086),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1151),
.A2(n_873),
.B(n_1196),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1055),
.A2(n_970),
.B(n_781),
.C(n_707),
.Y(n_1357)
);

BUFx12f_ASAP7_75t_L g1358 ( 
.A(n_1096),
.Y(n_1358)
);

INVx6_ASAP7_75t_SL g1359 ( 
.A(n_1074),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1202),
.A2(n_1199),
.B(n_1136),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1128),
.B(n_888),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1123),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_1123),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1302),
.A2(n_1232),
.B1(n_1345),
.B2(n_1327),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1358),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1247),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1225),
.A2(n_1312),
.B1(n_1322),
.B2(n_1232),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1362),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1231),
.B(n_1305),
.Y(n_1369)
);

BUFx10_ASAP7_75t_L g1370 ( 
.A(n_1244),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1265),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1271),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1278),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1305),
.B(n_1333),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1237),
.A2(n_1319),
.B1(n_1352),
.B2(n_1251),
.Y(n_1375)
);

AND2x4_ASAP7_75t_SL g1376 ( 
.A(n_1349),
.B(n_1363),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1247),
.B(n_1317),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1297),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_SL g1379 ( 
.A(n_1349),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1303),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1322),
.A2(n_1331),
.B(n_1321),
.Y(n_1381)
);

BUFx8_ASAP7_75t_L g1382 ( 
.A(n_1296),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1265),
.Y(n_1383)
);

OAI22x1_ASAP7_75t_SL g1384 ( 
.A1(n_1293),
.A2(n_1325),
.B1(n_1223),
.B2(n_1310),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1332),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1320),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1249),
.A2(n_1314),
.B1(n_1216),
.B2(n_1329),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1260),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1333),
.A2(n_1361),
.B1(n_1324),
.B2(n_1329),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1249),
.A2(n_1360),
.B1(n_1324),
.B2(n_1240),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1360),
.A2(n_1346),
.B1(n_1341),
.B2(n_1227),
.Y(n_1391)
);

BUFx2_ASAP7_75t_SL g1392 ( 
.A(n_1301),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1250),
.B(n_1325),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1221),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1257),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1211),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1341),
.A2(n_1346),
.B1(n_1227),
.B2(n_1361),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1299),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1274),
.Y(n_1399)
);

BUFx2_ASAP7_75t_SL g1400 ( 
.A(n_1343),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1238),
.A2(n_1229),
.B1(n_1277),
.B2(n_1261),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1238),
.A2(n_1277),
.B1(n_1280),
.B2(n_1295),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1255),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1236),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1276),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1335),
.A2(n_1357),
.B1(n_1342),
.B2(n_1353),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1284),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1266),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1272),
.B(n_1290),
.Y(n_1409)
);

CKINVDCx6p67_ASAP7_75t_R g1410 ( 
.A(n_1236),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_R g1411 ( 
.A1(n_1318),
.A2(n_1330),
.B1(n_1326),
.B2(n_1355),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1235),
.A2(n_1334),
.B1(n_1285),
.B2(n_1282),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1267),
.A2(n_1253),
.B1(n_1233),
.B2(n_1351),
.Y(n_1413)
);

OAI22x1_ASAP7_75t_L g1414 ( 
.A1(n_1338),
.A2(n_1323),
.B1(n_1287),
.B2(n_1348),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1252),
.A2(n_1243),
.B1(n_1263),
.B2(n_1289),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1267),
.A2(n_1253),
.B1(n_1233),
.B2(n_1350),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1288),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1233),
.A2(n_1337),
.B1(n_1354),
.B2(n_1315),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1298),
.A2(n_1313),
.B1(n_1304),
.B2(n_1300),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1215),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1235),
.A2(n_1347),
.B1(n_1339),
.B2(n_1279),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1294),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1259),
.A2(n_1275),
.B(n_1226),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1281),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1328),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1292),
.Y(n_1426)
);

BUFx4f_ASAP7_75t_L g1427 ( 
.A(n_1359),
.Y(n_1427)
);

BUFx4f_ASAP7_75t_SL g1428 ( 
.A(n_1359),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1264),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1286),
.B(n_1323),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1273),
.A2(n_1256),
.B1(n_1245),
.B2(n_1311),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_1254),
.Y(n_1432)
);

BUFx5_ASAP7_75t_L g1433 ( 
.A(n_1246),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1340),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1291),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1279),
.Y(n_1436)
);

INVx3_ASAP7_75t_SL g1437 ( 
.A(n_1339),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1268),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1323),
.A2(n_1347),
.B1(n_1259),
.B2(n_1269),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1239),
.B(n_1344),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1283),
.A2(n_1242),
.B1(n_1241),
.B2(n_1224),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1262),
.Y(n_1442)
);

CKINVDCx6p67_ASAP7_75t_R g1443 ( 
.A(n_1270),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1258),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1213),
.A2(n_1230),
.B1(n_1212),
.B2(n_1220),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1309),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1222),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1239),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1209),
.A2(n_1218),
.B1(n_1214),
.B2(n_1248),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1210),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1309),
.A2(n_1344),
.B1(n_1217),
.B2(n_1356),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1309),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1306),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1344),
.B(n_1219),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1307),
.A2(n_1308),
.B1(n_1316),
.B2(n_1336),
.Y(n_1455)
);

CKINVDCx6p67_ASAP7_75t_R g1456 ( 
.A(n_1219),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1231),
.A2(n_1345),
.B1(n_970),
.B2(n_1312),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1345),
.A2(n_1322),
.B(n_970),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1236),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1345),
.A2(n_1231),
.B1(n_1322),
.B2(n_1352),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1358),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_1358),
.Y(n_1463)
);

BUFx10_ASAP7_75t_L g1464 ( 
.A(n_1362),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1297),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1297),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1228),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1362),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1312),
.A2(n_970),
.B1(n_1055),
.B2(n_1134),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1345),
.A2(n_1055),
.B1(n_1225),
.B2(n_970),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1260),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1265),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1231),
.A2(n_1345),
.B1(n_970),
.B2(n_1312),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1362),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1247),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1234),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1302),
.A2(n_970),
.B1(n_1055),
.B2(n_1232),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1231),
.B(n_1305),
.Y(n_1483)
);

BUFx4f_ASAP7_75t_L g1484 ( 
.A(n_1371),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1431),
.A2(n_1451),
.B(n_1423),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1408),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1430),
.B(n_1440),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1441),
.A2(n_1449),
.B(n_1451),
.Y(n_1488)
);

CKINVDCx8_ASAP7_75t_R g1489 ( 
.A(n_1400),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1444),
.B(n_1435),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1454),
.B(n_1397),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1460),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1397),
.B(n_1414),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1369),
.B(n_1483),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1441),
.A2(n_1445),
.B(n_1409),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1387),
.B(n_1413),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1435),
.Y(n_1497)
);

INVx4_ASAP7_75t_L g1498 ( 
.A(n_1443),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1435),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1438),
.Y(n_1500)
);

INVxp33_ASAP7_75t_L g1501 ( 
.A(n_1393),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1445),
.A2(n_1409),
.B(n_1421),
.Y(n_1502)
);

CKINVDCx11_ASAP7_75t_R g1503 ( 
.A(n_1462),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1457),
.B(n_1474),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1380),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1452),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1471),
.A2(n_1367),
.B1(n_1458),
.B2(n_1457),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1442),
.B(n_1377),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1369),
.B(n_1483),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1470),
.A2(n_1477),
.B1(n_1482),
.B2(n_1480),
.Y(n_1511)
);

AO21x2_ASAP7_75t_L g1512 ( 
.A1(n_1431),
.A2(n_1453),
.B(n_1432),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1406),
.B(n_1415),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1391),
.B(n_1389),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1470),
.A2(n_1466),
.B1(n_1478),
.B2(n_1475),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1385),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1389),
.A2(n_1381),
.B(n_1458),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1413),
.B(n_1416),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1450),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_SL g1520 ( 
.A(n_1398),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1390),
.A2(n_1381),
.B(n_1401),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1468),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1377),
.B(n_1420),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1374),
.B(n_1461),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1474),
.A2(n_1439),
.A3(n_1374),
.B(n_1456),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1399),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1450),
.Y(n_1527)
);

AO21x2_ASAP7_75t_L g1528 ( 
.A1(n_1461),
.A2(n_1395),
.B(n_1417),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1375),
.B(n_1459),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1405),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1416),
.B(n_1418),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1447),
.A2(n_1429),
.B1(n_1436),
.B2(n_1450),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1402),
.A2(n_1364),
.B(n_1412),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1418),
.B(n_1448),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1376),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1433),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1437),
.B(n_1378),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1433),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1433),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1433),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1366),
.B(n_1479),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1433),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1455),
.Y(n_1543)
);

INVx4_ASAP7_75t_L g1544 ( 
.A(n_1434),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1426),
.B(n_1481),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1455),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1419),
.B(n_1386),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1410),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1373),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1419),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1465),
.Y(n_1551)
);

CKINVDCx11_ASAP7_75t_R g1552 ( 
.A(n_1463),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1467),
.B(n_1422),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1422),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1472),
.A2(n_1428),
.B1(n_1383),
.B2(n_1473),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1411),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1379),
.A2(n_1383),
.B(n_1473),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1427),
.B(n_1394),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1379),
.A2(n_1473),
.B(n_1371),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1427),
.A2(n_1424),
.B(n_1372),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_SL g1561 ( 
.A(n_1472),
.B(n_1392),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1472),
.B(n_1425),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1396),
.B(n_1476),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1487),
.B(n_1373),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1511),
.A2(n_1515),
.B1(n_1504),
.B2(n_1508),
.Y(n_1565)
);

AO32x2_ASAP7_75t_L g1566 ( 
.A1(n_1505),
.A2(n_1368),
.A3(n_1384),
.B1(n_1370),
.B2(n_1404),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1528),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1528),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1501),
.B(n_1464),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1495),
.B(n_1407),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1532),
.A2(n_1428),
.B1(n_1469),
.B2(n_1382),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1494),
.B(n_1382),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1529),
.A2(n_1388),
.B1(n_1403),
.B2(n_1464),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1495),
.B(n_1365),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1513),
.A2(n_1514),
.B(n_1521),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1537),
.B(n_1534),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1488),
.A2(n_1502),
.B(n_1543),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1513),
.A2(n_1556),
.B(n_1514),
.C(n_1524),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1505),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1535),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1506),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1492),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1543),
.A2(n_1546),
.B(n_1506),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1509),
.B(n_1491),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1521),
.A2(n_1513),
.B1(n_1533),
.B2(n_1556),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1516),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1507),
.Y(n_1587)
);

BUFx4f_ASAP7_75t_SL g1588 ( 
.A(n_1535),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1510),
.B(n_1554),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1531),
.A2(n_1496),
.B(n_1518),
.C(n_1493),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1523),
.B(n_1517),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1523),
.B(n_1517),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1485),
.A2(n_1517),
.B(n_1521),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1531),
.A2(n_1496),
.B(n_1518),
.C(n_1493),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_R g1595 ( 
.A(n_1503),
.B(n_1552),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_SL g1597 ( 
.A1(n_1555),
.A2(n_1527),
.B(n_1519),
.C(n_1563),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1489),
.A2(n_1484),
.B1(n_1521),
.B2(n_1533),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1498),
.B(n_1533),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1536),
.A2(n_1540),
.B(n_1538),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1485),
.A2(n_1546),
.B1(n_1561),
.B2(n_1553),
.C(n_1547),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1485),
.A2(n_1561),
.B1(n_1547),
.B2(n_1551),
.C(n_1545),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1533),
.A2(n_1527),
.B(n_1519),
.C(n_1560),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1541),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1489),
.A2(n_1484),
.B1(n_1548),
.B2(n_1549),
.Y(n_1606)
);

AO32x2_ASAP7_75t_L g1607 ( 
.A1(n_1497),
.A2(n_1499),
.A3(n_1525),
.B1(n_1512),
.B2(n_1544),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1535),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_R g1609 ( 
.A(n_1520),
.B(n_1548),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1549),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1507),
.A2(n_1500),
.B(n_1540),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1548),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1581),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1611),
.Y(n_1614)
);

OR2x2_ASAP7_75t_SL g1615 ( 
.A(n_1582),
.B(n_1522),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1581),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1611),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1490),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1611),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1587),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1577),
.B(n_1525),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1577),
.B(n_1525),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1584),
.B(n_1525),
.Y(n_1624)
);

CKINVDCx20_ASAP7_75t_R g1625 ( 
.A(n_1612),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1601),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1589),
.B(n_1512),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1596),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1583),
.B(n_1525),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1600),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1583),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1583),
.B(n_1486),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1500),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1592),
.B(n_1539),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1576),
.B(n_1542),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1570),
.B(n_1605),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1564),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1565),
.A2(n_1562),
.B1(n_1522),
.B2(n_1526),
.C(n_1530),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1599),
.B(n_1605),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1579),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1586),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1638),
.B(n_1603),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1613),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1637),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1613),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1629),
.B(n_1578),
.C(n_1602),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1624),
.B(n_1607),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1607),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1621),
.B(n_1622),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1621),
.B(n_1607),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1638),
.A2(n_1575),
.B1(n_1599),
.B2(n_1598),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1616),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1618),
.B(n_1574),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1621),
.B(n_1607),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1633),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1625),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1637),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1636),
.A2(n_1590),
.B1(n_1594),
.B2(n_1585),
.Y(n_1661)
);

INVx3_ASAP7_75t_SL g1662 ( 
.A(n_1615),
.Y(n_1662)
);

BUFx2_ASAP7_75t_SL g1663 ( 
.A(n_1631),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1629),
.A2(n_1593),
.B(n_1604),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1568),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1623),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1642),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1614),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1627),
.B(n_1567),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1623),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1614),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1620),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1620),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1617),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1635),
.B(n_1640),
.Y(n_1675)
);

OAI31xp33_ASAP7_75t_L g1676 ( 
.A1(n_1639),
.A2(n_1590),
.A3(n_1594),
.B(n_1578),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1617),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1615),
.B(n_1567),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1628),
.B(n_1574),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1644),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1669),
.B(n_1641),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1652),
.B(n_1628),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1644),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1665),
.B(n_1619),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1668),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1669),
.B(n_1641),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1662),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1659),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1665),
.B(n_1672),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1659),
.B(n_1595),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1646),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1648),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1662),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1659),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1653),
.B(n_1640),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1661),
.B(n_1569),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1657),
.B(n_1631),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1657),
.B(n_1631),
.Y(n_1704)
);

NOR2x1_ASAP7_75t_L g1705 ( 
.A(n_1647),
.B(n_1626),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1662),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1649),
.B(n_1635),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1668),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1668),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1656),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1648),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1649),
.B(n_1635),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1680),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1680),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1706),
.B(n_1660),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1705),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1684),
.B(n_1661),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1686),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1701),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1706),
.B(n_1656),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1683),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1683),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1686),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1692),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1691),
.B(n_1678),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1691),
.B(n_1678),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1705),
.B(n_1647),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1692),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1699),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1681),
.B(n_1658),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1696),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1699),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1699),
.B(n_1675),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1689),
.B(n_1660),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1693),
.B(n_1610),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1689),
.B(n_1660),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1696),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1681),
.B(n_1673),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.B(n_1702),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1697),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1687),
.B(n_1675),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1702),
.B(n_1673),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1697),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1675),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1711),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1698),
.B(n_1654),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1707),
.B(n_1660),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1707),
.B(n_1645),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1710),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1711),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1707),
.B(n_1645),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1645),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1715),
.B(n_1710),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_SL g1757 ( 
.A(n_1727),
.B(n_1690),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1719),
.B(n_1572),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1720),
.B(n_1710),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1715),
.B(n_1710),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1717),
.B(n_1732),
.Y(n_1761)
);

NAND2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1729),
.B(n_1580),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1749),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1734),
.B(n_1682),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1729),
.Y(n_1765)
);

NAND2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1732),
.B(n_1580),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1734),
.B(n_1682),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1721),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1721),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1736),
.B(n_1682),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1736),
.B(n_1688),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1720),
.B(n_1688),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1724),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1744),
.B(n_1685),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1748),
.B(n_1700),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1720),
.B(n_1688),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1724),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1745),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1750),
.B(n_1695),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1728),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1755),
.B(n_1703),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1685),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1747),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1716),
.A2(n_1664),
.B1(n_1704),
.B2(n_1703),
.C(n_1650),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1695),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1739),
.B(n_1685),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1728),
.Y(n_1787)
);

AND2x4_ASAP7_75t_SL g1788 ( 
.A(n_1753),
.B(n_1679),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1725),
.B(n_1694),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1733),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1725),
.B(n_1709),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1761),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1757),
.B(n_1735),
.Y(n_1793)
);

INVx6_ASAP7_75t_L g1794 ( 
.A(n_1759),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1783),
.A2(n_1781),
.B1(n_1775),
.B2(n_1778),
.C(n_1772),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1790),
.B(n_1726),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1768),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1768),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1784),
.B(n_1573),
.C(n_1664),
.D(n_1597),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1765),
.B(n_1573),
.C(n_1597),
.D(n_1726),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

O2A1O1Ixp5_ASAP7_75t_L g1802 ( 
.A1(n_1765),
.A2(n_1718),
.B(n_1723),
.C(n_1731),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1765),
.B(n_1753),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1789),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1758),
.B(n_1764),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1764),
.B(n_1754),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1767),
.B(n_1754),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1769),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1789),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1773),
.Y(n_1811)
);

NAND2x1p5_ASAP7_75t_L g1812 ( 
.A(n_1759),
.B(n_1608),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1776),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1773),
.A2(n_1571),
.B(n_1604),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1777),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1762),
.A2(n_1751),
.B1(n_1738),
.B2(n_1730),
.C(n_1679),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1767),
.B(n_1741),
.Y(n_1817)
);

NOR3xp33_ASAP7_75t_L g1818 ( 
.A(n_1777),
.B(n_1544),
.C(n_1751),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1794),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1805),
.B(n_1772),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1804),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1797),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1814),
.A2(n_1766),
.B1(n_1762),
.B2(n_1776),
.Y(n_1823)
);

OA211x2_ASAP7_75t_L g1824 ( 
.A1(n_1793),
.A2(n_1667),
.B(n_1762),
.C(n_1766),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1792),
.A2(n_1562),
.B1(n_1766),
.B2(n_1588),
.Y(n_1825)
);

OAI22x1_ASAP7_75t_SL g1826 ( 
.A1(n_1810),
.A2(n_1763),
.B1(n_1787),
.B2(n_1780),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1813),
.B(n_1776),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1814),
.A2(n_1788),
.B1(n_1771),
.B2(n_1770),
.Y(n_1828)
);

O2A1O1Ixp5_ASAP7_75t_L g1829 ( 
.A1(n_1802),
.A2(n_1763),
.B(n_1774),
.C(n_1760),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1798),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1792),
.A2(n_1780),
.B(n_1787),
.C(n_1774),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1794),
.B(n_1770),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1794),
.Y(n_1833)
);

AOI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1801),
.A2(n_1811),
.B(n_1809),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1806),
.B(n_1788),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1812),
.B(n_1771),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1815),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_L g1838 ( 
.A(n_1796),
.B(n_1609),
.Y(n_1838)
);

AOI32xp33_ASAP7_75t_L g1839 ( 
.A1(n_1818),
.A2(n_1760),
.A3(n_1756),
.B1(n_1785),
.B2(n_1779),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1803),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1829),
.A2(n_1799),
.B(n_1802),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1834),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1821),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1826),
.B(n_1800),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1819),
.B(n_1795),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1832),
.B(n_1820),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1819),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1820),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1833),
.B(n_1807),
.Y(n_1849)
);

NAND4xp25_ASAP7_75t_L g1850 ( 
.A(n_1835),
.B(n_1816),
.C(n_1808),
.D(n_1817),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1832),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1835),
.A2(n_1812),
.B(n_1756),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1822),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1846),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1847),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1847),
.B(n_1833),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1851),
.B(n_1840),
.Y(n_1857)
);

NOR2xp67_ASAP7_75t_L g1858 ( 
.A(n_1852),
.B(n_1823),
.Y(n_1858)
);

NOR2x1_ASAP7_75t_L g1859 ( 
.A(n_1842),
.B(n_1841),
.Y(n_1859)
);

OAI321xp33_ASAP7_75t_L g1860 ( 
.A1(n_1844),
.A2(n_1828),
.A3(n_1839),
.B1(n_1825),
.B2(n_1831),
.C(n_1836),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1844),
.B(n_1827),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1848),
.B(n_1836),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1845),
.B(n_1782),
.Y(n_1863)
);

O2A1O1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1860),
.A2(n_1843),
.B(n_1838),
.C(n_1853),
.Y(n_1864)
);

AOI221x1_ASAP7_75t_SL g1865 ( 
.A1(n_1862),
.A2(n_1849),
.B1(n_1850),
.B2(n_1837),
.C(n_1830),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1863),
.A2(n_1838),
.B1(n_1824),
.B2(n_1786),
.C(n_1782),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1861),
.A2(n_1786),
.B1(n_1791),
.B2(n_1785),
.C(n_1779),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1855),
.A2(n_1791),
.B1(n_1718),
.B2(n_1723),
.C(n_1746),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1854),
.B(n_1749),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1866),
.A2(n_1859),
.B(n_1858),
.C(n_1856),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1864),
.A2(n_1857),
.B(n_1562),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1867),
.A2(n_1606),
.B1(n_1588),
.B2(n_1663),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1869),
.A2(n_1868),
.B1(n_1865),
.B2(n_1663),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1869),
.B(n_1703),
.Y(n_1874)
);

NOR2xp67_ASAP7_75t_L g1875 ( 
.A(n_1869),
.B(n_1731),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1867),
.A2(n_1743),
.B1(n_1746),
.B2(n_1713),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1870),
.B(n_1562),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1874),
.Y(n_1878)
);

NAND4xp75_ASAP7_75t_L g1879 ( 
.A(n_1871),
.B(n_1743),
.C(n_1752),
.D(n_1740),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1873),
.B(n_1704),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1875),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1872),
.B(n_1562),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1881),
.B(n_1544),
.Y(n_1883)
);

OAI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1877),
.A2(n_1876),
.B1(n_1558),
.B2(n_1738),
.C(n_1737),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1878),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1883),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1886),
.A2(n_1885),
.B1(n_1882),
.B2(n_1884),
.Y(n_1887)
);

OAI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1887),
.A2(n_1880),
.B1(n_1879),
.B2(n_1714),
.Y(n_1888)
);

OA21x2_ASAP7_75t_L g1889 ( 
.A1(n_1887),
.A2(n_1722),
.B(n_1709),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1889),
.A2(n_1558),
.B1(n_1609),
.B2(n_1708),
.Y(n_1890)
);

CKINVDCx20_ASAP7_75t_R g1891 ( 
.A(n_1888),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1891),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1890),
.A2(n_1742),
.B1(n_1730),
.B2(n_1686),
.Y(n_1893)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1894 ( 
.A1(n_1892),
.A2(n_1655),
.B(n_1666),
.C(n_1670),
.D(n_1566),
.Y(n_1894)
);

NAND2x1_ASAP7_75t_L g1895 ( 
.A(n_1894),
.B(n_1893),
.Y(n_1895)
);

OAI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1895),
.A2(n_1708),
.B1(n_1742),
.B2(n_1709),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1896),
.A2(n_1708),
.B1(n_1674),
.B2(n_1671),
.C(n_1677),
.Y(n_1897)
);

OA22x2_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1671),
.B1(n_1674),
.B2(n_1677),
.Y(n_1898)
);


endmodule