module fake_jpeg_24741_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx10_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_25),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_15),
.B(n_26),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_20),
.B(n_27),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.C(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_77),
.C(n_19),
.Y(n_95)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_61),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_20),
.B(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_66),
.B1(n_24),
.B2(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_38),
.B1(n_32),
.B2(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_29),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_49),
.B(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_33),
.C(n_36),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_83),
.B1(n_79),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_71),
.B1(n_63),
.B2(n_74),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_89),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_51),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_36),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_106),
.B1(n_46),
.B2(n_81),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_82),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_111),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_60),
.B(n_59),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_114),
.B(n_116),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_58),
.B(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_78),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_65),
.B(n_46),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_87),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_1),
.C(n_2),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_98),
.Y(n_125)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_130),
.A3(n_18),
.B1(n_104),
.B2(n_28),
.C(n_21),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_88),
.B(n_30),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_101),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_42),
.B1(n_81),
.B2(n_19),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_30),
.C(n_21),
.Y(n_137)
);

OAI321xp33_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_100),
.A3(n_106),
.B1(n_112),
.B2(n_116),
.C(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_127),
.C(n_124),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_8),
.C(n_14),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_117),
.B1(n_119),
.B2(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_135),
.B1(n_129),
.B2(n_131),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_119),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_122),
.B(n_144),
.Y(n_153)
);

OAI21x1_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_143),
.B(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_155),
.C(n_18),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_156),
.B1(n_150),
.B2(n_145),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.C(n_160),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_18),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_7),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_9),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_8),
.A3(n_10),
.B1(n_9),
.B2(n_28),
.C1(n_5),
.C2(n_4),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_159),
.B(n_3),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_165),
.B1(n_2),
.B2(n_3),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_2),
.B(n_3),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.C(n_162),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_4),
.Y(n_169)
);


endmodule