module fake_jpeg_29858_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_22),
.B(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_30),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_36),
.B1(n_15),
.B2(n_27),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_15),
.B(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_28),
.C(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_36),
.C(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

OAI22x1_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_41),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_R g47 ( 
.A1(n_43),
.A2(n_13),
.B(n_11),
.C(n_17),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_34),
.C(n_33),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_46),
.C(n_47),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_28),
.C(n_43),
.Y(n_49)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_7),
.B(n_5),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_48),
.B(n_7),
.Y(n_51)
);


endmodule