module real_jpeg_2968_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_1),
.B(n_53),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_1),
.B(n_51),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_2),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_2),
.B(n_26),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_3),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_3),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_3),
.B(n_62),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_3),
.B(n_28),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_5),
.B(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_28),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_51),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_5),
.B(n_26),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_11),
.B(n_28),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_12),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_12),
.B(n_62),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_12),
.B(n_53),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_14),
.B(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_14),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_14),
.B(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_14),
.B(n_28),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_14),
.B(n_26),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_93),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_20),
.B(n_93),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_57),
.C(n_82),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_21),
.B(n_205),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_21),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_38),
.CI(n_42),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_38),
.C(n_42),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.C(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_23),
.A2(n_24),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_25),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_25),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_27),
.A2(n_72),
.B1(n_75),
.B2(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_29),
.B(n_128),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_31),
.B(n_35),
.Y(n_201)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_41),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_41),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_50),
.C(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_44),
.B(n_73),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_44),
.B(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_45),
.B(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_56),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_57),
.B(n_82),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_81),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_70),
.C(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_66),
.C(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.C(n_80),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_91),
.Y(n_82)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_83),
.B(n_87),
.CI(n_91),
.CON(n_195),
.SN(n_195)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_90),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_141),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_93),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_115),
.CI(n_116),
.CON(n_93),
.SN(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_126),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_203),
.B(n_207),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_191),
.B(n_202),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_163),
.B(n_190),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_154),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_154),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_138),
.CI(n_139),
.CON(n_155),
.SN(n_155)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_150),
.C(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_162),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_187),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_155),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_157),
.B1(n_162),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_184),
.B(n_189),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_175),
.B(n_183),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_171),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_198),
.C(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_206),
.Y(n_207)
);


endmodule