module real_aes_17082_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_656;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g660 ( .A(n_0), .Y(n_660) );
AND2x2_ASAP7_75t_L g491 ( .A(n_1), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g506 ( .A(n_1), .Y(n_506) );
AND2x2_ASAP7_75t_L g515 ( .A(n_1), .B(n_60), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_2), .Y(n_652) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g112 ( .A(n_4), .B(n_113), .Y(n_112) );
AOI21xp33_ASAP7_75t_L g537 ( .A1(n_5), .A2(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g577 ( .A(n_5), .Y(n_577) );
INVx1_ASAP7_75t_L g553 ( .A(n_6), .Y(n_553) );
INVx1_ASAP7_75t_L g575 ( .A(n_6), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_7), .A2(n_49), .B1(n_508), .B2(n_513), .Y(n_507) );
INVx1_ASAP7_75t_L g578 ( .A(n_7), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_8), .A2(n_61), .B1(n_495), .B2(n_498), .C(n_503), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_8), .A2(n_73), .B1(n_550), .B2(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g560 ( .A(n_9), .Y(n_560) );
OAI21x1_ASAP7_75t_L g93 ( .A1(n_10), .A2(n_24), .B(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_11), .B(n_198), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_12), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_13), .B(n_162), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_14), .B(n_91), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_15), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_16), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_17), .Y(n_137) );
INVx2_ASAP7_75t_L g562 ( .A(n_18), .Y(n_562) );
INVx1_ASAP7_75t_L g594 ( .A(n_18), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_18), .B(n_560), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_19), .B(n_113), .Y(n_183) );
INVx2_ASAP7_75t_L g669 ( .A(n_20), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_21), .B(n_187), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_22), .B(n_141), .Y(n_200) );
INVx1_ASAP7_75t_L g519 ( .A(n_23), .Y(n_519) );
AND2x2_ASAP7_75t_L g140 ( .A(n_25), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_26), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_27), .B(n_162), .Y(n_161) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_28), .A2(n_73), .B1(n_486), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_28), .A2(n_61), .B1(n_585), .B2(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g517 ( .A(n_29), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_30), .B(n_225), .Y(n_224) );
BUFx3_ASAP7_75t_L g554 ( .A(n_31), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_32), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_33), .A2(n_102), .B(n_111), .C(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g94 ( .A(n_34), .Y(n_94) );
AND2x4_ASAP7_75t_L g116 ( .A(n_35), .B(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_35), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_36), .A2(n_38), .B1(n_138), .B2(n_210), .Y(n_209) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_37), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_39), .B(n_91), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_40), .B(n_141), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_41), .Y(n_139) );
XNOR2xp5_ASAP7_75t_L g479 ( .A(n_42), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_43), .B(n_138), .Y(n_186) );
INVx1_ASAP7_75t_L g117 ( .A(n_44), .Y(n_117) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_45), .A2(n_64), .B1(n_522), .B2(n_526), .C(n_531), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_45), .A2(n_64), .B1(n_604), .B2(n_608), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_46), .Y(n_212) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_47), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_48), .B(n_91), .Y(n_188) );
INVx1_ASAP7_75t_L g599 ( .A(n_49), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_50), .B(n_98), .Y(n_160) );
NAND3xp33_ASAP7_75t_L g194 ( .A(n_51), .B(n_168), .C(n_187), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_52), .B(n_98), .Y(n_97) );
INVx2_ASAP7_75t_L g104 ( .A(n_53), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_54), .B(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_54), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_55), .B(n_113), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_56), .A2(n_74), .B1(n_625), .B2(n_635), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_57), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g623 ( .A(n_58), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_59), .A2(n_67), .B1(n_162), .B2(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g492 ( .A(n_60), .Y(n_492) );
BUFx3_ASAP7_75t_L g505 ( .A(n_60), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_62), .B(n_113), .Y(n_221) );
NAND2xp33_ASAP7_75t_SL g153 ( .A(n_63), .B(n_101), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_65), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g547 ( .A(n_66), .Y(n_547) );
INVx1_ASAP7_75t_L g557 ( .A(n_66), .Y(n_557) );
INVx1_ASAP7_75t_L g568 ( .A(n_66), .Y(n_568) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_68), .Y(n_662) );
NAND2xp33_ASAP7_75t_L g100 ( .A(n_69), .B(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_70), .B(n_141), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g149 ( .A(n_71), .B(n_101), .C(n_148), .Y(n_149) );
INVx1_ASAP7_75t_L g678 ( .A(n_71), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_72), .B(n_98), .Y(n_185) );
OAI211xp5_ASAP7_75t_L g483 ( .A1(n_74), .A2(n_484), .B(n_493), .C(n_516), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_75), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_76), .B(n_162), .Y(n_165) );
AOI21xp33_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_470), .B(n_478), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
AND2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_350), .Y(n_81) );
NOR3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_258), .C(n_309), .Y(n_82) );
OAI211xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_172), .B(n_227), .C(n_245), .Y(n_83) );
NAND3x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_118), .C(n_155), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g318 ( .A(n_86), .B(n_297), .Y(n_318) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND3x2_ASAP7_75t_L g238 ( .A(n_87), .B(n_239), .C(n_243), .Y(n_238) );
AND2x2_ASAP7_75t_L g273 ( .A(n_87), .B(n_257), .Y(n_273) );
AND2x2_ASAP7_75t_L g279 ( .A(n_87), .B(n_275), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_87), .B(n_243), .Y(n_420) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g322 ( .A(n_88), .B(n_243), .Y(n_322) );
AND2x2_ASAP7_75t_L g333 ( .A(n_88), .B(n_287), .Y(n_333) );
BUFx2_ASAP7_75t_L g339 ( .A(n_88), .Y(n_339) );
NAND2x1_ASAP7_75t_L g355 ( .A(n_88), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g361 ( .A(n_88), .B(n_362), .Y(n_361) );
INVx4_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx2_ASAP7_75t_L g255 ( .A(n_89), .Y(n_255) );
AND2x2_ASAP7_75t_L g286 ( .A(n_89), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g306 ( .A(n_89), .B(n_242), .Y(n_306) );
INVx1_ASAP7_75t_L g377 ( .A(n_89), .Y(n_377) );
AND2x4_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
INVx4_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x4_ASAP7_75t_SL g114 ( .A(n_92), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g144 ( .A(n_92), .Y(n_144) );
INVx2_ASAP7_75t_L g178 ( .A(n_92), .Y(n_178) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
OAI21x1_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_105), .B(n_114), .Y(n_95) );
AOI21xp5_ASAP7_75t_L g96 ( .A1(n_97), .A2(n_100), .B(n_102), .Y(n_96) );
OAI22xp33_ASAP7_75t_L g136 ( .A1(n_98), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_136) );
INVx3_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_99), .Y(n_101) );
INVx1_ASAP7_75t_L g111 ( .A(n_99), .Y(n_111) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_99), .Y(n_113) );
INVx2_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_99), .Y(n_138) );
INVx1_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_99), .Y(n_168) );
INVx1_ASAP7_75t_L g182 ( .A(n_99), .Y(n_182) );
INVx1_ASAP7_75t_L g210 ( .A(n_99), .Y(n_210) );
INVx2_ASAP7_75t_L g225 ( .A(n_101), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_102), .A2(n_151), .B(n_153), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_102), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_102), .A2(n_181), .B(n_183), .Y(n_180) );
BUFx4f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g109 ( .A(n_104), .Y(n_109) );
INVx1_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
BUFx8_ASAP7_75t_L g187 ( .A(n_104), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_108), .B1(n_110), .B2(n_112), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_107), .A2(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_113), .A2(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g198 ( .A(n_113), .Y(n_198) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_115), .A2(n_146), .B(n_150), .Y(n_145) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_115), .A2(n_159), .B(n_164), .Y(n_158) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_115), .A2(n_180), .B(n_184), .Y(n_179) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_115), .A2(n_192), .B(n_195), .Y(n_191) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_115), .A2(n_218), .B(n_222), .Y(n_217) );
BUFx10_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx10_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_117), .Y(n_647) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OR2x6_ASAP7_75t_L g354 ( .A(n_119), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g256 ( .A(n_120), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_120), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_143), .Y(n_120) );
INVx2_ASAP7_75t_L g244 ( .A(n_121), .Y(n_244) );
INVx1_ASAP7_75t_L g298 ( .A(n_121), .Y(n_298) );
AOI21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_128), .B(n_140), .Y(n_121) );
NOR2xp67_ASAP7_75t_SL g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_124), .A2(n_127), .A3(n_205), .B(n_211), .Y(n_204) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g142 ( .A(n_125), .Y(n_142) );
INVx2_ASAP7_75t_L g213 ( .A(n_125), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_126), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_131), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_131), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_134), .A2(n_206), .B1(n_208), .B2(n_209), .Y(n_205) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_138), .A2(n_193), .B(n_194), .Y(n_192) );
INVx2_ASAP7_75t_L g207 ( .A(n_138), .Y(n_207) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
INVx1_ASAP7_75t_L g242 ( .A(n_143), .Y(n_242) );
INVx2_ASAP7_75t_L g276 ( .A(n_143), .Y(n_276) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_154), .Y(n_143) );
INVx1_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_156), .A2(n_458), .B(n_462), .Y(n_457) );
BUFx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g297 ( .A(n_157), .B(n_298), .Y(n_297) );
OAI21xp33_ASAP7_75t_SL g157 ( .A1(n_158), .A2(n_170), .B(n_171), .Y(n_157) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_158), .A2(n_170), .B(n_171), .Y(n_241) );
INVx1_ASAP7_75t_L g476 ( .A(n_162), .Y(n_476) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_169), .Y(n_164) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI21x1_ASAP7_75t_L g216 ( .A1(n_170), .A2(n_217), .B(n_226), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_170), .A2(n_217), .B(n_226), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_201), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_174), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp67_ASAP7_75t_L g175 ( .A(n_176), .B(n_189), .Y(n_175) );
INVx3_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
AND2x2_ASAP7_75t_L g382 ( .A(n_176), .B(n_190), .Y(n_382) );
BUFx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g271 ( .A(n_177), .Y(n_271) );
OAI21x1_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_188), .Y(n_177) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_178), .A2(n_191), .B(n_200), .Y(n_190) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_178), .A2(n_179), .B(n_188), .Y(n_250) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_178), .A2(n_191), .B(n_200), .Y(n_253) );
INVx2_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
INVx6_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_L g218 ( .A1(n_187), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
AND2x4_ASAP7_75t_L g236 ( .A(n_189), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g295 ( .A(n_190), .Y(n_295) );
AND2x2_ASAP7_75t_L g312 ( .A(n_190), .B(n_204), .Y(n_312) );
AND2x2_ASAP7_75t_L g424 ( .A(n_190), .B(n_301), .Y(n_424) );
AND2x2_ASAP7_75t_L g446 ( .A(n_190), .B(n_215), .Y(n_446) );
AOI21x1_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .Y(n_195) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_203), .B(n_214), .Y(n_202) );
INVx1_ASAP7_75t_L g266 ( .A(n_203), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_203), .B(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g237 ( .A(n_204), .Y(n_237) );
OR2x2_ASAP7_75t_L g252 ( .A(n_204), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g270 ( .A(n_204), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g324 ( .A(n_204), .B(n_250), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_204), .B(n_253), .Y(n_366) );
OR2x2_ASAP7_75t_L g436 ( .A(n_204), .B(n_250), .Y(n_436) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_208), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx1_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
AND2x4_ASAP7_75t_L g282 ( .A(n_214), .B(n_236), .Y(n_282) );
AND2x2_ASAP7_75t_L g428 ( .A(n_214), .B(n_270), .Y(n_428) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx3_ASAP7_75t_L g230 ( .A(n_215), .Y(n_230) );
AND2x2_ASAP7_75t_L g290 ( .A(n_215), .B(n_249), .Y(n_290) );
INVx1_ASAP7_75t_L g343 ( .A(n_215), .Y(n_343) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_215), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_215), .B(n_253), .Y(n_384) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_215), .Y(n_394) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_231), .B(n_238), .Y(n_227) );
AND2x2_ASAP7_75t_L g426 ( .A(n_228), .B(n_331), .Y(n_426) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g293 ( .A(n_229), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_229), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_230), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g373 ( .A(n_230), .B(n_236), .Y(n_373) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_235), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g371 ( .A(n_235), .B(n_312), .Y(n_371) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_235), .Y(n_402) );
INVx2_ASAP7_75t_L g336 ( .A(n_236), .Y(n_336) );
AND2x2_ASAP7_75t_L g465 ( .A(n_237), .B(n_250), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_238), .A2(n_320), .B1(n_321), .B2(n_323), .C(n_325), .Y(n_319) );
AND2x2_ASAP7_75t_L g260 ( .A(n_239), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g321 ( .A(n_239), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
INVx2_ASAP7_75t_L g257 ( .A(n_240), .Y(n_257) );
OR2x2_ASAP7_75t_L g390 ( .A(n_240), .B(n_275), .Y(n_390) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
INVxp67_ASAP7_75t_L g317 ( .A(n_242), .Y(n_317) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g261 ( .A(n_244), .Y(n_261) );
AND2x2_ASAP7_75t_L g274 ( .A(n_244), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g281 ( .A(n_244), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
AND2x2_ASAP7_75t_L g404 ( .A(n_246), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g331 ( .A(n_248), .B(n_312), .Y(n_331) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_248), .Y(n_461) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g289 ( .A(n_251), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g439 ( .A(n_251), .Y(n_439) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g327 ( .A(n_252), .Y(n_327) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_252), .Y(n_401) );
AND2x2_ASAP7_75t_L g300 ( .A(n_253), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_254), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g296 ( .A(n_255), .B(n_297), .Y(n_296) );
OAI21xp33_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_278), .B(n_282), .Y(n_277) );
NAND4xp25_ASAP7_75t_L g258 ( .A(n_259), .B(n_277), .C(n_283), .D(n_291), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B(n_267), .Y(n_259) );
INVx2_ASAP7_75t_L g348 ( .A(n_261), .Y(n_348) );
AND2x2_ASAP7_75t_L g359 ( .A(n_261), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g369 ( .A(n_261), .B(n_286), .Y(n_369) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g445 ( .A(n_266), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_272), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI33xp33_ASAP7_75t_L g415 ( .A1(n_269), .A2(n_306), .A3(n_416), .B1(n_418), .B2(n_421), .B3(n_422), .Y(n_415) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g448 ( .A(n_270), .B(n_300), .Y(n_448) );
BUFx2_ASAP7_75t_L g303 ( .A(n_271), .Y(n_303) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_274), .B(n_286), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_275), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
INVx1_ASAP7_75t_L g362 ( .A(n_276), .Y(n_362) );
AND2x2_ASAP7_75t_L g376 ( .A(n_276), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g347 ( .A(n_279), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g399 ( .A(n_279), .Y(n_399) );
INVx1_ASAP7_75t_L g409 ( .A(n_280), .Y(n_409) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g285 ( .A(n_281), .Y(n_285) );
INVx1_ASAP7_75t_L g391 ( .A(n_281), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
OR2x2_ASAP7_75t_L g374 ( .A(n_285), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g345 ( .A(n_286), .B(n_329), .Y(n_345) );
AND2x2_ASAP7_75t_L g308 ( .A(n_287), .B(n_298), .Y(n_308) );
INVx2_ASAP7_75t_L g356 ( .A(n_287), .Y(n_356) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_296), .B1(n_299), .B2(n_304), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_294), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_296), .A2(n_379), .B1(n_383), .B2(n_385), .C(n_387), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_297), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g433 ( .A(n_297), .Y(n_433) );
AND2x2_ASAP7_75t_L g452 ( .A(n_297), .B(n_376), .Y(n_452) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g421 ( .A(n_300), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_300), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g407 ( .A(n_301), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_302), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g395 ( .A(n_302), .B(n_336), .Y(n_395) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_304), .A2(n_450), .B1(n_452), .B2(n_453), .Y(n_449) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OR2x2_ASAP7_75t_L g466 ( .A(n_307), .B(n_361), .Y(n_466) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g414 ( .A(n_308), .B(n_376), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B(n_319), .C(n_334), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
AND2x2_ASAP7_75t_L g393 ( .A(n_312), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g386 ( .A(n_318), .Y(n_386) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_324), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g383 ( .A(n_324), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g417 ( .A(n_324), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_324), .B(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B1(n_330), .B2(n_332), .Y(n_325) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI21xp33_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_337), .B(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_346), .B2(n_349), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_342), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_SL g427 ( .A1(n_345), .A2(n_428), .B(n_429), .C(n_437), .Y(n_427) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g442 ( .A(n_348), .B(n_376), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_410), .C(n_440), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_378), .C(n_398), .Y(n_351) );
O2A1O1Ixp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_357), .B(n_363), .C(n_367), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp33_ASAP7_75t_SL g429 ( .A1(n_355), .A2(n_430), .B1(n_432), .B2(n_434), .Y(n_429) );
INVx1_ASAP7_75t_SL g419 ( .A(n_356), .Y(n_419) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g432 ( .A(n_361), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_372), .B2(n_374), .Y(n_367) );
NAND2xp33_ASAP7_75t_SL g385 ( .A(n_368), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g451 ( .A(n_373), .Y(n_451) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g405 ( .A(n_376), .B(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_380), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g456 ( .A(n_381), .Y(n_456) );
INVx1_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B1(n_395), .B2(n_396), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2x1p5_ASAP7_75t_SL g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g397 ( .A(n_390), .Y(n_397) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g403 ( .A(n_394), .Y(n_403) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B(n_404), .C(n_408), .Y(n_398) );
NOR3x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .C(n_403), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_405), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_425), .C(n_427), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_449), .C(n_457), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx5_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AO21x1_ASAP7_75t_L g691 ( .A1(n_474), .A2(n_646), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_643), .B2(n_648), .C(n_684), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_480), .A2(n_685), .B1(n_686), .B2(n_689), .Y(n_684) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND4x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_548), .C(n_614), .D(n_638), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_521), .B(n_544), .Y(n_482) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_491), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx3_ASAP7_75t_L g513 ( .A(n_487), .Y(n_513) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x2_ASAP7_75t_L g497 ( .A(n_488), .B(n_490), .Y(n_497) );
INVx2_ASAP7_75t_L g502 ( .A(n_488), .Y(n_502) );
INVx1_ASAP7_75t_L g512 ( .A(n_488), .Y(n_512) );
BUFx2_ASAP7_75t_L g529 ( .A(n_488), .Y(n_529) );
NAND2x1_ASAP7_75t_L g536 ( .A(n_488), .B(n_490), .Y(n_536) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g501 ( .A(n_490), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g511 ( .A(n_490), .Y(n_511) );
INVx1_ASAP7_75t_L g633 ( .A(n_490), .Y(n_633) );
AND2x2_ASAP7_75t_L g518 ( .A(n_491), .B(n_510), .Y(n_518) );
AND2x4_ASAP7_75t_L g520 ( .A(n_491), .B(n_500), .Y(n_520) );
AND2x4_ASAP7_75t_SL g525 ( .A(n_491), .B(n_496), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_507), .B(n_514), .Y(n_493) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x6_ASAP7_75t_L g514 ( .A(n_496), .B(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g538 ( .A(n_501), .Y(n_538) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g541 ( .A(n_505), .Y(n_541) );
AND2x4_ASAP7_75t_L g540 ( .A(n_506), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g543 ( .A(n_509), .Y(n_543) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_510), .B(n_515), .Y(n_622) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_515), .B(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_517), .A2(n_519), .B1(n_639), .B2(n_642), .Y(n_638) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI211xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_537), .C(n_542), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_532), .A2(n_571), .B1(n_596), .B2(n_599), .C(n_600), .Y(n_595) );
INVx5_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_563), .C(n_603), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g602 ( .A(n_551), .Y(n_602) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
INVx1_ASAP7_75t_L g613 ( .A(n_552), .Y(n_613) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_553), .B(n_554), .Y(n_583) );
INVx1_ASAP7_75t_L g629 ( .A(n_553), .Y(n_629) );
INVx2_ASAP7_75t_L g576 ( .A(n_554), .Y(n_576) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_554), .Y(n_607) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_555), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_SL g609 ( .A(n_555), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
OR2x2_ASAP7_75t_L g621 ( .A(n_556), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g593 ( .A(n_557), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_558), .B(n_587), .Y(n_636) );
AND2x6_ASAP7_75t_L g668 ( .A(n_558), .B(n_605), .Y(n_668) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
NAND3x1_ASAP7_75t_L g592 ( .A(n_559), .B(n_593), .C(n_594), .Y(n_592) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp33_ASAP7_75t_SL g569 ( .A(n_560), .B(n_562), .Y(n_569) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_570), .B1(n_590), .B2(n_595), .Y(n_563) );
BUFx8_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
OR2x2_ASAP7_75t_L g619 ( .A(n_566), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_L g634 ( .A(n_567), .Y(n_634) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g674 ( .A(n_569), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_577), .B1(n_578), .B2(n_579), .C(n_584), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g642 ( .A(n_572), .B(n_641), .Y(n_642) );
BUFx8_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g589 ( .A(n_575), .Y(n_589) );
AND2x4_ASAP7_75t_L g587 ( .A(n_576), .B(n_588), .Y(n_587) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g598 ( .A(n_583), .Y(n_598) );
INVx8_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
INVx8_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_591), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
CKINVDCx8_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g618 ( .A(n_598), .Y(n_618) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_605), .B(n_671), .C(n_674), .Y(n_670) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_607), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_623), .B(n_624), .Y(n_614) );
INVx8_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OR2x2_ASAP7_75t_L g626 ( .A(n_619), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g641 ( .A(n_619), .Y(n_641) );
AND2x4_ASAP7_75t_L g625 ( .A(n_626), .B(n_630), .Y(n_625) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g637 ( .A(n_634), .Y(n_637) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x4_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
BUFx4f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g676 ( .A(n_645), .Y(n_676) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_647), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g692 ( .A(n_647), .B(n_676), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_663), .B1(n_677), .B2(n_679), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_649), .A2(n_664), .B1(n_677), .B2(n_680), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_658), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_655), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx12f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx8_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_670), .C(n_675), .Y(n_666) );
AND2x2_ASAP7_75t_L g683 ( .A(n_667), .B(n_670), .Y(n_683) );
INVx4_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx3_ASAP7_75t_L g673 ( .A(n_669), .Y(n_673) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g682 ( .A(n_675), .Y(n_682) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x6_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
endmodule