module fake_jpeg_26045_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_30),
.B1(n_32),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_19),
.B1(n_33),
.B2(n_26),
.Y(n_96)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_42),
.B1(n_37),
.B2(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_39),
.B1(n_36),
.B2(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_58),
.Y(n_95)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_18),
.B(n_17),
.C(n_20),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_24),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_61),
.B1(n_24),
.B2(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_24),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_72),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_18),
.B1(n_29),
.B2(n_33),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_42),
.B1(n_31),
.B2(n_27),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_91),
.B1(n_53),
.B2(n_54),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_39),
.B1(n_34),
.B2(n_35),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_89),
.B1(n_96),
.B2(n_26),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_36),
.B1(n_40),
.B2(n_38),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_40),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_98),
.B(n_26),
.C(n_36),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_97),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_40),
.B1(n_35),
.B2(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_29),
.B1(n_33),
.B2(n_19),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_26),
.B1(n_31),
.B2(n_27),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_47),
.B1(n_53),
.B2(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_47),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_12),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_40),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_104),
.B1(n_109),
.B2(n_115),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_85),
.A3(n_67),
.B1(n_66),
.B2(n_95),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_88),
.A3(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_61),
.C(n_38),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_117),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_27),
.B1(n_31),
.B2(n_38),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_38),
.B1(n_36),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_119),
.B1(n_115),
.B2(n_100),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_36),
.B1(n_25),
.B2(n_23),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_89),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_36),
.B1(n_62),
.B2(n_26),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_65),
.B1(n_74),
.B2(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_92),
.B1(n_82),
.B2(n_93),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_92),
.B1(n_75),
.B2(n_98),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_98),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_143),
.B(n_145),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_70),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_141),
.Y(n_188)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_69),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_14),
.B(n_15),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_15),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_69),
.B1(n_94),
.B2(n_86),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_150),
.B1(n_152),
.B2(n_108),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_36),
.B1(n_71),
.B2(n_25),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_111),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_71),
.B1(n_25),
.B2(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_64),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_114),
.B1(n_116),
.B2(n_112),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_108),
.B(n_64),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_71),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_106),
.B(n_8),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_178),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_126),
.B1(n_117),
.B2(n_110),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_171),
.B1(n_183),
.B2(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_172),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_110),
.B(n_114),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_173),
.B(n_174),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_112),
.B(n_116),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_180),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_184),
.B1(n_185),
.B2(n_3),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_157),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_122),
.B1(n_127),
.B2(n_111),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_179),
.A2(n_140),
.B1(n_149),
.B2(n_138),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_122),
.B(n_78),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_181),
.A2(n_192),
.B(n_6),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_127),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_0),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_22),
.B1(n_64),
.B2(n_2),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_11),
.C(n_9),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_147),
.C(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_5),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_155),
.B(n_129),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_194),
.A2(n_195),
.B(n_196),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_131),
.B(n_154),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_203),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_213),
.B1(n_176),
.B2(n_189),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_8),
.C(n_7),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_209),
.C(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_192),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_0),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_7),
.C(n_8),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g213 ( 
.A1(n_159),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_183),
.B1(n_160),
.B2(n_162),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_3),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_3),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_217),
.B(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_4),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_190),
.B1(n_191),
.B2(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

XOR2x2_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_164),
.Y(n_226)
);

XOR2x1_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_219),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_201),
.B1(n_196),
.B2(n_206),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_235),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_170),
.C(n_168),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_195),
.C(n_207),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_173),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_200),
.C(n_204),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_242),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_167),
.B1(n_184),
.B2(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_174),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_259),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_258),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_197),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_200),
.B(n_217),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_255),
.A2(n_262),
.B(n_215),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_229),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_212),
.C(n_198),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_231),
.C(n_236),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_243),
.B1(n_214),
.B2(n_238),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_210),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_277),
.C(n_208),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_276),
.B1(n_249),
.B2(n_248),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_216),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_160),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_230),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_243),
.B1(n_234),
.B2(n_239),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_211),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_256),
.C(n_247),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_249),
.B1(n_244),
.B2(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_247),
.C(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_245),
.C(n_244),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_245),
.C(n_237),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_235),
.B(n_242),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_263),
.A2(n_202),
.B1(n_227),
.B2(n_213),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_273),
.B1(n_276),
.B2(n_202),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_272),
.B(n_270),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_294),
.B(n_290),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_266),
.B1(n_264),
.B2(n_222),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_299),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_284),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_230),
.B1(n_199),
.B2(n_232),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_288),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_308),
.B1(n_299),
.B2(n_295),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_287),
.B(n_221),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_301),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_310),
.B(n_303),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_309),
.B1(n_313),
.B2(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_213),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_6),
.C(n_289),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_6),
.Y(n_319)
);


endmodule