module fake_netlist_6_4106_n_1158 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1158);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1158;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_1074;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_1075;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1146;
wire n_1141;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_1107;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_108),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_74),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_101),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_19),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_86),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_75),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_65),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_111),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

BUFx8_ASAP7_75t_SL g236 ( 
.A(n_117),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_105),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_91),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_115),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_116),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_140),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_102),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_164),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_64),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_47),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_152),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_50),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_14),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_56),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_72),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_118),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_109),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_76),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_73),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_77),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_158),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_70),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_125),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_123),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_16),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_0),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_7),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_185),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_120),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_12),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_213),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_28),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_38),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_129),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_221),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_217),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_226),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_240),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_260),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_216),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_236),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_236),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_269),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_257),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_284),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_218),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_219),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_228),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_231),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_232),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_229),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

NAND2xp33_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_232),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_245),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_307),
.A2(n_262),
.B1(n_234),
.B2(n_238),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_325),
.A2(n_283),
.B1(n_280),
.B2(n_276),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_287),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_289),
.A2(n_312),
.B1(n_300),
.B2(n_303),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_323),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_288),
.B(n_231),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_323),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_235),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_306),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_335),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_242),
.Y(n_365)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_243),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_289),
.A2(n_271),
.B1(n_268),
.B2(n_266),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_295),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_296),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_305),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_294),
.Y(n_380)
);

OAI22x1_ASAP7_75t_R g381 ( 
.A1(n_316),
.A2(n_264),
.B1(n_247),
.B2(n_261),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_301),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_239),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_301),
.A2(n_321),
.B(n_320),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_290),
.B(n_292),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_351),
.Y(n_391)
);

NOR2x1p5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_316),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_382),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_326),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_337),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_386),
.B(n_326),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_353),
.Y(n_397)
);

AND3x2_ASAP7_75t_L g398 ( 
.A(n_343),
.B(n_333),
.C(n_291),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_344),
.B(n_328),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_351),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_344),
.A2(n_330),
.B1(n_315),
.B2(n_328),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_344),
.B(n_291),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_378),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_350),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

AO21x2_ASAP7_75t_L g413 ( 
.A1(n_341),
.A2(n_232),
.B(n_315),
.Y(n_413)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_336),
.A2(n_232),
.B(n_250),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_357),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_371),
.B(n_317),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

CKINVDCx11_ASAP7_75t_R g423 ( 
.A(n_347),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_251),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_366),
.B(n_317),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_387),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_387),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_352),
.B(n_293),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_364),
.A2(n_384),
.B1(n_371),
.B2(n_367),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_365),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_365),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_369),
.B(n_299),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_366),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_355),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

NOR2x1p5_ASAP7_75t_L g447 ( 
.A(n_355),
.B(n_252),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_339),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_339),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_337),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_253),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_338),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_337),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_373),
.B(n_299),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_342),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_341),
.B(n_254),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_373),
.B(n_390),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_348),
.B(n_239),
.Y(n_463)
);

AND3x2_ASAP7_75t_L g464 ( 
.A(n_343),
.B(n_263),
.C(n_232),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g465 ( 
.A1(n_362),
.A2(n_258),
.B(n_256),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_411),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_423),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_422),
.B(n_365),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_363),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_397),
.B(n_353),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

XNOR2x2_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_381),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_370),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_412),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_418),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_360),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_430),
.B(n_372),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_418),
.B(n_390),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_391),
.B(n_374),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_401),
.B(n_366),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_405),
.Y(n_486)
);

XNOR2x2_ASAP7_75t_L g487 ( 
.A(n_404),
.B(n_463),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_428),
.B(n_366),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_432),
.B(n_390),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_456),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_432),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_459),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_459),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_411),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_391),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_458),
.B(n_345),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_433),
.B(n_346),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_452),
.B(n_358),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_443),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_403),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_439),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_408),
.B(n_358),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_408),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_403),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_458),
.B(n_361),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_452),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_431),
.A2(n_361),
.B(n_340),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_445),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_446),
.Y(n_520)
);

XNOR2x2_ASAP7_75t_L g521 ( 
.A(n_438),
.B(n_1),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_396),
.B(n_259),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_368),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_449),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_393),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_449),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_417),
.A2(n_340),
.B(n_380),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_394),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_435),
.B(n_368),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_455),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_411),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_419),
.B(n_263),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_419),
.B(n_340),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_413),
.B(n_368),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_455),
.B(n_33),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_425),
.Y(n_540)
);

AND2x2_ASAP7_75t_SL g541 ( 
.A(n_427),
.B(n_368),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_1),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_437),
.B(n_368),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_448),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_439),
.B(n_342),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_420),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_437),
.B(n_354),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_L g552 ( 
.A(n_506),
.B(n_461),
.C(n_414),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_488),
.B(n_439),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_515),
.B(n_413),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_468),
.A2(n_447),
.B1(n_392),
.B2(n_441),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_413),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_513),
.B(n_465),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_514),
.B(n_439),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_513),
.B(n_465),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_469),
.A2(n_465),
.B1(n_399),
.B2(n_402),
.Y(n_560)
);

AND2x4_ASAP7_75t_SL g561 ( 
.A(n_503),
.B(n_509),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_398),
.C(n_464),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_488),
.B(n_406),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_471),
.B(n_436),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_469),
.A2(n_399),
.B1(n_402),
.B2(n_400),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_496),
.B(n_406),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_480),
.B(n_392),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_541),
.A2(n_447),
.B1(n_436),
.B2(n_441),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_476),
.B(n_407),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_472),
.B(n_417),
.Y(n_571)
);

OAI22x1_ASAP7_75t_R g572 ( 
.A1(n_467),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_572)
);

BUFx2_ASAP7_75t_R g573 ( 
.A(n_470),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_491),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_417),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_502),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_477),
.B(n_411),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_429),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

OAI221xp5_ASAP7_75t_L g580 ( 
.A1(n_481),
.A2(n_400),
.B1(n_453),
.B2(n_450),
.C(n_415),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_537),
.A2(n_429),
.B(n_415),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_484),
.B(n_429),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_486),
.B(n_429),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_492),
.B(n_407),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_468),
.A2(n_537),
.B1(n_479),
.B2(n_474),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_504),
.A2(n_483),
.B1(n_533),
.B2(n_485),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_523),
.B(n_416),
.Y(n_587)
);

BUFx4f_ASAP7_75t_SL g588 ( 
.A(n_531),
.Y(n_588)
);

BUFx8_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

AND2x6_ASAP7_75t_SL g590 ( 
.A(n_543),
.B(n_2),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_474),
.A2(n_453),
.B1(n_421),
.B2(n_416),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_517),
.B(n_414),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_497),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_518),
.A2(n_421),
.B(n_454),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_521),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_487),
.B(n_442),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_493),
.A2(n_457),
.B1(n_454),
.B2(n_442),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_494),
.B(n_442),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_482),
.B(n_457),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_495),
.B(n_442),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_498),
.B(n_395),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_512),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_478),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_395),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_528),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_479),
.B(n_395),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_476),
.B(n_395),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_549),
.B(n_34),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_539),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_489),
.B(n_490),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_522),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_480),
.B(n_3),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_519),
.B(n_395),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_489),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_520),
.B(n_424),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_424),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_489),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_574),
.B(n_536),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_614),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_589),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_574),
.B(n_490),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_561),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_585),
.B(n_490),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_567),
.B(n_507),
.Y(n_627)
);

O2A1O1Ixp5_ASAP7_75t_L g628 ( 
.A1(n_555),
.A2(n_529),
.B(n_526),
.C(n_530),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_579),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_597),
.B(n_507),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_619),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_597),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_571),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_562),
.B(n_473),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_605),
.B(n_4),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_594),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_616),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_607),
.Y(n_640)
);

INVx8_ASAP7_75t_L g641 ( 
.A(n_616),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_593),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_586),
.B(n_510),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_596),
.B(n_604),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_613),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_616),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_525),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_575),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_567),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_616),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_R g652 ( 
.A(n_558),
.B(n_538),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_584),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_598),
.B(n_525),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_578),
.B(n_540),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_557),
.B(n_544),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_564),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_R g658 ( 
.A(n_588),
.B(n_542),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_577),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_588),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_SL g661 ( 
.A(n_559),
.B(n_572),
.C(n_566),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_554),
.B(n_601),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_582),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_610),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_603),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_552),
.B(n_510),
.Y(n_667)
);

NOR3xp33_ASAP7_75t_SL g668 ( 
.A(n_590),
.B(n_546),
.C(n_545),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_583),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_608),
.B(n_550),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_600),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_SL g672 ( 
.A(n_553),
.B(n_529),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_552),
.A2(n_532),
.B1(n_527),
.B2(n_547),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_573),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_602),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_615),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_SL g677 ( 
.A(n_563),
.B(n_501),
.C(n_466),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_606),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_617),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_618),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_560),
.B(n_565),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_611),
.B(n_532),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_609),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_580),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_591),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_569),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_595),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_688),
.A2(n_581),
.A3(n_518),
.B(n_551),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_650),
.B(n_570),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_671),
.A2(n_560),
.B(n_534),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_654),
.B(n_592),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_681),
.A2(n_548),
.B(n_599),
.C(n_460),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_662),
.A2(n_460),
.B(n_424),
.Y(n_695)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_667),
.A2(n_460),
.B(n_424),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_632),
.B(n_5),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_671),
.A2(n_628),
.B(n_673),
.Y(n_698)
);

BUFx4f_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_686),
.A2(n_460),
.B1(n_424),
.B2(n_380),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_633),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_671),
.A2(n_460),
.B(n_354),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_632),
.B(n_5),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_6),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_670),
.A2(n_354),
.B(n_36),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_656),
.B(n_653),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_642),
.B(n_6),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_688),
.A2(n_380),
.B(n_342),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_644),
.A2(n_380),
.B(n_342),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_625),
.A2(n_380),
.B(n_354),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_650),
.B(n_35),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_659),
.A2(n_354),
.B(n_40),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_685),
.A2(n_41),
.B(n_37),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_681),
.A2(n_43),
.B(n_42),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_620),
.B(n_8),
.Y(n_715)
);

AO31x2_ASAP7_75t_L g716 ( 
.A1(n_687),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_629),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_643),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_645),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_682),
.B(n_9),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_672),
.A2(n_342),
.B(n_12),
.C(n_13),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_659),
.A2(n_46),
.B(n_45),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_672),
.A2(n_49),
.B(n_48),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_641),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_646),
.Y(n_725)
);

AND3x2_ASAP7_75t_L g726 ( 
.A(n_622),
.B(n_10),
.C(n_13),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_635),
.A2(n_52),
.B(n_51),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_623),
.B(n_14),
.Y(n_728)
);

AO21x1_ASAP7_75t_L g729 ( 
.A1(n_687),
.A2(n_15),
.B(n_16),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_624),
.B(n_15),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_623),
.B(n_17),
.Y(n_731)
);

AOI21xp33_ASAP7_75t_L g732 ( 
.A1(n_621),
.A2(n_17),
.B(n_18),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_640),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_665),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_627),
.B(n_215),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_641),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_648),
.A2(n_54),
.B(n_53),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_634),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_664),
.A2(n_675),
.B(n_649),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_664),
.A2(n_57),
.B(n_55),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_635),
.A2(n_649),
.B(n_657),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_686),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_641),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_675),
.A2(n_657),
.B(n_676),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_634),
.B(n_20),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_636),
.B(n_21),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_669),
.A2(n_130),
.B(n_212),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_684),
.A2(n_128),
.B(n_211),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_663),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_678),
.A2(n_127),
.B(n_208),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_661),
.B(n_21),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_663),
.B(n_22),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_SL g753 ( 
.A1(n_720),
.A2(n_637),
.B1(n_674),
.B2(n_665),
.C(n_680),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_743),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_718),
.Y(n_755)
);

AO31x2_ASAP7_75t_L g756 ( 
.A1(n_694),
.A2(n_684),
.A3(n_679),
.B(n_630),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_734),
.A2(n_627),
.B1(n_660),
.B2(n_624),
.Y(n_757)
);

OA22x2_ASAP7_75t_L g758 ( 
.A1(n_726),
.A2(n_637),
.B1(n_633),
.B2(n_627),
.Y(n_758)
);

OA21x2_ASAP7_75t_L g759 ( 
.A1(n_710),
.A2(n_677),
.B(n_655),
.Y(n_759)
);

AO31x2_ASAP7_75t_L g760 ( 
.A1(n_708),
.A2(n_638),
.A3(n_651),
.B(n_639),
.Y(n_760)
);

AND3x2_ASAP7_75t_L g761 ( 
.A(n_714),
.B(n_660),
.C(n_651),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_714),
.A2(n_683),
.B(n_668),
.C(n_666),
.Y(n_762)
);

AO31x2_ASAP7_75t_L g763 ( 
.A1(n_695),
.A2(n_639),
.A3(n_648),
.B(n_666),
.Y(n_763)
);

OA21x2_ASAP7_75t_L g764 ( 
.A1(n_710),
.A2(n_683),
.B(n_648),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_743),
.Y(n_765)
);

CKINVDCx11_ASAP7_75t_R g766 ( 
.A(n_749),
.Y(n_766)
);

INVx3_ASAP7_75t_SL g767 ( 
.A(n_701),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_741),
.A2(n_666),
.B(n_641),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_713),
.A2(n_666),
.B(n_647),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_713),
.A2(n_666),
.B(n_647),
.C(n_631),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_735),
.A2(n_631),
.B1(n_648),
.B2(n_647),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_738),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_712),
.A2(n_648),
.B(n_652),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_742),
.A2(n_648),
.B1(n_658),
.B2(n_25),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_706),
.A2(n_214),
.B(n_132),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_702),
.A2(n_124),
.B(n_204),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_743),
.B(n_719),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_692),
.A2(n_206),
.B(n_122),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_721),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_705),
.A2(n_696),
.B(n_698),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_737),
.A2(n_133),
.B(n_202),
.Y(n_781)
);

OAI21x1_ASAP7_75t_L g782 ( 
.A1(n_739),
.A2(n_121),
.B(n_201),
.Y(n_782)
);

AO21x1_ASAP7_75t_L g783 ( 
.A1(n_737),
.A2(n_723),
.B(n_715),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_749),
.B(n_58),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_707),
.B(n_23),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_744),
.A2(n_134),
.B(n_200),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_700),
.A2(n_119),
.B(n_199),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_722),
.A2(n_114),
.B(n_197),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_748),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_740),
.A2(n_113),
.B(n_194),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_691),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_709),
.A2(n_112),
.B(n_193),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_693),
.A2(n_203),
.B(n_110),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_746),
.B(n_26),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_725),
.Y(n_796)
);

AO31x2_ASAP7_75t_L g797 ( 
.A1(n_729),
.A2(n_135),
.A3(n_191),
.B(n_190),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_690),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_727),
.A2(n_192),
.B(n_106),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_697),
.B(n_27),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_699),
.Y(n_801)
);

AND3x1_ASAP7_75t_L g802 ( 
.A(n_751),
.B(n_28),
.C(n_29),
.Y(n_802)
);

AO31x2_ASAP7_75t_L g803 ( 
.A1(n_704),
.A2(n_107),
.A3(n_188),
.B(n_187),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_699),
.Y(n_804)
);

NAND3x1_ASAP7_75t_L g805 ( 
.A(n_752),
.B(n_29),
.C(n_30),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_728),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_736),
.B(n_59),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_731),
.Y(n_808)
);

AOI221x1_ASAP7_75t_L g809 ( 
.A1(n_732),
.A2(n_703),
.B1(n_745),
.B2(n_690),
.C(n_735),
.Y(n_809)
);

AO31x2_ASAP7_75t_L g810 ( 
.A1(n_689),
.A2(n_136),
.A3(n_184),
.B(n_183),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_738),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_711),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_812)
);

CKINVDCx11_ASAP7_75t_R g813 ( 
.A(n_711),
.Y(n_813)
);

NAND2x1p5_ASAP7_75t_L g814 ( 
.A(n_736),
.B(n_60),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_733),
.B(n_189),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_747),
.A2(n_61),
.B(n_62),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_724),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_SL g818 ( 
.A1(n_724),
.A2(n_63),
.B(n_66),
.C(n_67),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_730),
.B(n_68),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_750),
.A2(n_69),
.B(n_71),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_758),
.A2(n_716),
.B1(n_689),
.B2(n_80),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_791),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_783),
.A2(n_716),
.B1(n_79),
.B2(n_81),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_806),
.B(n_716),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_794),
.B(n_785),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_801),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_812),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_755),
.Y(n_829)
);

BUFx4f_ASAP7_75t_SL g830 ( 
.A(n_801),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_774),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_774),
.A2(n_819),
.B1(n_781),
.B2(n_808),
.Y(n_832)
);

BUFx8_ASAP7_75t_SL g833 ( 
.A(n_804),
.Y(n_833)
);

BUFx10_ASAP7_75t_L g834 ( 
.A(n_784),
.Y(n_834)
);

BUFx8_ASAP7_75t_L g835 ( 
.A(n_772),
.Y(n_835)
);

AND2x4_ASAP7_75t_SL g836 ( 
.A(n_765),
.B(n_88),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_802),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_837)
);

INVx6_ASAP7_75t_L g838 ( 
.A(n_813),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_795),
.Y(n_839)
);

CKINVDCx11_ASAP7_75t_R g840 ( 
.A(n_766),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_767),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_SL g842 ( 
.A1(n_800),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_796),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_811),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_798),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_761),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_809),
.B(n_99),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_757),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_817),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_753),
.B(n_100),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_756),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_754),
.Y(n_852)
);

INVx6_ASAP7_75t_L g853 ( 
.A(n_777),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_756),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_793),
.A2(n_103),
.B1(n_137),
.B2(n_138),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_815),
.A2(n_775),
.B1(n_771),
.B2(n_799),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_809),
.B(n_139),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_762),
.B(n_141),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_760),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_769),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_760),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_807),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_760),
.Y(n_863)
);

CKINVDCx6p67_ASAP7_75t_R g864 ( 
.A(n_805),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_SL g865 ( 
.A1(n_787),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_865)
);

BUFx4f_ASAP7_75t_SL g866 ( 
.A(n_814),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_810),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_759),
.B(n_149),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_759),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_768),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_778),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_871)
);

BUFx8_ASAP7_75t_L g872 ( 
.A(n_779),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_763),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_770),
.A2(n_162),
.B1(n_165),
.B2(n_167),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_764),
.Y(n_875)
);

OAI22xp33_ASAP7_75t_L g876 ( 
.A1(n_820),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_764),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_773),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_763),
.B(n_179),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_782),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_780),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_803),
.B(n_181),
.Y(n_883)
);

CKINVDCx6p67_ASAP7_75t_R g884 ( 
.A(n_803),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_797),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_872),
.A2(n_786),
.B1(n_790),
.B2(n_788),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_851),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_873),
.Y(n_888)
);

BUFx2_ASAP7_75t_SL g889 ( 
.A(n_841),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_854),
.Y(n_890)
);

BUFx2_ASAP7_75t_SL g891 ( 
.A(n_858),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_859),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_873),
.A2(n_816),
.B(n_792),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_822),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_881),
.A2(n_816),
.B(n_792),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_861),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_823),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_844),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_839),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_825),
.B(n_797),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_845),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_843),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_825),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_875),
.B(n_786),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_872),
.A2(n_776),
.B1(n_789),
.B2(n_818),
.Y(n_905)
);

INVx4_ASAP7_75t_SL g906 ( 
.A(n_858),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_875),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_882),
.A2(n_182),
.B(n_867),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_878),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_863),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_885),
.Y(n_911)
);

AO21x2_ASAP7_75t_L g912 ( 
.A1(n_847),
.A2(n_857),
.B(n_880),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_829),
.B(n_884),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_849),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_835),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_880),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_868),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_868),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_883),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_826),
.B(n_857),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_847),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_821),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_824),
.A2(n_856),
.B(n_874),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_853),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_832),
.B(n_834),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_874),
.A2(n_877),
.B(n_879),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_835),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_853),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_834),
.B(n_850),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_853),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_828),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_862),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_828),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_876),
.A2(n_837),
.B(n_869),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_838),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_837),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_852),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_864),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_899),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_887),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_929),
.A2(n_925),
.B(n_900),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_899),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_904),
.B(n_831),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_899),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_907),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_904),
.B(n_846),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_907),
.B(n_860),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_897),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_887),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_887),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_920),
.B(n_838),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_897),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_907),
.B(n_870),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_890),
.Y(n_954)
);

OA21x2_ASAP7_75t_L g955 ( 
.A1(n_893),
.A2(n_871),
.B(n_848),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_894),
.B(n_827),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_890),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_894),
.B(n_827),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_890),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_935),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_893),
.A2(n_855),
.B(n_865),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_903),
.B(n_842),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_902),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_910),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_902),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_902),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_892),
.B(n_838),
.Y(n_967)
);

AO21x2_ASAP7_75t_L g968 ( 
.A1(n_893),
.A2(n_866),
.B(n_833),
.Y(n_968)
);

AOI221xp5_ASAP7_75t_L g969 ( 
.A1(n_922),
.A2(n_830),
.B1(n_836),
.B2(n_840),
.C(n_936),
.Y(n_969)
);

OA21x2_ASAP7_75t_L g970 ( 
.A1(n_895),
.A2(n_908),
.B(n_896),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_895),
.A2(n_911),
.B(n_909),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_903),
.B(n_900),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_909),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_967),
.B(n_945),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_967),
.B(n_945),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_972),
.B(n_912),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_967),
.B(n_888),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_972),
.B(n_912),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_965),
.B(n_888),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_965),
.B(n_920),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_939),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_940),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_940),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_965),
.B(n_912),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_940),
.Y(n_985)
);

AND2x4_ASAP7_75t_SL g986 ( 
.A(n_964),
.B(n_930),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_964),
.B(n_912),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_943),
.A2(n_922),
.B1(n_925),
.B2(n_936),
.C(n_931),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_963),
.B(n_916),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_940),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_939),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_942),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_963),
.B(n_916),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_942),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_956),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_966),
.B(n_919),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_960),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_968),
.B(n_913),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_944),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_974),
.B(n_968),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_974),
.B(n_968),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_981),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_981),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_980),
.B(n_901),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_980),
.B(n_995),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_983),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_983),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_991),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_975),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_975),
.B(n_968),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_991),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_998),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_994),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_987),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_977),
.B(n_941),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_998),
.B(n_960),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1008),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_1012),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_1009),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1006),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1016),
.B(n_998),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1016),
.B(n_997),
.Y(n_1022)
);

INVxp33_ASAP7_75t_L g1023 ( 
.A(n_1016),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1008),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1002),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1003),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_R g1027 ( 
.A(n_1012),
.B(n_938),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1011),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1000),
.B(n_997),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1013),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1022),
.B(n_1021),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1019),
.B(n_1015),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1029),
.B(n_1015),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_1005),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1029),
.B(n_1022),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_1023),
.A2(n_988),
.B(n_929),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1021),
.B(n_1000),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_1026),
.B(n_1004),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1018),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1023),
.B(n_1001),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1036),
.A2(n_1027),
.B1(n_1001),
.B2(n_1010),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_1039),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1040),
.B(n_1010),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_1036),
.B(n_1018),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1035),
.A2(n_891),
.B1(n_969),
.B2(n_935),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1034),
.B(n_1028),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1032),
.A2(n_891),
.B1(n_1030),
.B2(n_938),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_1043),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1045),
.A2(n_1033),
.B(n_1038),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_1041),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1047),
.Y(n_1052)
);

NAND2x1p5_ASAP7_75t_L g1053 ( 
.A(n_1048),
.B(n_935),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1042),
.B(n_1037),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1044),
.B(n_1017),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1046),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1043),
.B(n_1024),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1049),
.B(n_1020),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_SL g1060 ( 
.A(n_1050),
.B(n_969),
.C(n_951),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1051),
.B(n_1020),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1050),
.A2(n_927),
.B1(n_928),
.B2(n_934),
.Y(n_1063)
);

AOI31xp33_ASAP7_75t_L g1064 ( 
.A1(n_1056),
.A2(n_927),
.A3(n_915),
.B(n_928),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_1052),
.B(n_889),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1057),
.B(n_987),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1054),
.A2(n_934),
.B1(n_889),
.B2(n_924),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1065),
.A2(n_1053),
.B1(n_1055),
.B2(n_924),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1061),
.B(n_1014),
.Y(n_1069)
);

OAI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1063),
.A2(n_960),
.B1(n_930),
.B2(n_958),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1059),
.Y(n_1071)
);

AOI22x1_ASAP7_75t_L g1072 ( 
.A1(n_1064),
.A2(n_930),
.B1(n_937),
.B2(n_958),
.Y(n_1072)
);

OAI33xp33_ASAP7_75t_L g1073 ( 
.A1(n_1062),
.A2(n_976),
.A3(n_978),
.B1(n_956),
.B2(n_993),
.B3(n_962),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1067),
.B(n_941),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_1066),
.A2(n_937),
.B(n_932),
.C(n_924),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1069),
.A2(n_1060),
.B(n_905),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1071),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1068),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1070),
.A2(n_930),
.B1(n_934),
.B2(n_932),
.Y(n_1079)
);

AOI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1074),
.A2(n_923),
.B(n_933),
.C(n_931),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1078),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1077),
.B(n_1076),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1079),
.Y(n_1083)
);

CKINVDCx16_ASAP7_75t_R g1084 ( 
.A(n_1080),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1077),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1078),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_L g1087 ( 
.A(n_1081),
.B(n_1072),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_1085),
.B(n_1075),
.C(n_1073),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1086),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1084),
.A2(n_986),
.B1(n_937),
.B2(n_932),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1082),
.B(n_1083),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1082),
.A2(n_1007),
.B(n_1006),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_1091),
.B(n_962),
.C(n_921),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_1089),
.B(n_1007),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_SL g1095 ( 
.A(n_1088),
.B(n_917),
.C(n_921),
.Y(n_1095)
);

OAI221xp5_ASAP7_75t_L g1096 ( 
.A1(n_1087),
.A2(n_917),
.B1(n_976),
.B2(n_978),
.C(n_933),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_1090),
.B(n_901),
.C(n_886),
.Y(n_1097)
);

OAI211xp5_ASAP7_75t_L g1098 ( 
.A1(n_1094),
.A2(n_1092),
.B(n_984),
.C(n_955),
.Y(n_1098)
);

NOR4xp25_ASAP7_75t_L g1099 ( 
.A(n_1096),
.B(n_999),
.C(n_994),
.D(n_984),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_961),
.C(n_908),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1095),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_986),
.B1(n_982),
.B2(n_992),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_L g1103 ( 
.A(n_1096),
.B(n_961),
.C(n_908),
.Y(n_1103)
);

NOR4xp25_ASAP7_75t_L g1104 ( 
.A(n_1096),
.B(n_999),
.C(n_982),
.D(n_979),
.Y(n_1104)
);

OAI211xp5_ASAP7_75t_L g1105 ( 
.A1(n_1094),
.A2(n_955),
.B(n_979),
.C(n_977),
.Y(n_1105)
);

NOR2xp67_ASAP7_75t_L g1106 ( 
.A(n_1098),
.B(n_1105),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1101),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1104),
.B(n_993),
.Y(n_1108)
);

OAI311xp33_ASAP7_75t_L g1109 ( 
.A1(n_1099),
.A2(n_946),
.A3(n_943),
.B1(n_913),
.C1(n_953),
.Y(n_1109)
);

AND3x2_ASAP7_75t_L g1110 ( 
.A(n_1100),
.B(n_898),
.C(n_946),
.Y(n_1110)
);

OAI321xp33_ASAP7_75t_L g1111 ( 
.A1(n_1102),
.A2(n_946),
.A3(n_943),
.B1(n_918),
.B2(n_953),
.C(n_948),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1103),
.Y(n_1112)
);

NAND3x1_ASAP7_75t_SL g1113 ( 
.A(n_1101),
.B(n_953),
.C(n_947),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1101),
.B(n_982),
.Y(n_1114)
);

NAND4xp75_ASAP7_75t_L g1115 ( 
.A(n_1114),
.B(n_955),
.C(n_989),
.D(n_947),
.Y(n_1115)
);

AND3x4_ASAP7_75t_L g1116 ( 
.A(n_1106),
.B(n_918),
.C(n_919),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1107),
.A2(n_934),
.B(n_923),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1113),
.Y(n_1118)
);

OAI21xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1108),
.A2(n_923),
.B(n_926),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1112),
.B(n_996),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_1110),
.B(n_1109),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1111),
.B(n_996),
.Y(n_1122)
);

NOR3x1_ASAP7_75t_L g1123 ( 
.A(n_1108),
.B(n_961),
.C(n_926),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1107),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1107),
.B(n_989),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1107),
.A2(n_926),
.B(n_918),
.Y(n_1126)
);

OR4x1_ASAP7_75t_L g1127 ( 
.A(n_1113),
.B(n_952),
.C(n_948),
.D(n_973),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1124),
.A2(n_990),
.B1(n_985),
.B2(n_919),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_SL g1129 ( 
.A1(n_1118),
.A2(n_955),
.B1(n_990),
.B2(n_985),
.Y(n_1129)
);

AOI31xp33_ASAP7_75t_L g1130 ( 
.A1(n_1121),
.A2(n_947),
.A3(n_952),
.B(n_906),
.Y(n_1130)
);

OAI221xp5_ASAP7_75t_L g1131 ( 
.A1(n_1125),
.A2(n_955),
.B1(n_914),
.B2(n_966),
.C(n_973),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1116),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1120),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1122),
.B(n_906),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1115),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1117),
.B(n_906),
.C(n_914),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1133),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1130),
.Y(n_1138)
);

NAND4xp25_ASAP7_75t_L g1139 ( 
.A(n_1134),
.B(n_1123),
.C(n_1126),
.D(n_1127),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1132),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1135),
.A2(n_1119),
.B1(n_911),
.B2(n_944),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1135),
.A2(n_914),
.B1(n_959),
.B2(n_957),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1137),
.A2(n_1136),
.B1(n_1129),
.B2(n_1128),
.Y(n_1143)
);

OAI22x1_ASAP7_75t_L g1144 ( 
.A1(n_1138),
.A2(n_1131),
.B1(n_970),
.B2(n_959),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1140),
.A2(n_959),
.B1(n_954),
.B2(n_957),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1143),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1146),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1147),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1148),
.A2(n_1141),
.B1(n_1142),
.B2(n_1139),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1148),
.A2(n_1144),
.B1(n_1145),
.B2(n_906),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1148),
.A2(n_970),
.B1(n_971),
.B2(n_906),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1150),
.B(n_970),
.Y(n_1152)
);

XNOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1149),
.B(n_970),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1151),
.B(n_971),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1152),
.B(n_954),
.Y(n_1155)
);

XNOR2x1_ASAP7_75t_L g1156 ( 
.A(n_1153),
.B(n_970),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_1154),
.B(n_959),
.C(n_954),
.Y(n_1157)
);

AOI211xp5_ASAP7_75t_L g1158 ( 
.A1(n_1157),
.A2(n_1155),
.B(n_950),
.C(n_949),
.Y(n_1158)
);


endmodule