module fake_jpeg_15204_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_0),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_1),
.B(n_2),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_17),
.B1(n_34),
.B2(n_33),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_40),
.C(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_8),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_59),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_1),
.B(n_4),
.Y(n_72)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_4),
.Y(n_74)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_42),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_21),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_45),
.A3(n_42),
.B1(n_36),
.B2(n_23),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_78),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_46),
.B(n_15),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_73),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_9),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_9),
.Y(n_91)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_64),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_89),
.B1(n_77),
.B2(n_78),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_99),
.B1(n_84),
.B2(n_86),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_11),
.B(n_12),
.C(n_14),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_87),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_90),
.B1(n_99),
.B2(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_25),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_26),
.C(n_28),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_29),
.B(n_35),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_94),
.Y(n_112)
);


endmodule