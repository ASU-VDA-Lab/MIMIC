module fake_jpeg_1191_n_172 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_0),
.B(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_41),
.Y(n_84)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_36),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_40),
.Y(n_94)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_69),
.B1(n_16),
.B2(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_53),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_37),
.B1(n_51),
.B2(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_4),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_61),
.Y(n_88)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_66),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_56),
.Y(n_93)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_58),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_19),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_71),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_32),
.A2(n_11),
.B(n_9),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_24),
.B(n_10),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_72),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_18),
.A2(n_16),
.B1(n_24),
.B2(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_41),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_96),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_11),
.B1(n_58),
.B2(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_38),
.A2(n_45),
.B1(n_65),
.B2(n_59),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_36),
.C(n_49),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_94),
.C(n_84),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_42),
.B1(n_37),
.B2(n_61),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_34),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_34),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_95),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_124),
.C(n_84),
.Y(n_126)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_79),
.B1(n_85),
.B2(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_118),
.Y(n_128)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_121),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_122),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_75),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_87),
.C(n_94),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_132),
.C(n_117),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_86),
.B(n_93),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_102),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_98),
.B(n_83),
.C(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_107),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_124),
.C(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_126),
.C(n_137),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_112),
.B1(n_110),
.B2(n_113),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_147),
.B(n_136),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_110),
.B1(n_123),
.B2(n_114),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_130),
.B(n_138),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_123),
.B(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_162),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_147),
.B1(n_153),
.B2(n_144),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_131),
.C(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_158),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_167),
.B1(n_165),
.B2(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_150),
.B(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_109),
.C(n_97),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_92),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_171),
.Y(n_172)
);


endmodule