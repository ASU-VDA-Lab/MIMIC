module fake_jpeg_31081_n_405 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_405);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_0),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_20),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_45),
.Y(n_83)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_40),
.B1(n_48),
.B2(n_45),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_118),
.B1(n_120),
.B2(n_38),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_93),
.Y(n_158)
);

CKINVDCx11_ASAP7_75t_R g100 ( 
.A(n_55),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_116),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_61),
.A2(n_40),
.B1(n_48),
.B2(n_45),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_64),
.A2(n_40),
.B1(n_48),
.B2(n_32),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_84),
.B1(n_82),
.B2(n_78),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_121),
.B1(n_114),
.B2(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_155),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_131),
.B(n_140),
.Y(n_178)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_80),
.B1(n_51),
.B2(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_138),
.B1(n_152),
.B2(n_92),
.Y(n_166)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_77),
.B1(n_72),
.B2(n_66),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_94),
.B(n_73),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_76),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_67),
.B1(n_58),
.B2(n_53),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_154),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_32),
.B1(n_56),
.B2(n_70),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_26),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_23),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_97),
.B(n_36),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_21),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_172),
.B1(n_175),
.B2(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_121),
.B1(n_114),
.B2(n_103),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_104),
.B1(n_119),
.B2(n_111),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_130),
.A2(n_118),
.B1(n_123),
.B2(n_102),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_24),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_30),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_195),
.Y(n_212)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_188),
.Y(n_228)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_131),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_198),
.Y(n_214)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_155),
.B(n_149),
.C(n_154),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_154),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_147),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_205),
.Y(n_217)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_149),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_157),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_149),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_22),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_22),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_164),
.B1(n_172),
.B2(n_163),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_213),
.B1(n_216),
.B2(n_220),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_195),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_164),
.B1(n_166),
.B2(n_111),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_186),
.C(n_181),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_227),
.C(n_71),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_196),
.B1(n_199),
.B2(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_219),
.B(n_207),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_161),
.B1(n_162),
.B2(n_119),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_229),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_173),
.B(n_156),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_225),
.B(n_167),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_156),
.B(n_162),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_160),
.C(n_173),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_68),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_190),
.B1(n_189),
.B2(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_243),
.B1(n_249),
.B2(n_158),
.Y(n_273)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_233),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_216),
.A2(n_190),
.B(n_188),
.C(n_192),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_252),
.B(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_192),
.B1(n_191),
.B2(n_189),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_246),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_241),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_191),
.B1(n_182),
.B2(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_248),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_170),
.B1(n_202),
.B2(n_177),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_170),
.B1(n_176),
.B2(n_174),
.Y(n_244)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_176),
.B1(n_177),
.B2(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_210),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_150),
.B1(n_151),
.B2(n_139),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_193),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_167),
.B(n_146),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_23),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_223),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_259),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_256),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_234),
.B(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_269),
.C(n_271),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_222),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_237),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_223),
.C(n_218),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_218),
.C(n_132),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_SL g272 ( 
.A1(n_234),
.A2(n_136),
.B(n_153),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_127),
.B1(n_153),
.B2(n_146),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_280),
.B1(n_254),
.B2(n_127),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_35),
.B(n_188),
.C(n_158),
.D(n_36),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_230),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_231),
.A2(n_137),
.B1(n_145),
.B2(n_110),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_238),
.C(n_239),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_237),
.C(n_249),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_242),
.B(n_46),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_46),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_16),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_264),
.A2(n_234),
.B1(n_240),
.B2(n_245),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_290),
.B1(n_298),
.B2(n_261),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_271),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_234),
.B1(n_244),
.B2(n_237),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_292),
.B(n_145),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_302),
.Y(n_309)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_243),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_251),
.C(n_235),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_304),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_297),
.B(n_305),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_255),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_268),
.B1(n_283),
.B2(n_279),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_30),
.B1(n_24),
.B2(n_42),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_39),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_117),
.C(n_135),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_269),
.B(n_19),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_258),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_262),
.B1(n_268),
.B2(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_311),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_314),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_293),
.B1(n_307),
.B2(n_292),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_322),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_289),
.A2(n_277),
.B1(n_278),
.B2(n_283),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_10),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_241),
.B1(n_110),
.B2(n_42),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_326),
.B(n_62),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_329),
.A2(n_13),
.B(n_20),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_286),
.C(n_296),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_331),
.C(n_339),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_286),
.C(n_304),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_309),
.A2(n_285),
.B(n_284),
.C(n_49),
.Y(n_333)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

OAI321xp33_ASAP7_75t_L g335 ( 
.A1(n_309),
.A2(n_284),
.A3(n_18),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_335)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_337),
.B(n_308),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_83),
.C(n_47),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_340),
.B(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_42),
.C(n_47),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_343),
.C(n_317),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_47),
.C(n_95),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_91),
.C(n_87),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_346),
.B(n_329),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_115),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_319),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_348),
.B(n_355),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_315),
.Y(n_349)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_328),
.Y(n_350)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_338),
.A2(n_314),
.B(n_324),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_358),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_359),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_325),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_338),
.A2(n_323),
.B1(n_310),
.B2(n_321),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_356),
.B1(n_351),
.B2(n_361),
.Y(n_371)
);

OA22x2_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_322),
.B1(n_323),
.B2(n_115),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_341),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_366),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_333),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_330),
.C(n_331),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_369),
.C(n_372),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_339),
.B(n_343),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_354),
.B(n_332),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_336),
.C(n_337),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_9),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_332),
.C(n_91),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_363),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_375),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_353),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_376),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_380),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_9),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_8),
.Y(n_385)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_373),
.A2(n_10),
.B(n_20),
.Y(n_382)
);

AOI31xp67_ASAP7_75t_L g391 ( 
.A1(n_382),
.A2(n_8),
.A3(n_18),
.B(n_4),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_369),
.B1(n_365),
.B2(n_98),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_383),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_365),
.A2(n_7),
.B(n_18),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_384),
.A2(n_5),
.B(n_6),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_392),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_377),
.A2(n_93),
.B1(n_87),
.B2(n_3),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

O2A1O1Ixp33_ASAP7_75t_SL g396 ( 
.A1(n_391),
.A2(n_12),
.B(n_14),
.C(n_1),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_378),
.B(n_379),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_393),
.A2(n_390),
.B(n_388),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g394 ( 
.A(n_387),
.B(n_378),
.CI(n_5),
.CON(n_394),
.SN(n_394)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_12),
.C(n_14),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_396),
.B(n_385),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_398),
.A2(n_399),
.B(n_400),
.C(n_397),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_395),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_402),
.A2(n_93),
.B(n_1),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_403),
.A2(n_1),
.B(n_2),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_2),
.C(n_231),
.Y(n_405)
);


endmodule