module fake_jpeg_10558_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.C(n_26),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_22),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_17),
.B1(n_28),
.B2(n_20),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_50),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_21),
.B1(n_27),
.B2(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_63),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_34),
.B1(n_21),
.B2(n_27),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_83),
.B1(n_92),
.B2(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_34),
.B1(n_51),
.B2(n_20),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_98),
.B1(n_32),
.B2(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_84),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_52),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_97),
.B1(n_62),
.B2(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_38),
.B1(n_37),
.B2(n_26),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_31),
.B1(n_33),
.B2(n_23),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_106),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_58),
.B1(n_59),
.B2(n_48),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_98),
.B1(n_87),
.B2(n_80),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_87),
.CI(n_75),
.CON(n_106),
.SN(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_116),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_62),
.A3(n_60),
.B1(n_42),
.B2(n_41),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_121),
.B(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_19),
.B1(n_73),
.B2(n_91),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_19),
.B(n_42),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_87),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_47),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_145),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_131),
.B1(n_144),
.B2(n_68),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_80),
.B1(n_90),
.B2(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_96),
.B1(n_85),
.B2(n_90),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_154),
.B1(n_100),
.B2(n_112),
.Y(n_169)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_84),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_140),
.B(n_99),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_1),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_90),
.B1(n_78),
.B2(n_95),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_50),
.B1(n_67),
.B2(n_23),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_150),
.B1(n_111),
.B2(n_116),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_104),
.B1(n_121),
.B2(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_155),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_110),
.A2(n_73),
.B1(n_97),
.B2(n_33),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_100),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_160),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_168),
.C(n_172),
.Y(n_192)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_113),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_33),
.B1(n_31),
.B2(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_176),
.B(n_178),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_114),
.B(n_115),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_184),
.B(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_109),
.C(n_102),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_106),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_175),
.B(n_10),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_130),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_73),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_132),
.A2(n_102),
.B1(n_106),
.B2(n_55),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_138),
.B1(n_139),
.B2(n_133),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_57),
.B(n_18),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_165),
.Y(n_216)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_207),
.B1(n_214),
.B2(n_176),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_140),
.C(n_138),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_216),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_139),
.B(n_146),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_178),
.B(n_171),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_146),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_140),
.C(n_18),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_174),
.C(n_166),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_202),
.A2(n_186),
.B(n_177),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_18),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_33),
.B1(n_31),
.B2(n_24),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_31),
.B1(n_24),
.B2(n_1),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_163),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_175),
.C(n_180),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_228),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_196),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_161),
.A3(n_171),
.B1(n_187),
.B2(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_227),
.B(n_231),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_171),
.B(n_161),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_159),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_158),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_184),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_232),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_157),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_238),
.B1(n_241),
.B2(n_208),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_191),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_157),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_1),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_214),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_190),
.B1(n_194),
.B2(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_192),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_261),
.C(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_216),
.B1(n_210),
.B2(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_239),
.B1(n_219),
.B2(n_217),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_262),
.B1(n_242),
.B2(n_221),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_226),
.A2(n_188),
.B1(n_199),
.B2(n_177),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_220),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_200),
.C(n_204),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_228),
.C(n_232),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_164),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_24),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_223),
.Y(n_265)
);

OAI211xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_244),
.B(n_259),
.C(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_276),
.C(n_277),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_229),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_269),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_225),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_241),
.C(n_229),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_234),
.C(n_24),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_24),
.C(n_2),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_252),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_9),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_255),
.B(n_264),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_291),
.B(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_258),
.B1(n_251),
.B2(n_245),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_305)
);

XOR2x2_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_243),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_267),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_8),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_268),
.A2(n_254),
.B(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_247),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_299),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_270),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_301),
.B(n_306),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_298),
.A2(n_303),
.B(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_250),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_277),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_9),
.B(n_3),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_11),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_12),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_5),
.A3(n_6),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_SL g307 ( 
.A(n_298),
.B(n_283),
.C(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_289),
.B1(n_291),
.B2(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_314),
.Y(n_320)
);

AO221x1_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_289),
.B1(n_290),
.B2(n_281),
.C(n_7),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_312),
.A2(n_16),
.B(n_2),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_6),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_319),
.B(n_321),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_13),
.Y(n_317)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_315),
.B(n_309),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_322),
.B(n_310),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_320),
.B(n_16),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_323),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_2),
.Y(n_329)
);


endmodule