module fake_jpeg_12649_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_15),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_0),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_3),
.B(n_4),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_80),
.Y(n_88)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_5),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_6),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_78),
.A2(n_70),
.B1(n_50),
.B2(n_69),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_86),
.B(n_89),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_58),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_10),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_69),
.B1(n_62),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_69),
.B1(n_66),
.B2(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_68),
.B1(n_61),
.B2(n_52),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_6),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_68),
.B1(n_61),
.B2(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_71),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_56),
.B1(n_55),
.B2(n_53),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_56),
.B1(n_54),
.B2(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_72),
.B1(n_55),
.B2(n_54),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_57),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_25),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_17),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_8),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_9),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_29),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_83),
.B(n_12),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_125),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_127),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_31),
.B(n_47),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_24),
.B(n_36),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_28),
.B(n_46),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_38),
.B(n_41),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_11),
.C(n_12),
.Y(n_125)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_32),
.C(n_45),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_132),
.C(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_42),
.B1(n_48),
.B2(n_119),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_34),
.C(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_13),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_136),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_17),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_145),
.C(n_146),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_97),
.B1(n_118),
.B2(n_110),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_148),
.B(n_145),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_35),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_144),
.B1(n_149),
.B2(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_120),
.B1(n_133),
.B2(n_122),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_22),
.C(n_23),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_124),
.C(n_129),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_157),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_126),
.B(n_130),
.C(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_160),
.B1(n_151),
.B2(n_155),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_141),
.B(n_137),
.C(n_140),
.D(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_164),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_156),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_159),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_166),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_161),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_161),
.B(n_154),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_158),
.Y(n_171)
);


endmodule