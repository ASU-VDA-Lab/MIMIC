module fake_jpeg_930_n_220 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_220);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_46),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_23),
.A2(n_6),
.B(n_1),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_54),
.B(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_23),
.A2(n_8),
.B(n_1),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_31),
.B1(n_13),
.B2(n_29),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_88),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_65),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_31),
.C(n_30),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_11),
.C(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_36),
.A2(n_13),
.B1(n_27),
.B2(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_84),
.B1(n_85),
.B2(n_61),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_32),
.B(n_29),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_89),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_40),
.A2(n_24),
.B1(n_2),
.B2(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_11),
.B1(n_12),
.B2(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_24),
.B1(n_0),
.B2(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_2),
.B1(n_5),
.B2(n_8),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_9),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_62),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_43),
.B1(n_50),
.B2(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_41),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_41),
.CON(n_102),
.SN(n_102)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_105),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_11),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_116),
.C(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_59),
.B1(n_55),
.B2(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_112),
.B1(n_116),
.B2(n_94),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_109),
.B(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_55),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_71),
.B1(n_76),
.B2(n_78),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_57),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_90),
.C(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_74),
.A3(n_56),
.B1(n_58),
.B2(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_123),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_91),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_71),
.B1(n_92),
.B2(n_60),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_134),
.B1(n_140),
.B2(n_133),
.Y(n_156)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_136),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_106),
.B(n_102),
.C(n_99),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_135),
.B(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_139),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_96),
.B1(n_104),
.B2(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_144),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_97),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_121),
.B(n_122),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_111),
.C(n_101),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_155),
.C(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_100),
.B1(n_101),
.B2(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_142),
.B1(n_139),
.B2(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_162),
.B1(n_137),
.B2(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_133),
.B1(n_123),
.B2(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_134),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.C(n_162),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_150),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_124),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_153),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_138),
.B(n_137),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_146),
.B1(n_154),
.B2(n_157),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_156),
.B1(n_146),
.B2(n_161),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_187),
.B1(n_170),
.B2(n_167),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_189),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_148),
.B1(n_147),
.B2(n_158),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_158),
.C(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_168),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_177),
.C(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_195),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_166),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_182),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.C(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_182),
.C(n_187),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_181),
.B(n_185),
.Y(n_205)
);

OAI31xp33_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_181),
.A3(n_198),
.B(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_204),
.B(n_192),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_206),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_218),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_216),
.Y(n_220)
);


endmodule