module fake_ariane_3311_n_3280 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_844, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_3280);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_3280;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3063;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2663;
wire n_2233;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_3207;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_3003;
wire n_2874;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_3126;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3119;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1468;
wire n_1253;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2930;
wire n_2871;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_1623;
wire n_990;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_3052;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3179;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_3260;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_1708;
wire n_3085;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_1373;
wire n_1975;
wire n_1081;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3097;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2723;
wire n_2928;
wire n_1118;
wire n_943;
wire n_2905;
wire n_2884;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_961;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_3107;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2890;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_3184;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2796;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_2647;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_2935;
wire n_2401;
wire n_889;
wire n_3255;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_3243;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_1968;
wire n_918;
wire n_1885;
wire n_3251;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3241;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_3106;
wire n_2977;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3269;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3248;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_3091;
wire n_1024;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_898;
wire n_857;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3111;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_3146;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_3143;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_3196;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_2052;
wire n_1091;
wire n_2485;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2275;
wire n_2205;
wire n_2183;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_1474;
wire n_937;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_2573;
wire n_2940;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx2_ASAP7_75t_SL g845 ( 
.A(n_737),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_216),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_135),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_453),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_663),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_831),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_685),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_586),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_722),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_561),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_354),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_689),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_757),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_752),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_533),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_378),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_326),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_800),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_803),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_781),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_690),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_802),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_150),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_822),
.Y(n_868)
);

BUFx2_ASAP7_75t_SL g869 ( 
.A(n_431),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_603),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_680),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_306),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_707),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_693),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_605),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_513),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_351),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_475),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_710),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_103),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_735),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_279),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_323),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_202),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_482),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_843),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_804),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_216),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_145),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_62),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_264),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_233),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_794),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_713),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_450),
.Y(n_895)
);

BUFx10_ASAP7_75t_L g896 ( 
.A(n_696),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_695),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_294),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_799),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_747),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_708),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_347),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_753),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_359),
.Y(n_904)
);

CKINVDCx14_ASAP7_75t_R g905 ( 
.A(n_675),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_725),
.Y(n_906)
);

CKINVDCx16_ASAP7_75t_R g907 ( 
.A(n_805),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_811),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_821),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_523),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_582),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_571),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_499),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_748),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_14),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_681),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_32),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_762),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_389),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_232),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_705),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_808),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_827),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_739),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_578),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_46),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_62),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_785),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_796),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_186),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_809),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_699),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_510),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_755),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_300),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_203),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_730),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_333),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_203),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_241),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_678),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_773),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_742),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_149),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_97),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_780),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_238),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_311),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_296),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_517),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_836),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_823),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_638),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_209),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_63),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_229),
.Y(n_956)
);

CKINVDCx14_ASAP7_75t_R g957 ( 
.A(n_492),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_782),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_740),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_691),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_338),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_383),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_127),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_682),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_656),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_824),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_826),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_278),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_686),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_606),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_194),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_784),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_763),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_697),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_400),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_348),
.Y(n_976)
);

BUFx10_ASAP7_75t_L g977 ( 
.A(n_118),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_834),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_779),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_50),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_724),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_790),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_674),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_819),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_716),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_698),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_404),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_246),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_621),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_635),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_734),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_720),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_502),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_761),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_840),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_759),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_266),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_495),
.Y(n_998)
);

CKINVDCx16_ASAP7_75t_R g999 ( 
.A(n_727),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_770),
.Y(n_1000)
);

BUFx5_ASAP7_75t_L g1001 ( 
.A(n_797),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_835),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_688),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_294),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_267),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_837),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_327),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_583),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_365),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_50),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_556),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_618),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_668),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_462),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_832),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_130),
.Y(n_1016)
);

BUFx10_ASAP7_75t_L g1017 ( 
.A(n_741),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_376),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_442),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_812),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_158),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_666),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_738),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_354),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_552),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_590),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_193),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_694),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_700),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_486),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_501),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_454),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_191),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_111),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_772),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_99),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_324),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_160),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_473),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_732),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_174),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_719),
.Y(n_1042)
);

INVxp67_ASAP7_75t_SL g1043 ( 
.A(n_665),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_650),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_342),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_426),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_112),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_745),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_795),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_478),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_706),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_65),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_428),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_71),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_711),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_801),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_768),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_448),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_828),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_70),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_170),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_153),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_193),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_212),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_149),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_810),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_673),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_701),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_756),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_628),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_197),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_558),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_408),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_787),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_124),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_189),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_751),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_441),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_677),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_788),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_446),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_769),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_102),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_119),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_80),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_798),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_703),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_791),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_536),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_728),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_664),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_744),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_422),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_332),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_786),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_765),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_764),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_133),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_192),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_60),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_676),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_721),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_715),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_298),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_778),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_279),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_315),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_152),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_430),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_310),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_143),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_733),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_344),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_709),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_539),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_411),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_26),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_283),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_340),
.Y(n_1119)
);

CKINVDCx14_ASAP7_75t_R g1120 ( 
.A(n_670),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_304),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_818),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_270),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_25),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_654),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_736),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_766),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_87),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_371),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_217),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_188),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_151),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_458),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_85),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_683),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_645),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_208),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_530),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_692),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_783),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_749),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_46),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_412),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_7),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_833),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_684),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_521),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_793),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_639),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_518),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_459),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_51),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_789),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_310),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_96),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_440),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_420),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_807),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_601),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_78),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_726),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_101),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_838),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_83),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_472),
.Y(n_1165)
);

BUFx10_ASAP7_75t_L g1166 ( 
.A(n_717),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_232),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_311),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_436),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_415),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_468),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_52),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_702),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_750),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_643),
.Y(n_1175)
);

BUFx10_ASAP7_75t_L g1176 ( 
.A(n_820),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_687),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_101),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_184),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_90),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_206),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_775),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_581),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_135),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_91),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_540),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_365),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_548),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_557),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_815),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_758),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_776),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_319),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_516),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_141),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_382),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_63),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_114),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_209),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_777),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_69),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_704),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_672),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_842),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_792),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_839),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_559),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_351),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_439),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_550),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_471),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_218),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_679),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_187),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_401),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_369),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_110),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_729),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_333),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_570),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_731),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_714),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_661),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_144),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_806),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_142),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_274),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_817),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_646),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_125),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_814),
.Y(n_1231)
);

INVxp33_ASAP7_75t_SL g1232 ( 
.A(n_111),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_830),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_607),
.Y(n_1234)
);

CKINVDCx16_ASAP7_75t_R g1235 ( 
.A(n_542),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_610),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_575),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_173),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_573),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_332),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_774),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_281),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_760),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_166),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_153),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_267),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_553),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_22),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_555),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_825),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_816),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_813),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_55),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_314),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_278),
.Y(n_1255)
);

CKINVDCx14_ASAP7_75t_R g1256 ( 
.A(n_746),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_754),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_140),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_207),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_718),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_363),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_528),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_144),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_290),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_743),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_25),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_96),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_712),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_767),
.Y(n_1269)
);

BUFx10_ASAP7_75t_L g1270 ( 
.A(n_651),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_366),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_829),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_316),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_118),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_723),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_771),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_346),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_587),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_276),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_104),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_223),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_358),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_445),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_647),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_414),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_342),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_629),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_846),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1075),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_860),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1034),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1010),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_880),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1093),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1142),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_900),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1248),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_953),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1006),
.Y(n_1299)
);

INVxp33_ASAP7_75t_SL g1300 ( 
.A(n_847),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_889),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_891),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1014),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_902),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_907),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1069),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_919),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_920),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_939),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1072),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1103),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_963),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_968),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_976),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1127),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1007),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1033),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1037),
.Y(n_1318)
);

INVxp33_ASAP7_75t_L g1319 ( 
.A(n_884),
.Y(n_1319)
);

INVxp33_ASAP7_75t_SL g1320 ( 
.A(n_855),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1038),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_956),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1054),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_999),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_940),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1153),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1061),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1062),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_956),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1063),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1183),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1065),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1024),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_1203),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1071),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1210),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1073),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1228),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1229),
.Y(n_1339)
);

INVxp33_ASAP7_75t_SL g1340 ( 
.A(n_877),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1076),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1233),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1085),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1099),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1241),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1108),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1262),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1111),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1232),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_882),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_883),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1118),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1123),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1128),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1129),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1130),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_888),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_890),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1132),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1322),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1329),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1288),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1333),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1290),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1333),
.B(n_1190),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1303),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1293),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1301),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1302),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1304),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1311),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1306),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1292),
.B(n_1170),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1305),
.B(n_1235),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1307),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1308),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1309),
.Y(n_1377)
);

XOR2xp5_ASAP7_75t_L g1378 ( 
.A(n_1296),
.B(n_861),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1289),
.A2(n_872),
.B1(n_949),
.B2(n_935),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1294),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1312),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1350),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1313),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1325),
.B(n_973),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1314),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1316),
.A2(n_849),
.B(n_848),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1341),
.B(n_1191),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1291),
.B(n_1196),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1317),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1324),
.B(n_896),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1318),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1321),
.B(n_1323),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1327),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1328),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1295),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1300),
.B(n_905),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1330),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1332),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1319),
.B(n_957),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1335),
.B(n_852),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1351),
.B(n_1217),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1337),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1298),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1343),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1344),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1310),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1346),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1348),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1352),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1357),
.B(n_1259),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1315),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1299),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1353),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1354),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1331),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1355),
.B(n_853),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1356),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1359),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1358),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1297),
.B(n_1120),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1385),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1361),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1389),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1393),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1399),
.B(n_1320),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1397),
.Y(n_1426)
);

NAND2xp33_ASAP7_75t_L g1427 ( 
.A(n_1419),
.B(n_1349),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1371),
.B(n_1326),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1398),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1396),
.A2(n_1340),
.B1(n_1144),
.B2(n_1172),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1402),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1404),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1418),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1382),
.B(n_1336),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1370),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1362),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1363),
.Y(n_1437)
);

NAND2xp33_ASAP7_75t_L g1438 ( 
.A(n_1380),
.B(n_956),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1363),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1364),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1367),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1360),
.B(n_1256),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1368),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1395),
.B(n_898),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1370),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1375),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1369),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1381),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1366),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1375),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1394),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1374),
.B(n_1345),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1372),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1376),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1405),
.Y(n_1455)
);

XNOR2xp5_ASAP7_75t_L g1456 ( 
.A(n_1378),
.B(n_1338),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1407),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1376),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1377),
.B(n_863),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1384),
.B(n_1147),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1401),
.A2(n_1193),
.B1(n_961),
.B2(n_1121),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1420),
.B(n_1339),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1373),
.B(n_1342),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1379),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1408),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1387),
.B(n_915),
.C(n_904),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1383),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1383),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1413),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1410),
.B(n_1347),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1406),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_L g1472 ( 
.A(n_1414),
.B(n_1052),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1391),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1391),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1411),
.A2(n_867),
.B1(n_987),
.B2(n_947),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1409),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1388),
.B(n_1134),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1409),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1417),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1417),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1392),
.Y(n_1481)
);

OAI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1390),
.A2(n_1334),
.B1(n_1084),
.B2(n_1187),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_L g1483 ( 
.A(n_1416),
.B(n_1052),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1386),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1400),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1365),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1403),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1412),
.A2(n_1045),
.B1(n_917),
.B2(n_930),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_L g1489 ( 
.A(n_1415),
.B(n_1052),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1385),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1396),
.B(n_926),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1366),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1361),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1361),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1436),
.Y(n_1495)
);

AO22x2_ASAP7_75t_L g1496 ( 
.A1(n_1464),
.A2(n_1487),
.B1(n_1475),
.B2(n_1456),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1440),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1441),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1443),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1492),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_L g1501 ( 
.A(n_1485),
.B(n_936),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1453),
.B(n_927),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1447),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1449),
.B(n_988),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1462),
.B(n_955),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1425),
.B(n_1286),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1486),
.B(n_938),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1471),
.B(n_955),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1448),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1451),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1463),
.B(n_1094),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1422),
.Y(n_1512)
);

AO22x2_ASAP7_75t_L g1513 ( 
.A1(n_1428),
.A2(n_1104),
.B1(n_1164),
.B2(n_1162),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1455),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1457),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1465),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1481),
.B(n_944),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1493),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1469),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1446),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1460),
.B(n_945),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1494),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1480),
.B(n_1281),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1430),
.A2(n_1043),
.B1(n_951),
.B2(n_1177),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1424),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1437),
.B(n_1179),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1446),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1426),
.Y(n_1528)
);

AO22x2_ASAP7_75t_L g1529 ( 
.A1(n_1461),
.A2(n_1184),
.B1(n_1195),
.B2(n_1180),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1429),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1433),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1488),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1421),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1423),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1444),
.B(n_869),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1491),
.A2(n_962),
.B1(n_971),
.B2(n_954),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1452),
.B(n_1434),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1442),
.B(n_975),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1439),
.B(n_1199),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1470),
.B(n_977),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1444),
.B(n_977),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1480),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1431),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1427),
.B(n_1273),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1477),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1454),
.B(n_1201),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1432),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1480),
.B(n_1208),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1435),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1490),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1445),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1473),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1459),
.B(n_1274),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1476),
.B(n_980),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1450),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1458),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1467),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1468),
.B(n_1004),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1474),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1478),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1479),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1484),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1466),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1483),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1489),
.B(n_1224),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1472),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1482),
.A2(n_896),
.B1(n_1166),
.B2(n_1017),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1438),
.B(n_1004),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1446),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1436),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1449),
.B(n_1227),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1449),
.B(n_1230),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1425),
.B(n_997),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1436),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1492),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1425),
.B(n_1005),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1481),
.B(n_1009),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1430),
.B(n_1018),
.C(n_1016),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1436),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1492),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1449),
.B(n_1240),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1436),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1446),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1436),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1481),
.B(n_1027),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1436),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1449),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1422),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1449),
.B(n_1271),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1453),
.B(n_1083),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1481),
.B(n_1036),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1422),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1436),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1453),
.B(n_1083),
.Y(n_1594)
);

BUFx10_ASAP7_75t_L g1595 ( 
.A(n_1492),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1492),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1446),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1425),
.B(n_1280),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1422),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1425),
.B(n_1041),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1422),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1422),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1492),
.B(n_1017),
.Y(n_1603)
);

INVx4_ASAP7_75t_SL g1604 ( 
.A(n_1449),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1446),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1436),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1422),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1422),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1446),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1446),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1449),
.B(n_1244),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1425),
.B(n_1047),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1436),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1436),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1492),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1436),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1425),
.B(n_1060),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1422),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1425),
.B(n_1064),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1449),
.B(n_1258),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1422),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1425),
.B(n_1098),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1436),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1481),
.B(n_1100),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1446),
.Y(n_1625)
);

AO22x2_ASAP7_75t_L g1626 ( 
.A1(n_1464),
.A2(n_1279),
.B1(n_1282),
.B2(n_1277),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1436),
.Y(n_1627)
);

INVx3_ASAP7_75t_R g1628 ( 
.A(n_1453),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1492),
.Y(n_1629)
);

CKINVDCx11_ASAP7_75t_R g1630 ( 
.A(n_1453),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1422),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1436),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1425),
.B(n_1266),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1422),
.Y(n_1634)
);

OA22x2_ASAP7_75t_L g1635 ( 
.A1(n_1461),
.A2(n_1107),
.B1(n_1110),
.B2(n_1106),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1580),
.Y(n_1636)
);

NOR3xp33_ASAP7_75t_SL g1637 ( 
.A(n_1629),
.B(n_1116),
.C(n_1113),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1630),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1496),
.A2(n_1176),
.B1(n_1257),
.B2(n_1166),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1537),
.B(n_1117),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1512),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1587),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1285),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1545),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1517),
.B(n_1119),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1495),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1575),
.Y(n_1647)
);

BUFx10_ASAP7_75t_L g1648 ( 
.A(n_1544),
.Y(n_1648)
);

BUFx4f_ASAP7_75t_L g1649 ( 
.A(n_1589),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1506),
.A2(n_1137),
.B1(n_1143),
.B2(n_1124),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1595),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1497),
.Y(n_1652)
);

NOR2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1596),
.B(n_1152),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1527),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1573),
.B(n_1154),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1498),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1499),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1527),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1615),
.B(n_1155),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1500),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1518),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1576),
.A2(n_1252),
.B(n_859),
.C(n_866),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1558),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1505),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1569),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1628),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1503),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1532),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1577),
.A2(n_854),
.B(n_850),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1520),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1535),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1598),
.B(n_1600),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1509),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1508),
.B(n_892),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1569),
.Y(n_1675)
);

NOR2xp67_ASAP7_75t_L g1676 ( 
.A(n_1542),
.B(n_1272),
.Y(n_1676)
);

INVx6_ASAP7_75t_L g1677 ( 
.A(n_1571),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1626),
.A2(n_1257),
.B1(n_1270),
.B2(n_1176),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1585),
.B(n_1157),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1591),
.B(n_1160),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1529),
.A2(n_1635),
.B1(n_1510),
.B2(n_1515),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1612),
.B(n_1167),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1522),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1588),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1514),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1583),
.B(n_948),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1583),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1624),
.B(n_1168),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1619),
.B(n_1178),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1603),
.B(n_1181),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1597),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1516),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1519),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1597),
.B(n_1021),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1592),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1622),
.B(n_1185),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1599),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1563),
.B(n_1197),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_SL g1699 ( 
.A(n_1617),
.B(n_1212),
.C(n_1198),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1507),
.B(n_1214),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1601),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1570),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1574),
.B(n_1215),
.Y(n_1703)
);

AOI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1534),
.A2(n_870),
.B(n_864),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1579),
.B(n_1582),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1584),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1586),
.B(n_1219),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1602),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1609),
.B(n_1238),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1501),
.A2(n_893),
.B1(n_897),
.B2(n_895),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1593),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1609),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1610),
.B(n_1242),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1606),
.B(n_1245),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1610),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1524),
.A2(n_903),
.B(n_942),
.C(n_906),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1572),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1613),
.B(n_1246),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1578),
.B(n_1253),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1625),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1614),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1616),
.B(n_1254),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1623),
.B(n_1255),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1607),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1627),
.B(n_1261),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1632),
.Y(n_1726)
);

BUFx4f_ASAP7_75t_L g1727 ( 
.A(n_1581),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1608),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1538),
.A2(n_950),
.B(n_943),
.Y(n_1729)
);

INVx5_ASAP7_75t_L g1730 ( 
.A(n_1625),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1543),
.Y(n_1731)
);

NOR2x2_ASAP7_75t_L g1732 ( 
.A(n_1533),
.B(n_1131),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1547),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1540),
.B(n_1263),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1521),
.A2(n_964),
.B(n_974),
.C(n_958),
.Y(n_1735)
);

NOR2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1590),
.B(n_1264),
.Y(n_1736)
);

INVx5_ASAP7_75t_L g1737 ( 
.A(n_1611),
.Y(n_1737)
);

AND2x6_ASAP7_75t_SL g1738 ( 
.A(n_1620),
.B(n_978),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1550),
.B(n_1525),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1594),
.B(n_1267),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1528),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1551),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1504),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1526),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1618),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1530),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1605),
.B(n_1216),
.Y(n_1747)
);

CKINVDCx20_ASAP7_75t_R g1748 ( 
.A(n_1541),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1551),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1559),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1633),
.A2(n_1553),
.B1(n_1568),
.B2(n_1536),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_L g1752 ( 
.A(n_1502),
.B(n_1552),
.C(n_1554),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1621),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1531),
.B(n_1226),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_R g1755 ( 
.A(n_1559),
.B(n_856),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1523),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1631),
.B(n_1634),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1556),
.B(n_979),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1562),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1560),
.B(n_986),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1549),
.B(n_1270),
.Y(n_1761)
);

BUFx12f_ASAP7_75t_L g1762 ( 
.A(n_1511),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1555),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1548),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1557),
.A2(n_996),
.B(n_995),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1539),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1561),
.B(n_1003),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1564),
.B(n_1019),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1566),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1546),
.B(n_857),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1565),
.B(n_875),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1567),
.B(n_862),
.Y(n_1772)
);

OR2x2_ASAP7_75t_SL g1773 ( 
.A(n_1513),
.B(n_1020),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1587),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1587),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1512),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1512),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1545),
.B(n_0),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1495),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1587),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1512),
.Y(n_1781)
);

AND2x4_ASAP7_75t_SL g1782 ( 
.A(n_1595),
.B(n_1022),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1517),
.B(n_1250),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1558),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1537),
.A2(n_1029),
.B1(n_1031),
.B2(n_1025),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1495),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1587),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1517),
.B(n_1265),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1517),
.B(n_1035),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1512),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1517),
.B(n_1039),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1580),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1587),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1558),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1495),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1537),
.A2(n_1057),
.B1(n_1059),
.B2(n_1049),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1512),
.Y(n_1797)
);

INVx5_ASAP7_75t_L g1798 ( 
.A(n_1595),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1495),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1587),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1512),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1587),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1517),
.B(n_1067),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1537),
.B(n_1068),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1495),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1587),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1495),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1512),
.Y(n_1808)
);

INVx4_ASAP7_75t_L g1809 ( 
.A(n_1629),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1496),
.A2(n_910),
.B1(n_1095),
.B2(n_1032),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1517),
.A2(n_1077),
.B1(n_1082),
.B2(n_1070),
.Y(n_1811)
);

NOR3xp33_ASAP7_75t_SL g1812 ( 
.A(n_1629),
.B(n_868),
.C(n_865),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1495),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1587),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1512),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1517),
.B(n_1126),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1587),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1587),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1587),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1495),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1512),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1629),
.Y(n_1822)
);

AND2x2_ASAP7_75t_SL g1823 ( 
.A(n_1603),
.B(n_1044),
.Y(n_1823)
);

INVx5_ASAP7_75t_L g1824 ( 
.A(n_1595),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1537),
.B(n_871),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1537),
.A2(n_1139),
.B1(n_1141),
.B2(n_1136),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1495),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1580),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1587),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1495),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1517),
.B(n_1161),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1672),
.B(n_1284),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1646),
.Y(n_1833)
);

AND2x6_ASAP7_75t_L g1834 ( 
.A(n_1652),
.B(n_1163),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1741),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1746),
.Y(n_1836)
);

O2A1O1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1640),
.A2(n_1204),
.B(n_1211),
.C(n_1200),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1656),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1657),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1667),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1775),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1644),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1682),
.B(n_873),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1673),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1696),
.B(n_874),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1647),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1804),
.B(n_876),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1677),
.B(n_845),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1664),
.A2(n_1251),
.B1(n_1221),
.B2(n_993),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1775),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1641),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1715),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1661),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1823),
.B(n_1269),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1648),
.B(n_1275),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1683),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1645),
.B(n_0),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1715),
.Y(n_1858)
);

INVx5_ASAP7_75t_L g1859 ( 
.A(n_1806),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1783),
.A2(n_1058),
.B(n_1148),
.C(n_922),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1685),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1734),
.B(n_1655),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1692),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1689),
.B(n_1),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1660),
.B(n_878),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1693),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1668),
.B(n_1236),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1717),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1787),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1702),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1706),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1727),
.B(n_1225),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1730),
.B(n_1670),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1711),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1788),
.B(n_1789),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1721),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1791),
.B(n_1),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1726),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1792),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1806),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1740),
.B(n_1674),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1803),
.B(n_2),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1663),
.B(n_2),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1816),
.B(n_3),
.Y(n_1884)
);

CKINVDCx8_ASAP7_75t_R g1885 ( 
.A(n_1638),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1779),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1684),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1695),
.Y(n_1888)
);

BUFx8_ASAP7_75t_L g1889 ( 
.A(n_1814),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1831),
.B(n_3),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1730),
.B(n_886),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1830),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1737),
.B(n_1243),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1786),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1795),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1636),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1697),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1799),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1705),
.B(n_4),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1744),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1700),
.B(n_4),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1805),
.Y(n_1902)
);

NAND2xp33_ASAP7_75t_L g1903 ( 
.A(n_1798),
.B(n_1001),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1807),
.B(n_5),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1813),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1814),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1701),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1762),
.B(n_887),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1819),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1820),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1819),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1827),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1784),
.B(n_879),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1829),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1731),
.B(n_5),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1828),
.Y(n_1916)
);

INVx4_ASAP7_75t_L g1917 ( 
.A(n_1829),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1794),
.B(n_6),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1774),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1733),
.B(n_6),
.Y(n_1920)
);

INVx5_ASAP7_75t_L g1921 ( 
.A(n_1798),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1708),
.Y(n_1922)
);

BUFx3_ASAP7_75t_L g1923 ( 
.A(n_1793),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1724),
.Y(n_1924)
);

AND3x1_ASAP7_75t_L g1925 ( 
.A(n_1637),
.B(n_1699),
.C(n_1812),
.Y(n_1925)
);

INVx5_ASAP7_75t_L g1926 ( 
.A(n_1824),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1759),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1809),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1675),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1802),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1675),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1681),
.B(n_7),
.Y(n_1932)
);

O2A1O1Ixp5_ASAP7_75t_L g1933 ( 
.A1(n_1729),
.A2(n_1825),
.B(n_1811),
.C(n_1662),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1737),
.B(n_1283),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1649),
.B(n_8),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1739),
.Y(n_1936)
);

NOR2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1822),
.B(n_881),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1728),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1761),
.B(n_8),
.Y(n_1939)
);

INVx4_ASAP7_75t_L g1940 ( 
.A(n_1824),
.Y(n_1940)
);

INVxp67_ASAP7_75t_L g1941 ( 
.A(n_1778),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1751),
.B(n_1826),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1748),
.A2(n_899),
.B1(n_901),
.B2(n_885),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1742),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1757),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1686),
.B(n_894),
.Y(n_1946)
);

BUFx8_ASAP7_75t_SL g1947 ( 
.A(n_1800),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1745),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1763),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1750),
.Y(n_1950)
);

BUFx12f_ASAP7_75t_L g1951 ( 
.A(n_1671),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1769),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1752),
.B(n_908),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1753),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1712),
.Y(n_1955)
);

AND2x4_ASAP7_75t_SL g1956 ( 
.A(n_1818),
.B(n_851),
.Y(n_1956)
);

NOR2xp67_ASAP7_75t_L g1957 ( 
.A(n_1642),
.B(n_909),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1776),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1780),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1817),
.B(n_1237),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1749),
.Y(n_1961)
);

AND2x6_ASAP7_75t_L g1962 ( 
.A(n_1651),
.B(n_984),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1777),
.Y(n_1963)
);

A2O1A1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1785),
.A2(n_1151),
.B(n_1234),
.C(n_1149),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1796),
.B(n_9),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1781),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1790),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1743),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1686),
.B(n_9),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1716),
.B(n_10),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1797),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1801),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1808),
.Y(n_1973)
);

INVx4_ASAP7_75t_L g1974 ( 
.A(n_1694),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1719),
.B(n_1703),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1815),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1873),
.B(n_1766),
.Y(n_1977)
);

INVx1_ASAP7_75t_SL g1978 ( 
.A(n_1879),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1846),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1858),
.Y(n_1980)
);

AND2x6_ASAP7_75t_L g1981 ( 
.A(n_1936),
.B(n_1821),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1835),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1885),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1944),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1842),
.B(n_1694),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1847),
.A2(n_1810),
.B1(n_1639),
.B2(n_1678),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1836),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1881),
.B(n_1935),
.Y(n_1988)
);

NAND2x1p5_ASAP7_75t_L g1989 ( 
.A(n_1859),
.B(n_1654),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1868),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1969),
.B(n_1736),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1833),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1942),
.A2(n_1650),
.B1(n_1772),
.B2(n_1747),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1851),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1843),
.A2(n_1710),
.B1(n_1764),
.B2(n_1690),
.Y(n_1995)
);

INVx4_ASAP7_75t_L g1996 ( 
.A(n_1950),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1834),
.A2(n_1770),
.B1(n_1755),
.B2(n_1765),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1875),
.B(n_1658),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1889),
.Y(n_1999)
);

AOI21xp33_ASAP7_75t_L g2000 ( 
.A1(n_1845),
.A2(n_1698),
.B(n_1735),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1838),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1968),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1862),
.B(n_1687),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1859),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1839),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1840),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1947),
.Y(n_2007)
);

OR2x6_ASAP7_75t_L g2008 ( 
.A(n_1946),
.B(n_1666),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1941),
.B(n_1782),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1853),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1844),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1856),
.Y(n_2012)
);

A2O1A1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_1837),
.A2(n_1679),
.B(n_1688),
.C(n_1680),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1921),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1861),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1887),
.Y(n_2016)
);

A2O1A1Ixp33_ASAP7_75t_SL g2017 ( 
.A1(n_1864),
.A2(n_1669),
.B(n_1714),
.C(n_1707),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1900),
.B(n_1773),
.Y(n_2018)
);

BUFx4f_ASAP7_75t_L g2019 ( 
.A(n_1951),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1975),
.B(n_1738),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1921),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1863),
.Y(n_2022)
);

BUFx8_ASAP7_75t_L g2023 ( 
.A(n_1896),
.Y(n_2023)
);

BUFx8_ASAP7_75t_SL g2024 ( 
.A(n_1916),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1866),
.Y(n_2025)
);

AOI222xp33_ASAP7_75t_L g2026 ( 
.A1(n_1932),
.A2(n_1834),
.B1(n_1965),
.B2(n_1854),
.C1(n_1865),
.C2(n_1871),
.Y(n_2026)
);

O2A1O1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1939),
.A2(n_1659),
.B(n_1722),
.C(n_1718),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1869),
.B(n_1691),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1877),
.A2(n_1725),
.B1(n_1723),
.B2(n_1676),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_1841),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1888),
.Y(n_2031)
);

INVx5_ASAP7_75t_L g2032 ( 
.A(n_1926),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1897),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1926),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1870),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1930),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1907),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1945),
.B(n_1834),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_1906),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_1953),
.A2(n_1643),
.B1(n_1653),
.B2(n_1709),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_1929),
.Y(n_2041)
);

OR2x6_ASAP7_75t_L g2042 ( 
.A(n_1946),
.B(n_1974),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1882),
.A2(n_1713),
.B1(n_1768),
.B2(n_1720),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1874),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1876),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1878),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_1906),
.Y(n_2047)
);

A2O1A1Ixp33_ASAP7_75t_L g2048 ( 
.A1(n_1933),
.A2(n_1767),
.B(n_1758),
.C(n_1760),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1955),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1955),
.B(n_1665),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1867),
.B(n_1756),
.Y(n_2051)
);

INVx4_ASAP7_75t_L g2052 ( 
.A(n_1909),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1886),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1909),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1892),
.B(n_1754),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1922),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1894),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1883),
.B(n_1771),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1924),
.Y(n_2059)
);

OR2x6_ASAP7_75t_L g2060 ( 
.A(n_1908),
.B(n_1732),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1895),
.B(n_1704),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1976),
.A2(n_1268),
.B1(n_858),
.B2(n_921),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1898),
.B(n_10),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1884),
.A2(n_1890),
.B(n_1901),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1938),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1918),
.B(n_11),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1902),
.Y(n_2067)
);

A2O1A1Ixp33_ASAP7_75t_L g2068 ( 
.A1(n_1857),
.A2(n_912),
.B(n_913),
.C(n_911),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1919),
.B(n_423),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1905),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1832),
.A2(n_858),
.B(n_851),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1948),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1954),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1899),
.A2(n_1860),
.B(n_1903),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1910),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1943),
.B(n_1913),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1904),
.A2(n_916),
.B1(n_918),
.B2(n_914),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1961),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1958),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1911),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1912),
.B(n_11),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1927),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1949),
.Y(n_2083)
);

INVxp67_ASAP7_75t_SL g2084 ( 
.A(n_1952),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_1961),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1850),
.B(n_12),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1915),
.A2(n_1249),
.B(n_858),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1923),
.B(n_424),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1967),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1880),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1929),
.B(n_12),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1963),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1931),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1972),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1931),
.B(n_1962),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1917),
.B(n_923),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1920),
.A2(n_925),
.B1(n_928),
.B2(n_924),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1973),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1914),
.B(n_13),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1970),
.A2(n_921),
.B(n_851),
.Y(n_2100)
);

NAND2x1p5_ASAP7_75t_L g2101 ( 
.A(n_1852),
.B(n_921),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_1928),
.B(n_425),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1971),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1966),
.Y(n_2104)
);

A2O1A1Ixp33_ASAP7_75t_L g2105 ( 
.A1(n_1964),
.A2(n_931),
.B(n_933),
.C(n_929),
.Y(n_2105)
);

OAI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_1849),
.A2(n_941),
.B1(n_946),
.B2(n_937),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1940),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1959),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1956),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1957),
.B(n_1231),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1891),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1962),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1962),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1848),
.B(n_13),
.Y(n_2114)
);

BUFx8_ASAP7_75t_L g2115 ( 
.A(n_1908),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1848),
.B(n_1925),
.Y(n_2116)
);

OAI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1855),
.A2(n_934),
.B1(n_959),
.B2(n_952),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_1937),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1893),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_1872),
.A2(n_966),
.B1(n_1133),
.B2(n_932),
.Y(n_2120)
);

INVxp67_ASAP7_75t_SL g2121 ( 
.A(n_1934),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1960),
.A2(n_960),
.B1(n_967),
.B2(n_965),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1835),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_2002),
.Y(n_2124)
);

OAI21x1_ASAP7_75t_L g2125 ( 
.A1(n_2100),
.A2(n_1001),
.B(n_429),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1988),
.B(n_14),
.Y(n_2126)
);

CKINVDCx20_ASAP7_75t_R g2127 ( 
.A(n_1983),
.Y(n_2127)
);

OAI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2076),
.A2(n_966),
.B1(n_1133),
.B2(n_932),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2085),
.Y(n_2129)
);

AO21x1_ASAP7_75t_L g2130 ( 
.A1(n_2064),
.A2(n_1001),
.B(n_15),
.Y(n_2130)
);

OAI21x1_ASAP7_75t_L g2131 ( 
.A1(n_2087),
.A2(n_1001),
.B(n_432),
.Y(n_2131)
);

OAI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_1995),
.A2(n_966),
.B1(n_1133),
.B2(n_932),
.Y(n_2132)
);

INVx6_ASAP7_75t_L g2133 ( 
.A(n_2032),
.Y(n_2133)
);

INVxp33_ASAP7_75t_L g2134 ( 
.A(n_2051),
.Y(n_2134)
);

INVx1_ASAP7_75t_SL g2135 ( 
.A(n_2030),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_2061),
.A2(n_1001),
.B(n_433),
.Y(n_2136)
);

AOI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_2048),
.A2(n_1189),
.B(n_1135),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_2074),
.A2(n_434),
.B(n_427),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1982),
.Y(n_2139)
);

OAI21x1_ASAP7_75t_L g2140 ( 
.A1(n_2071),
.A2(n_437),
.B(n_435),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2066),
.B(n_15),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2123),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2103),
.Y(n_2143)
);

OA21x2_ASAP7_75t_L g2144 ( 
.A1(n_2038),
.A2(n_970),
.B(n_969),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_L g2145 ( 
.A1(n_1992),
.A2(n_443),
.B(n_438),
.Y(n_2145)
);

NOR2x1_ASAP7_75t_SL g2146 ( 
.A(n_2032),
.B(n_1135),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1987),
.Y(n_2147)
);

OAI21x1_ASAP7_75t_L g2148 ( 
.A1(n_2001),
.A2(n_447),
.B(n_444),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1977),
.B(n_16),
.Y(n_2149)
);

CKINVDCx14_ASAP7_75t_R g2150 ( 
.A(n_1999),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2104),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1994),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2005),
.Y(n_2153)
);

OAI21x1_ASAP7_75t_L g2154 ( 
.A1(n_2006),
.A2(n_451),
.B(n_449),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2011),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2015),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2020),
.A2(n_1249),
.B1(n_1189),
.B2(n_1135),
.Y(n_2157)
);

OA21x2_ASAP7_75t_L g2158 ( 
.A1(n_2000),
.A2(n_2084),
.B(n_2025),
.Y(n_2158)
);

A2O1A1Ixp33_ASAP7_75t_L g2159 ( 
.A1(n_2027),
.A2(n_981),
.B(n_982),
.C(n_972),
.Y(n_2159)
);

OAI21x1_ASAP7_75t_L g2160 ( 
.A1(n_2022),
.A2(n_455),
.B(n_452),
.Y(n_2160)
);

OAI21x1_ASAP7_75t_L g2161 ( 
.A1(n_2035),
.A2(n_457),
.B(n_456),
.Y(n_2161)
);

OAI21x1_ASAP7_75t_L g2162 ( 
.A1(n_2044),
.A2(n_461),
.B(n_460),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1984),
.B(n_16),
.Y(n_2163)
);

INVx2_ASAP7_75t_SL g2164 ( 
.A(n_2004),
.Y(n_2164)
);

OAI21x1_ASAP7_75t_SL g2165 ( 
.A1(n_2029),
.A2(n_17),
.B(n_18),
.Y(n_2165)
);

OAI21x1_ASAP7_75t_L g2166 ( 
.A1(n_2045),
.A2(n_464),
.B(n_463),
.Y(n_2166)
);

OR2x6_ASAP7_75t_L g2167 ( 
.A(n_2060),
.B(n_1189),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2026),
.A2(n_985),
.B1(n_989),
.B2(n_983),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2046),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2081),
.B(n_17),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2047),
.B(n_2004),
.Y(n_2171)
);

OAI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2060),
.A2(n_1249),
.B1(n_991),
.B2(n_992),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1991),
.B(n_18),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2053),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2010),
.Y(n_2175)
);

OR2x6_ASAP7_75t_L g2176 ( 
.A(n_2042),
.B(n_465),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2057),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_2049),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2067),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_1990),
.B(n_19),
.Y(n_2180)
);

O2A1O1Ixp33_ASAP7_75t_SL g2181 ( 
.A1(n_2013),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_2181)
);

OAI21x1_ASAP7_75t_L g2182 ( 
.A1(n_2070),
.A2(n_467),
.B(n_466),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2114),
.B(n_20),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_2024),
.Y(n_2184)
);

OA21x2_ASAP7_75t_L g2185 ( 
.A1(n_2075),
.A2(n_2083),
.B(n_2082),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_1986),
.A2(n_994),
.B1(n_998),
.B2(n_990),
.Y(n_2186)
);

AO21x2_ASAP7_75t_L g2187 ( 
.A1(n_2017),
.A2(n_1002),
.B(n_1000),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2050),
.B(n_21),
.Y(n_2188)
);

OAI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_1997),
.A2(n_1011),
.B1(n_1013),
.B2(n_1008),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_2112),
.A2(n_2113),
.B(n_2092),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_SL g2191 ( 
.A1(n_2063),
.A2(n_22),
.B(n_23),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_2042),
.B(n_23),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1996),
.B(n_24),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_L g2194 ( 
.A1(n_2043),
.A2(n_470),
.B(n_469),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2012),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1998),
.B(n_24),
.Y(n_2196)
);

AOI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_1981),
.A2(n_1015),
.B1(n_1023),
.B2(n_1012),
.Y(n_2197)
);

BUFx12f_ASAP7_75t_L g2198 ( 
.A(n_2007),
.Y(n_2198)
);

OAI21x1_ASAP7_75t_L g2199 ( 
.A1(n_2055),
.A2(n_476),
.B(n_474),
.Y(n_2199)
);

NAND2x1p5_ASAP7_75t_L g2200 ( 
.A(n_2049),
.B(n_477),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2016),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_2101),
.A2(n_480),
.B(n_479),
.Y(n_2202)
);

INVxp67_ASAP7_75t_SL g2203 ( 
.A(n_2036),
.Y(n_2203)
);

OAI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_2003),
.A2(n_1028),
.B(n_1026),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_SL g2205 ( 
.A1(n_2091),
.A2(n_26),
.B(n_27),
.Y(n_2205)
);

NOR2x1_ASAP7_75t_L g2206 ( 
.A(n_2021),
.B(n_1030),
.Y(n_2206)
);

NOR2xp67_ASAP7_75t_SL g2207 ( 
.A(n_2116),
.B(n_1223),
.Y(n_2207)
);

O2A1O1Ixp5_ASAP7_75t_L g2208 ( 
.A1(n_2121),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_SL g2209 ( 
.A1(n_2118),
.A2(n_28),
.B(n_29),
.Y(n_2209)
);

OAI22xp33_ASAP7_75t_L g2210 ( 
.A1(n_2018),
.A2(n_1042),
.B1(n_1046),
.B2(n_1040),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2031),
.Y(n_2211)
);

OAI21x1_ASAP7_75t_L g2212 ( 
.A1(n_2095),
.A2(n_483),
.B(n_481),
.Y(n_2212)
);

BUFx8_ASAP7_75t_L g2213 ( 
.A(n_2078),
.Y(n_2213)
);

OAI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2068),
.A2(n_1050),
.B(n_1048),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2033),
.Y(n_2215)
);

OA21x2_ASAP7_75t_L g2216 ( 
.A1(n_2105),
.A2(n_1053),
.B(n_1051),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2037),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_2056),
.A2(n_485),
.B(n_484),
.Y(n_2218)
);

OA21x2_ASAP7_75t_L g2219 ( 
.A1(n_2062),
.A2(n_1056),
.B(n_1055),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2090),
.B(n_30),
.Y(n_2220)
);

AO21x1_ASAP7_75t_L g2221 ( 
.A1(n_2077),
.A2(n_30),
.B(n_31),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_SL g2222 ( 
.A1(n_2119),
.A2(n_1985),
.B1(n_1978),
.B2(n_1979),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_2028),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2126),
.B(n_2086),
.Y(n_2224)
);

CKINVDCx11_ASAP7_75t_R g2225 ( 
.A(n_2127),
.Y(n_2225)
);

OAI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_2186),
.A2(n_1993),
.B1(n_2040),
.B2(n_2097),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2143),
.Y(n_2227)
);

O2A1O1Ixp33_ASAP7_75t_SL g2228 ( 
.A1(n_2159),
.A2(n_2014),
.B(n_2110),
.C(n_2034),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2151),
.Y(n_2229)
);

AOI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2181),
.A2(n_2106),
.B1(n_2117),
.B2(n_2009),
.C(n_2099),
.Y(n_2230)
);

AO31x2_ASAP7_75t_L g2231 ( 
.A1(n_2130),
.A2(n_2059),
.A3(n_2072),
.B(n_2065),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2185),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_2203),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2153),
.Y(n_2234)
);

AOI22xp33_ASAP7_75t_L g2235 ( 
.A1(n_2221),
.A2(n_1981),
.B1(n_2115),
.B2(n_2079),
.Y(n_2235)
);

NAND2xp33_ASAP7_75t_R g2236 ( 
.A(n_2167),
.B(n_2008),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2155),
.Y(n_2237)
);

AOI22xp33_ASAP7_75t_SL g2238 ( 
.A1(n_2222),
.A2(n_1981),
.B1(n_2058),
.B2(n_2111),
.Y(n_2238)
);

AOI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2137),
.A2(n_2102),
.B(n_2088),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2156),
.Y(n_2240)
);

AOI21x1_ASAP7_75t_L g2241 ( 
.A1(n_2158),
.A2(n_2008),
.B(n_2109),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2128),
.A2(n_2069),
.B(n_2120),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2169),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2142),
.Y(n_2244)
);

INVx4_ASAP7_75t_L g2245 ( 
.A(n_2184),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_2178),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2124),
.B(n_2108),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_2133),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2152),
.Y(n_2249)
);

BUFx2_ASAP7_75t_L g2250 ( 
.A(n_2223),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2174),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2175),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2177),
.Y(n_2253)
);

OAI22xp5_ASAP7_75t_SL g2254 ( 
.A1(n_2150),
.A2(n_2052),
.B1(n_2054),
.B2(n_2039),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2168),
.A2(n_2019),
.B1(n_2122),
.B2(n_1980),
.Y(n_2255)
);

A2O1A1Ixp33_ASAP7_75t_L g2256 ( 
.A1(n_2204),
.A2(n_2096),
.B(n_2041),
.C(n_2093),
.Y(n_2256)
);

AOI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_2157),
.A2(n_2089),
.B1(n_2094),
.B2(n_2073),
.Y(n_2257)
);

NAND2x1p5_ASAP7_75t_L g2258 ( 
.A(n_2135),
.B(n_2078),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2179),
.B(n_2023),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2180),
.B(n_2098),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2132),
.A2(n_1989),
.B(n_2080),
.Y(n_2261)
);

CKINVDCx11_ASAP7_75t_R g2262 ( 
.A(n_2198),
.Y(n_2262)
);

INVx4_ASAP7_75t_L g2263 ( 
.A(n_2133),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2208),
.B(n_2107),
.C(n_1074),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_SL g2265 ( 
.A1(n_2165),
.A2(n_2107),
.B1(n_1078),
.B2(n_1079),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2139),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2147),
.B(n_2134),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2195),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2201),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2211),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2213),
.Y(n_2271)
);

OAI221xp5_ASAP7_75t_L g2272 ( 
.A1(n_2193),
.A2(n_1081),
.B1(n_1086),
.B2(n_1080),
.C(n_1066),
.Y(n_2272)
);

OAI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2194),
.A2(n_1088),
.B(n_1087),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2176),
.A2(n_2167),
.B1(n_2192),
.B2(n_2149),
.Y(n_2274)
);

NAND2xp33_ASAP7_75t_R g2275 ( 
.A(n_2176),
.B(n_32),
.Y(n_2275)
);

AO21x2_ASAP7_75t_L g2276 ( 
.A1(n_2136),
.A2(n_1213),
.B(n_1209),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2197),
.A2(n_1125),
.B1(n_1159),
.B2(n_1101),
.Y(n_2277)
);

NAND2x1p5_ASAP7_75t_L g2278 ( 
.A(n_2171),
.B(n_487),
.Y(n_2278)
);

BUFx2_ASAP7_75t_L g2279 ( 
.A(n_2233),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2251),
.Y(n_2280)
);

NOR3xp33_ASAP7_75t_SL g2281 ( 
.A(n_2275),
.B(n_2163),
.C(n_2210),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_SL g2282 ( 
.A1(n_2226),
.A2(n_2170),
.B1(n_2191),
.B2(n_2205),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2234),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2237),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_2225),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_2250),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_2238),
.A2(n_2144),
.B1(n_2216),
.B2(n_2215),
.Y(n_2287)
);

CKINVDCx16_ASAP7_75t_R g2288 ( 
.A(n_2271),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2240),
.B(n_2196),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2268),
.Y(n_2290)
);

BUFx2_ASAP7_75t_L g2291 ( 
.A(n_2247),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2243),
.B(n_2141),
.Y(n_2292)
);

AND4x1_ASAP7_75t_L g2293 ( 
.A(n_2274),
.B(n_2207),
.C(n_2206),
.D(n_2173),
.Y(n_2293)
);

AOI211xp5_ASAP7_75t_L g2294 ( 
.A1(n_2272),
.A2(n_2172),
.B(n_2255),
.C(n_2239),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2253),
.Y(n_2295)
);

AO21x1_ASAP7_75t_L g2296 ( 
.A1(n_2259),
.A2(n_2220),
.B(n_2189),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2235),
.A2(n_2217),
.B1(n_2219),
.B2(n_2183),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_2262),
.Y(n_2298)
);

CKINVDCx16_ASAP7_75t_R g2299 ( 
.A(n_2254),
.Y(n_2299)
);

HB1xp67_ASAP7_75t_L g2300 ( 
.A(n_2267),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2266),
.B(n_2129),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2265),
.A2(n_2200),
.B1(n_2188),
.B2(n_2214),
.Y(n_2302)
);

AO32x2_ASAP7_75t_L g2303 ( 
.A1(n_2248),
.A2(n_2164),
.A3(n_2190),
.B1(n_2209),
.B2(n_2187),
.Y(n_2303)
);

OR2x6_ASAP7_75t_L g2304 ( 
.A(n_2263),
.B(n_2199),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_2246),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2260),
.B(n_31),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2269),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2270),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_SL g2309 ( 
.A(n_2264),
.B(n_1090),
.C(n_1089),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_2245),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2224),
.B(n_2145),
.Y(n_2311)
);

CKINVDCx16_ASAP7_75t_R g2312 ( 
.A(n_2236),
.Y(n_2312)
);

HB1xp67_ASAP7_75t_L g2313 ( 
.A(n_2231),
.Y(n_2313)
);

OR2x6_ASAP7_75t_L g2314 ( 
.A(n_2261),
.B(n_2212),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2258),
.B(n_2229),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_2256),
.B(n_33),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2227),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_2241),
.A2(n_2138),
.B(n_2125),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2232),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2244),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2228),
.B(n_33),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2249),
.B(n_34),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2252),
.B(n_2148),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2231),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2230),
.A2(n_1092),
.B1(n_1096),
.B2(n_1091),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2278),
.B(n_2154),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2276),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_2257),
.Y(n_2328)
);

AOI21x1_ASAP7_75t_L g2329 ( 
.A1(n_2273),
.A2(n_2131),
.B(n_2160),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_2242),
.Y(n_2330)
);

A2O1A1Ixp33_ASAP7_75t_L g2331 ( 
.A1(n_2277),
.A2(n_2166),
.B(n_2182),
.C(n_2162),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_2225),
.Y(n_2332)
);

CKINVDCx12_ASAP7_75t_R g2333 ( 
.A(n_2254),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_2225),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2268),
.Y(n_2335)
);

O2A1O1Ixp33_ASAP7_75t_L g2336 ( 
.A1(n_2226),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2280),
.Y(n_2337)
);

AO31x2_ASAP7_75t_L g2338 ( 
.A1(n_2324),
.A2(n_2146),
.A3(n_2161),
.B(n_2218),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2290),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2283),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2286),
.B(n_2202),
.Y(n_2341)
);

OR2x2_ASAP7_75t_L g2342 ( 
.A(n_2300),
.B(n_35),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2284),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2279),
.B(n_2140),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2295),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2307),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2308),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2291),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2319),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2288),
.B(n_36),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2305),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2311),
.B(n_37),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2335),
.Y(n_2353)
);

INVxp67_ASAP7_75t_SL g2354 ( 
.A(n_2313),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2317),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2289),
.B(n_2301),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2315),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2320),
.Y(n_2358)
);

INVx5_ASAP7_75t_L g2359 ( 
.A(n_2314),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2292),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2323),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2322),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2330),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2299),
.B(n_37),
.Y(n_2364)
);

CKINVDCx6p67_ASAP7_75t_R g2365 ( 
.A(n_2333),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2306),
.B(n_38),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2312),
.B(n_38),
.Y(n_2367)
);

BUFx3_ASAP7_75t_L g2368 ( 
.A(n_2285),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2298),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2327),
.B(n_39),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2330),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2303),
.Y(n_2372)
);

OR2x2_ASAP7_75t_L g2373 ( 
.A(n_2296),
.B(n_39),
.Y(n_2373)
);

INVx5_ASAP7_75t_L g2374 ( 
.A(n_2314),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2332),
.B(n_40),
.Y(n_2375)
);

BUFx3_ASAP7_75t_L g2376 ( 
.A(n_2334),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2304),
.B(n_40),
.Y(n_2377)
);

HB1xp67_ASAP7_75t_L g2378 ( 
.A(n_2304),
.Y(n_2378)
);

BUFx3_ASAP7_75t_L g2379 ( 
.A(n_2310),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2326),
.B(n_41),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2281),
.B(n_41),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2303),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2316),
.B(n_42),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_2309),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2321),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2282),
.B(n_42),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2318),
.Y(n_2387)
);

INVx2_ASAP7_75t_SL g2388 ( 
.A(n_2293),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2294),
.B(n_43),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2328),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2331),
.A2(n_1102),
.B(n_1097),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2329),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2302),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2325),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2336),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2297),
.Y(n_2396)
);

INVx1_ASAP7_75t_SL g2397 ( 
.A(n_2287),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2286),
.B(n_43),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2280),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2290),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2286),
.B(n_44),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2280),
.Y(n_2402)
);

BUFx4f_ASAP7_75t_L g2403 ( 
.A(n_2330),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2279),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_2279),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2286),
.B(n_44),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2299),
.B(n_45),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2279),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2286),
.B(n_45),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2299),
.B(n_47),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2286),
.B(n_47),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2280),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2280),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2279),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2279),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2290),
.Y(n_2416)
);

BUFx2_ASAP7_75t_L g2417 ( 
.A(n_2279),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_SL g2418 ( 
.A(n_2385),
.B(n_2403),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2348),
.B(n_48),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2356),
.B(n_2362),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2349),
.Y(n_2421)
);

AOI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2391),
.A2(n_2395),
.B(n_2383),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2404),
.B(n_48),
.Y(n_2423)
);

OAI221xp5_ASAP7_75t_SL g2424 ( 
.A1(n_2373),
.A2(n_2386),
.B1(n_2389),
.B2(n_2381),
.C(n_2407),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_2365),
.B(n_49),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_2351),
.Y(n_2426)
);

NAND4xp25_ASAP7_75t_L g2427 ( 
.A(n_2398),
.B(n_2409),
.C(n_2411),
.D(n_2401),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2405),
.B(n_49),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2408),
.B(n_51),
.Y(n_2429)
);

OAI21xp5_ASAP7_75t_L g2430 ( 
.A1(n_2410),
.A2(n_2364),
.B(n_2393),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2417),
.B(n_52),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2414),
.B(n_53),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2415),
.B(n_53),
.Y(n_2433)
);

OAI221xp5_ASAP7_75t_SL g2434 ( 
.A1(n_2377),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.C(n_57),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2360),
.B(n_54),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2337),
.B(n_56),
.Y(n_2436)
);

NAND3xp33_ASAP7_75t_L g2437 ( 
.A(n_2382),
.B(n_1109),
.C(n_1105),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2357),
.B(n_57),
.Y(n_2438)
);

OA21x2_ASAP7_75t_L g2439 ( 
.A1(n_2372),
.A2(n_1114),
.B(n_1112),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2399),
.B(n_58),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2378),
.B(n_58),
.Y(n_2441)
);

OAI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2394),
.A2(n_1122),
.B1(n_1138),
.B2(n_1115),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2368),
.B(n_59),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2402),
.B(n_2412),
.Y(n_2444)
);

OAI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_2388),
.A2(n_2380),
.B1(n_2342),
.B2(n_2397),
.Y(n_2445)
);

OAI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2359),
.A2(n_1171),
.B1(n_1140),
.B2(n_1146),
.Y(n_2446)
);

AOI211xp5_ASAP7_75t_L g2447 ( 
.A1(n_2350),
.A2(n_69),
.B(n_77),
.C(n_59),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2413),
.B(n_60),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_SL g2449 ( 
.A1(n_2341),
.A2(n_1150),
.B(n_1145),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2352),
.B(n_61),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2359),
.B(n_1156),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2340),
.B(n_61),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_L g2453 ( 
.A1(n_2396),
.A2(n_1165),
.B1(n_1169),
.B2(n_1158),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2343),
.B(n_64),
.Y(n_2454)
);

OAI21xp33_ASAP7_75t_L g2455 ( 
.A1(n_2352),
.A2(n_64),
.B(n_65),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2345),
.B(n_66),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2376),
.B(n_66),
.Y(n_2457)
);

NAND3xp33_ASAP7_75t_L g2458 ( 
.A(n_2392),
.B(n_1174),
.C(n_1173),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2361),
.B(n_67),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2354),
.B(n_67),
.Y(n_2460)
);

OAI22xp5_ASAP7_75t_L g2461 ( 
.A1(n_2406),
.A2(n_1182),
.B1(n_1186),
.B2(n_1175),
.Y(n_2461)
);

OAI21xp5_ASAP7_75t_SL g2462 ( 
.A1(n_2375),
.A2(n_68),
.B(n_70),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2374),
.B(n_1188),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2370),
.B(n_68),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2358),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2363),
.B(n_2371),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2379),
.B(n_71),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2374),
.B(n_2369),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2344),
.B(n_2366),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2387),
.B(n_72),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2339),
.B(n_72),
.Y(n_2471)
);

OAI221xp5_ASAP7_75t_L g2472 ( 
.A1(n_2367),
.A2(n_1202),
.B1(n_1205),
.B2(n_1194),
.C(n_1192),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2346),
.B(n_73),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2347),
.B(n_73),
.Y(n_2474)
);

OAI21xp5_ASAP7_75t_SL g2475 ( 
.A1(n_2390),
.A2(n_74),
.B(n_75),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2353),
.B(n_74),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2400),
.B(n_75),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2416),
.B(n_76),
.Y(n_2478)
);

AOI221xp5_ASAP7_75t_L g2479 ( 
.A1(n_2384),
.A2(n_1218),
.B1(n_1220),
.B2(n_1207),
.C(n_1206),
.Y(n_2479)
);

OAI221xp5_ASAP7_75t_SL g2480 ( 
.A1(n_2355),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2338),
.B(n_79),
.Y(n_2481)
);

OAI221xp5_ASAP7_75t_L g2482 ( 
.A1(n_2338),
.A2(n_1247),
.B1(n_1260),
.B2(n_1239),
.C(n_1222),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2348),
.B(n_80),
.Y(n_2483)
);

OAI21xp5_ASAP7_75t_SL g2484 ( 
.A1(n_2389),
.A2(n_81),
.B(n_82),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2348),
.B(n_81),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2348),
.B(n_82),
.Y(n_2486)
);

NAND3xp33_ASAP7_75t_L g2487 ( 
.A(n_2385),
.B(n_1278),
.C(n_1276),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2385),
.B(n_1287),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2361),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2348),
.B(n_83),
.Y(n_2490)
);

AOI221xp5_ASAP7_75t_SL g2491 ( 
.A1(n_2385),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.C(n_87),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2385),
.B(n_84),
.Y(n_2492)
);

AOI221xp5_ASAP7_75t_L g2493 ( 
.A1(n_2385),
.A2(n_89),
.B1(n_86),
.B2(n_88),
.C(n_90),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2348),
.B(n_88),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2348),
.B(n_89),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2348),
.B(n_91),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2348),
.B(n_92),
.Y(n_2497)
);

OAI21xp33_ASAP7_75t_L g2498 ( 
.A1(n_2389),
.A2(n_92),
.B(n_93),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2348),
.B(n_93),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2385),
.B(n_94),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2348),
.B(n_94),
.Y(n_2501)
);

NAND3xp33_ASAP7_75t_L g2502 ( 
.A(n_2385),
.B(n_95),
.C(n_97),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2348),
.B(n_95),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2365),
.B(n_98),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2385),
.B(n_98),
.C(n_99),
.Y(n_2505)
);

INVxp67_ASAP7_75t_L g2506 ( 
.A(n_2404),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2348),
.B(n_100),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2348),
.B(n_100),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2348),
.B(n_102),
.Y(n_2509)
);

OAI221xp5_ASAP7_75t_SL g2510 ( 
.A1(n_2383),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.C(n_106),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2385),
.B(n_105),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2348),
.B(n_106),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2365),
.B(n_107),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2348),
.B(n_107),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2385),
.B(n_108),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2348),
.B(n_108),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2348),
.B(n_109),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2348),
.B(n_109),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2348),
.B(n_110),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2348),
.B(n_112),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2348),
.B(n_113),
.Y(n_2521)
);

OAI21xp5_ASAP7_75t_SL g2522 ( 
.A1(n_2389),
.A2(n_113),
.B(n_114),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2348),
.B(n_115),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_SL g2524 ( 
.A(n_2386),
.B(n_115),
.C(n_116),
.Y(n_2524)
);

OAI21xp5_ASAP7_75t_SL g2525 ( 
.A1(n_2389),
.A2(n_116),
.B(n_117),
.Y(n_2525)
);

NAND4xp25_ASAP7_75t_L g2526 ( 
.A(n_2386),
.B(n_120),
.C(n_117),
.D(n_119),
.Y(n_2526)
);

NAND2xp33_ASAP7_75t_SL g2527 ( 
.A(n_2405),
.B(n_120),
.Y(n_2527)
);

OAI221xp5_ASAP7_75t_L g2528 ( 
.A1(n_2385),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_124),
.Y(n_2528)
);

OAI221xp5_ASAP7_75t_SL g2529 ( 
.A1(n_2383),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_125),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2348),
.B(n_126),
.Y(n_2530)
);

NAND3xp33_ASAP7_75t_L g2531 ( 
.A(n_2385),
.B(n_126),
.C(n_127),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2348),
.B(n_128),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2421),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2468),
.B(n_128),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2426),
.B(n_129),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2426),
.B(n_2506),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_2444),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2489),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2475),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2469),
.B(n_131),
.Y(n_2540)
);

NAND3xp33_ASAP7_75t_L g2541 ( 
.A(n_2447),
.B(n_132),
.C(n_133),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2465),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2470),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2420),
.B(n_132),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2428),
.B(n_134),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2471),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2466),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_2445),
.B(n_134),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2431),
.B(n_136),
.Y(n_2549)
);

HB1xp67_ASAP7_75t_L g2550 ( 
.A(n_2481),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2485),
.B(n_136),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2490),
.B(n_137),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2456),
.Y(n_2553)
);

NAND2x1p5_ASAP7_75t_L g2554 ( 
.A(n_2438),
.B(n_137),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2499),
.B(n_138),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2460),
.B(n_138),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2473),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2427),
.B(n_139),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2501),
.B(n_2507),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2441),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2514),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2476),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2516),
.B(n_139),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2477),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2418),
.B(n_140),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2517),
.B(n_141),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2518),
.B(n_142),
.Y(n_2567)
);

INVx3_ASAP7_75t_L g2568 ( 
.A(n_2519),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2474),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2419),
.B(n_143),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2520),
.B(n_145),
.Y(n_2571)
);

OR2x2_ASAP7_75t_L g2572 ( 
.A(n_2483),
.B(n_146),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2436),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2452),
.B(n_146),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2454),
.B(n_147),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2440),
.Y(n_2576)
);

OR2x2_ASAP7_75t_L g2577 ( 
.A(n_2486),
.B(n_147),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2448),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2435),
.Y(n_2579)
);

OAI221xp5_ASAP7_75t_L g2580 ( 
.A1(n_2484),
.A2(n_151),
.B1(n_148),
.B2(n_150),
.C(n_152),
.Y(n_2580)
);

NAND2x1_ASAP7_75t_SL g2581 ( 
.A(n_2467),
.B(n_148),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2521),
.B(n_154),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2478),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2523),
.B(n_2532),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2459),
.B(n_154),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2494),
.B(n_155),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2495),
.B(n_2496),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2497),
.B(n_155),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2503),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2508),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2509),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2512),
.Y(n_2592)
);

OAI21xp5_ASAP7_75t_SL g2593 ( 
.A1(n_2462),
.A2(n_156),
.B(n_157),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2530),
.B(n_156),
.Y(n_2594)
);

INVx1_ASAP7_75t_SL g2595 ( 
.A(n_2450),
.Y(n_2595)
);

AND2x4_ASAP7_75t_SL g2596 ( 
.A(n_2443),
.B(n_157),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2423),
.B(n_158),
.Y(n_2597)
);

AND2x4_ASAP7_75t_SL g2598 ( 
.A(n_2457),
.B(n_2425),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2429),
.B(n_159),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2430),
.B(n_159),
.Y(n_2600)
);

INVxp67_ASAP7_75t_SL g2601 ( 
.A(n_2439),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2432),
.B(n_2433),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2464),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2504),
.B(n_160),
.Y(n_2604)
);

OR2x2_ASAP7_75t_L g2605 ( 
.A(n_2424),
.B(n_161),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2439),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2422),
.B(n_161),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2513),
.B(n_162),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2492),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2491),
.B(n_162),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2498),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2500),
.B(n_163),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2522),
.B(n_164),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2511),
.B(n_165),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2502),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2451),
.B(n_2463),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2515),
.B(n_166),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2449),
.B(n_167),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2525),
.B(n_167),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2488),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2455),
.B(n_168),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2524),
.B(n_168),
.Y(n_2622)
);

NAND2x1p5_ASAP7_75t_L g2623 ( 
.A(n_2527),
.B(n_169),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_SL g2624 ( 
.A1(n_2505),
.A2(n_169),
.B(n_170),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2531),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2437),
.B(n_171),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2528),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2482),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2526),
.B(n_171),
.Y(n_2629)
);

AND2x4_ASAP7_75t_L g2630 ( 
.A(n_2458),
.B(n_172),
.Y(n_2630)
);

INVxp67_ASAP7_75t_L g2631 ( 
.A(n_2487),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2461),
.B(n_172),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2493),
.B(n_173),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2453),
.B(n_174),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2472),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2442),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2480),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2434),
.B(n_175),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2510),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2529),
.B(n_176),
.Y(n_2640)
);

OR2x2_ASAP7_75t_L g2641 ( 
.A(n_2446),
.B(n_177),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2479),
.B(n_178),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2420),
.B(n_178),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2468),
.B(n_179),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2420),
.B(n_179),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2468),
.B(n_180),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2420),
.B(n_180),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2420),
.B(n_181),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2468),
.B(n_181),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2468),
.B(n_182),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2468),
.B(n_182),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2420),
.B(n_183),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2421),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2421),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2468),
.B(n_183),
.Y(n_2655)
);

BUFx2_ASAP7_75t_L g2656 ( 
.A(n_2468),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2489),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2468),
.B(n_184),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2421),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2421),
.Y(n_2660)
);

BUFx2_ASAP7_75t_L g2661 ( 
.A(n_2468),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2420),
.B(n_185),
.Y(n_2662)
);

INVxp67_ASAP7_75t_SL g2663 ( 
.A(n_2481),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2468),
.B(n_185),
.Y(n_2664)
);

NAND3xp33_ASAP7_75t_L g2665 ( 
.A(n_2447),
.B(n_186),
.C(n_187),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2506),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2468),
.B(n_188),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2468),
.B(n_189),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2468),
.B(n_190),
.Y(n_2669)
);

OR2x2_ASAP7_75t_L g2670 ( 
.A(n_2603),
.B(n_190),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2533),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2653),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2656),
.B(n_191),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2656),
.B(n_192),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2661),
.B(n_194),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2663),
.B(n_195),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2654),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2661),
.B(n_195),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2550),
.B(n_196),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2659),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2579),
.B(n_196),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2536),
.B(n_197),
.Y(n_2682)
);

INVx2_ASAP7_75t_SL g2683 ( 
.A(n_2650),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2666),
.B(n_198),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2553),
.B(n_198),
.Y(n_2685)
);

NAND2x1_ASAP7_75t_L g2686 ( 
.A(n_2568),
.B(n_199),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2560),
.B(n_199),
.Y(n_2687)
);

NOR2xp67_ASAP7_75t_L g2688 ( 
.A(n_2537),
.B(n_200),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2660),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2542),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2559),
.B(n_200),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2595),
.B(n_201),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2547),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2561),
.B(n_201),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2557),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2602),
.B(n_202),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2589),
.B(n_204),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2590),
.B(n_204),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2538),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2562),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2657),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_2573),
.B(n_205),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2546),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2591),
.B(n_205),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2576),
.B(n_206),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2606),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2578),
.B(n_2564),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2592),
.B(n_207),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2543),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2587),
.B(n_208),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2544),
.B(n_210),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2609),
.B(n_210),
.Y(n_2712)
);

CKINVDCx16_ASAP7_75t_R g2713 ( 
.A(n_2658),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2584),
.B(n_211),
.Y(n_2714)
);

HB1xp67_ASAP7_75t_L g2715 ( 
.A(n_2615),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2643),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2534),
.B(n_211),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2625),
.B(n_212),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2644),
.B(n_213),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2645),
.B(n_213),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2646),
.B(n_2649),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2647),
.B(n_214),
.Y(n_2722)
);

AND2x4_ASAP7_75t_L g2723 ( 
.A(n_2583),
.B(n_214),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2648),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2652),
.B(n_2569),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2662),
.B(n_215),
.Y(n_2726)
);

AOI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2593),
.A2(n_218),
.B1(n_215),
.B2(n_217),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2554),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2651),
.B(n_219),
.Y(n_2729)
);

OR2x2_ASAP7_75t_L g2730 ( 
.A(n_2605),
.B(n_219),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2607),
.B(n_220),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2601),
.B(n_220),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2540),
.B(n_221),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2655),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2668),
.B(n_221),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2558),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2598),
.B(n_2631),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2627),
.B(n_222),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2570),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2535),
.B(n_222),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2572),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2637),
.B(n_223),
.Y(n_2742)
);

NOR2xp67_ASAP7_75t_L g2743 ( 
.A(n_2541),
.B(n_224),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2669),
.B(n_224),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2577),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2664),
.B(n_225),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2667),
.B(n_225),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2586),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2597),
.Y(n_2749)
);

AND2x4_ASAP7_75t_SL g2750 ( 
.A(n_2545),
.B(n_226),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2600),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2556),
.Y(n_2752)
);

INVxp67_ASAP7_75t_L g2753 ( 
.A(n_2639),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2599),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2574),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2551),
.B(n_226),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2575),
.Y(n_2757)
);

HB1xp67_ASAP7_75t_L g2758 ( 
.A(n_2552),
.Y(n_2758)
);

INVxp67_ASAP7_75t_SL g2759 ( 
.A(n_2581),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2555),
.B(n_227),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2588),
.B(n_2594),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2563),
.B(n_227),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2566),
.B(n_2567),
.Y(n_2763)
);

INVxp67_ASAP7_75t_SL g2764 ( 
.A(n_2548),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2571),
.B(n_228),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2582),
.B(n_228),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2610),
.Y(n_2767)
);

OR2x2_ASAP7_75t_L g2768 ( 
.A(n_2613),
.B(n_229),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2585),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2549),
.B(n_230),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2621),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2619),
.B(n_230),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2640),
.B(n_231),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2612),
.B(n_231),
.Y(n_2774)
);

BUFx2_ASAP7_75t_L g2775 ( 
.A(n_2614),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2629),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_R g2777 ( 
.A(n_2622),
.B(n_233),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2596),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2617),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2628),
.B(n_234),
.Y(n_2780)
);

NOR2x1p5_ASAP7_75t_L g2781 ( 
.A(n_2665),
.B(n_234),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2626),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2633),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2604),
.B(n_235),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2620),
.B(n_235),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2565),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2608),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2623),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2618),
.B(n_236),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2641),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2638),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_L g2792 ( 
.A(n_2616),
.B(n_236),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2635),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2539),
.B(n_237),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2632),
.B(n_237),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2630),
.B(n_238),
.Y(n_2796)
);

INVx4_ASAP7_75t_L g2797 ( 
.A(n_2634),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2580),
.B(n_239),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2624),
.B(n_239),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2636),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2642),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2611),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2533),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2656),
.B(n_240),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2533),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2603),
.B(n_240),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2656),
.B(n_241),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2533),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2663),
.B(n_242),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2663),
.B(n_242),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2533),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2663),
.B(n_243),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2533),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2560),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2603),
.B(n_243),
.Y(n_2815)
);

OR2x2_ASAP7_75t_L g2816 ( 
.A(n_2603),
.B(n_244),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2656),
.B(n_244),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2656),
.B(n_245),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2663),
.B(n_245),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2656),
.B(n_246),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2656),
.B(n_247),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2603),
.B(n_247),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2663),
.B(n_248),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2663),
.B(n_248),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2560),
.Y(n_2825)
);

OR2x2_ASAP7_75t_L g2826 ( 
.A(n_2603),
.B(n_249),
.Y(n_2826)
);

NAND2xp67_ASAP7_75t_SL g2827 ( 
.A(n_2536),
.B(n_249),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2560),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2663),
.B(n_250),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2663),
.B(n_250),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2656),
.B(n_251),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2656),
.B(n_251),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2656),
.B(n_252),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2533),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2533),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2656),
.B(n_252),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2533),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2533),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2603),
.B(n_253),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2560),
.Y(n_2840)
);

INVx2_ASAP7_75t_SL g2841 ( 
.A(n_2650),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2663),
.B(n_253),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2533),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2663),
.B(n_254),
.Y(n_2844)
);

OR2x2_ASAP7_75t_L g2845 ( 
.A(n_2603),
.B(n_254),
.Y(n_2845)
);

AND2x4_ASAP7_75t_L g2846 ( 
.A(n_2656),
.B(n_255),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2663),
.B(n_255),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2656),
.B(n_256),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2663),
.B(n_256),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2656),
.B(n_257),
.Y(n_2850)
);

INVxp67_ASAP7_75t_L g2851 ( 
.A(n_2656),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2560),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2663),
.B(n_257),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2656),
.B(n_258),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2533),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2663),
.B(n_258),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2663),
.B(n_259),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2663),
.B(n_259),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2656),
.B(n_260),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2656),
.B(n_260),
.Y(n_2860)
);

OR2x2_ASAP7_75t_L g2861 ( 
.A(n_2603),
.B(n_261),
.Y(n_2861)
);

OR2x2_ASAP7_75t_L g2862 ( 
.A(n_2603),
.B(n_261),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2758),
.B(n_2721),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2775),
.B(n_262),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2713),
.B(n_262),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2767),
.B(n_263),
.Y(n_2866)
);

OAI32xp33_ASAP7_75t_L g2867 ( 
.A1(n_2715),
.A2(n_265),
.A3(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2775),
.B(n_265),
.Y(n_2868)
);

AOI211xp5_ASAP7_75t_L g2869 ( 
.A1(n_2798),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_2869)
);

OAI211xp5_ASAP7_75t_L g2870 ( 
.A1(n_2727),
.A2(n_271),
.B(n_268),
.C(n_269),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2814),
.B(n_271),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2753),
.B(n_272),
.Y(n_2872)
);

NAND2x1p5_ASAP7_75t_L g2873 ( 
.A(n_2686),
.B(n_272),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2801),
.B(n_273),
.Y(n_2874)
);

OAI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2764),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2875)
);

XNOR2xp5_ASAP7_75t_L g2876 ( 
.A(n_2763),
.B(n_275),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2707),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2825),
.B(n_276),
.Y(n_2878)
);

OAI211xp5_ASAP7_75t_L g2879 ( 
.A1(n_2851),
.A2(n_281),
.B(n_277),
.C(n_280),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2706),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2828),
.B(n_277),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2734),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2671),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2761),
.B(n_280),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2736),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_2885)
);

OR2x2_ASAP7_75t_L g2886 ( 
.A(n_2752),
.B(n_2716),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2724),
.B(n_282),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2769),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2739),
.B(n_284),
.Y(n_2889)
);

NAND4xp75_ASAP7_75t_L g2890 ( 
.A(n_2743),
.B(n_287),
.C(n_285),
.D(n_286),
.Y(n_2890)
);

NAND4xp75_ASAP7_75t_SL g2891 ( 
.A(n_2674),
.B(n_287),
.C(n_285),
.D(n_286),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2672),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2725),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2677),
.Y(n_2894)
);

INVx3_ASAP7_75t_L g2895 ( 
.A(n_2778),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2680),
.Y(n_2896)
);

AOI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2802),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2725),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2689),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2690),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2803),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2776),
.A2(n_2759),
.B1(n_2783),
.B2(n_2781),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2797),
.Y(n_2903)
);

O2A1O1Ixp33_ASAP7_75t_L g2904 ( 
.A1(n_2676),
.A2(n_291),
.B(n_288),
.C(n_289),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2741),
.B(n_291),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2805),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2787),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2745),
.B(n_292),
.Y(n_2908)
);

AOI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2782),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2673),
.Y(n_2910)
);

INVxp67_ASAP7_75t_L g2911 ( 
.A(n_2737),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2840),
.B(n_2852),
.Y(n_2912)
);

OAI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2688),
.A2(n_302),
.B1(n_312),
.B2(n_293),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2748),
.B(n_295),
.Y(n_2914)
);

NAND2x1p5_ASAP7_75t_L g2915 ( 
.A(n_2846),
.B(n_2860),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2771),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2916)
);

AOI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2790),
.A2(n_300),
.B1(n_297),
.B2(n_299),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2808),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2811),
.Y(n_2919)
);

AOI221xp5_ASAP7_75t_L g2920 ( 
.A1(n_2800),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.C(n_303),
.Y(n_2920)
);

NOR4xp25_ASAP7_75t_L g2921 ( 
.A(n_2718),
.B(n_304),
.C(n_301),
.D(n_303),
.Y(n_2921)
);

NAND4xp75_ASAP7_75t_L g2922 ( 
.A(n_2799),
.B(n_307),
.C(n_305),
.D(n_306),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2675),
.B(n_305),
.Y(n_2923)
);

OR2x2_ASAP7_75t_L g2924 ( 
.A(n_2754),
.B(n_307),
.Y(n_2924)
);

HB1xp67_ASAP7_75t_L g2925 ( 
.A(n_2791),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2788),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2813),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2834),
.Y(n_2928)
);

OAI31xp33_ASAP7_75t_L g2929 ( 
.A1(n_2692),
.A2(n_312),
.A3(n_308),
.B(n_309),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2835),
.Y(n_2930)
);

NAND4xp75_ASAP7_75t_L g2931 ( 
.A(n_2794),
.B(n_313),
.C(n_308),
.D(n_309),
.Y(n_2931)
);

OA222x2_ASAP7_75t_L g2932 ( 
.A1(n_2684),
.A2(n_315),
.B1(n_317),
.B2(n_313),
.C1(n_314),
.C2(n_316),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2837),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2749),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2934)
);

OAI21xp33_ASAP7_75t_L g2935 ( 
.A1(n_2731),
.A2(n_318),
.B(n_320),
.Y(n_2935)
);

OAI33xp33_ASAP7_75t_L g2936 ( 
.A1(n_2695),
.A2(n_322),
.A3(n_324),
.B1(n_320),
.B2(n_321),
.B3(n_323),
.Y(n_2936)
);

AOI32xp33_ASAP7_75t_L g2937 ( 
.A1(n_2795),
.A2(n_325),
.A3(n_327),
.B1(n_322),
.B2(n_326),
.Y(n_2937)
);

OAI221xp5_ASAP7_75t_L g2938 ( 
.A1(n_2730),
.A2(n_2773),
.B1(n_2732),
.B2(n_2810),
.C(n_2809),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2683),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2779),
.Y(n_2940)
);

AOI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2786),
.A2(n_328),
.B1(n_321),
.B2(n_325),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2678),
.B(n_328),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2841),
.B(n_329),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2804),
.B(n_2807),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2817),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2818),
.B(n_329),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2820),
.B(n_330),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2838),
.Y(n_2948)
);

INVxp67_ASAP7_75t_L g2949 ( 
.A(n_2821),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2831),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2843),
.Y(n_2951)
);

NOR2xp33_ASAP7_75t_L g2952 ( 
.A(n_2755),
.B(n_330),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2855),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2832),
.B(n_331),
.Y(n_2954)
);

OAI33xp33_ASAP7_75t_L g2955 ( 
.A1(n_2700),
.A2(n_335),
.A3(n_337),
.B1(n_331),
.B2(n_334),
.B3(n_336),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2812),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2819),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2833),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2823),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2836),
.Y(n_2960)
);

AOI22xp5_ASAP7_75t_L g2961 ( 
.A1(n_2751),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2848),
.B(n_337),
.Y(n_2962)
);

O2A1O1Ixp5_ASAP7_75t_R g2963 ( 
.A1(n_2772),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2757),
.A2(n_343),
.B1(n_339),
.B2(n_341),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2824),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2850),
.B(n_341),
.Y(n_2966)
);

OAI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2854),
.A2(n_343),
.B(n_344),
.Y(n_2967)
);

HB1xp67_ASAP7_75t_L g2968 ( 
.A(n_2859),
.Y(n_2968)
);

OR2x2_ASAP7_75t_L g2969 ( 
.A(n_2709),
.B(n_345),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2691),
.B(n_2682),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2793),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_2971)
);

AOI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2789),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2728),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2702),
.B(n_349),
.Y(n_2974)
);

OR2x2_ASAP7_75t_L g2975 ( 
.A(n_2670),
.B(n_350),
.Y(n_2975)
);

OR3x2_ASAP7_75t_L g2976 ( 
.A(n_2768),
.B(n_352),
.C(n_353),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2687),
.B(n_2694),
.Y(n_2977)
);

INVxp67_ASAP7_75t_L g2978 ( 
.A(n_2806),
.Y(n_2978)
);

NAND4xp25_ASAP7_75t_L g2979 ( 
.A(n_2681),
.B(n_355),
.C(n_352),
.D(n_353),
.Y(n_2979)
);

OAI32xp33_ASAP7_75t_L g2980 ( 
.A1(n_2829),
.A2(n_357),
.A3(n_355),
.B1(n_356),
.B2(n_358),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2714),
.B(n_356),
.Y(n_2981)
);

AOI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2703),
.A2(n_2697),
.B1(n_2704),
.B2(n_2698),
.Y(n_2982)
);

OAI221xp5_ASAP7_75t_L g2983 ( 
.A1(n_2830),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.C(n_361),
.Y(n_2983)
);

XOR2x2_ASAP7_75t_L g2984 ( 
.A(n_2785),
.B(n_361),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2842),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2844),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2847),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2696),
.B(n_360),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2723),
.B(n_362),
.Y(n_2989)
);

INVx2_ASAP7_75t_SL g2990 ( 
.A(n_2750),
.Y(n_2990)
);

NAND4xp75_ASAP7_75t_L g2991 ( 
.A(n_2784),
.B(n_364),
.C(n_362),
.D(n_363),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2708),
.B(n_364),
.Y(n_2992)
);

NOR3xp33_ASAP7_75t_SL g2993 ( 
.A(n_2733),
.B(n_366),
.C(n_367),
.Y(n_2993)
);

NOR4xp25_ASAP7_75t_L g2994 ( 
.A(n_2738),
.B(n_369),
.C(n_367),
.D(n_368),
.Y(n_2994)
);

AOI32xp33_ASAP7_75t_L g2995 ( 
.A1(n_2849),
.A2(n_371),
.A3(n_373),
.B1(n_370),
.B2(n_372),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2780),
.A2(n_372),
.B1(n_368),
.B2(n_370),
.Y(n_2996)
);

INVx2_ASAP7_75t_SL g2997 ( 
.A(n_2740),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2853),
.Y(n_2998)
);

INVxp67_ASAP7_75t_L g2999 ( 
.A(n_2815),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2712),
.B(n_373),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2856),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2717),
.B(n_374),
.Y(n_3002)
);

HB1xp67_ASAP7_75t_L g3003 ( 
.A(n_2685),
.Y(n_3003)
);

AND2x2_ASAP7_75t_SL g3004 ( 
.A(n_2963),
.B(n_2719),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2864),
.Y(n_3005)
);

OAI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2902),
.A2(n_2857),
.B1(n_2858),
.B2(n_2679),
.Y(n_3006)
);

NAND2x1_ASAP7_75t_L g3007 ( 
.A(n_2895),
.B(n_2729),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2863),
.B(n_2735),
.Y(n_3008)
);

O2A1O1Ixp33_ASAP7_75t_L g3009 ( 
.A1(n_2869),
.A2(n_2904),
.B(n_2974),
.C(n_2994),
.Y(n_3009)
);

OR2x2_ASAP7_75t_L g3010 ( 
.A(n_2968),
.B(n_2705),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2886),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_SL g3012 ( 
.A(n_2865),
.B(n_2744),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2868),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2880),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2911),
.B(n_2711),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2864),
.B(n_2770),
.Y(n_3016)
);

AND3x2_ASAP7_75t_L g3017 ( 
.A(n_2921),
.B(n_2760),
.C(n_2756),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2883),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2970),
.B(n_2945),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2892),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2894),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2949),
.B(n_2762),
.Y(n_3022)
);

HB1xp67_ASAP7_75t_L g3023 ( 
.A(n_2925),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2896),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2899),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2977),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2900),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2901),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2950),
.B(n_2816),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2938),
.B(n_2722),
.Y(n_3030)
);

INVxp67_ASAP7_75t_SL g3031 ( 
.A(n_2876),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2958),
.B(n_2822),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2960),
.B(n_2826),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2903),
.B(n_2912),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_3003),
.B(n_2839),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2939),
.B(n_2765),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2977),
.B(n_2845),
.Y(n_3037)
);

AND2x4_ASAP7_75t_L g3038 ( 
.A(n_2910),
.B(n_2710),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2906),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_SL g3040 ( 
.A1(n_2952),
.A2(n_2796),
.B1(n_2774),
.B2(n_2792),
.Y(n_3040)
);

INVx2_ASAP7_75t_SL g3041 ( 
.A(n_2915),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2918),
.Y(n_3042)
);

AOI211xp5_ASAP7_75t_L g3043 ( 
.A1(n_2879),
.A2(n_2777),
.B(n_2720),
.C(n_2726),
.Y(n_3043)
);

OAI22xp33_ASAP7_75t_L g3044 ( 
.A1(n_2982),
.A2(n_2862),
.B1(n_2861),
.B2(n_2742),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2943),
.Y(n_3045)
);

OAI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2993),
.A2(n_2766),
.B(n_2747),
.Y(n_3046)
);

AND3x2_ASAP7_75t_L g3047 ( 
.A(n_2929),
.B(n_2746),
.C(n_2827),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2919),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2907),
.B(n_2693),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2927),
.Y(n_3050)
);

OR2x2_ASAP7_75t_L g3051 ( 
.A(n_2940),
.B(n_2699),
.Y(n_3051)
);

O2A1O1Ixp33_ASAP7_75t_L g3052 ( 
.A1(n_2967),
.A2(n_2701),
.B(n_378),
.C(n_375),
.Y(n_3052)
);

INVxp67_ASAP7_75t_L g3053 ( 
.A(n_2884),
.Y(n_3053)
);

INVx2_ASAP7_75t_SL g3054 ( 
.A(n_2943),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2990),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2978),
.B(n_377),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2944),
.B(n_2997),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_2956),
.B(n_377),
.Y(n_3058)
);

OAI22xp5_ASAP7_75t_L g3059 ( 
.A1(n_2976),
.A2(n_2866),
.B1(n_3001),
.B2(n_2959),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2999),
.B(n_379),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2928),
.Y(n_3061)
);

INVx1_ASAP7_75t_SL g3062 ( 
.A(n_3002),
.Y(n_3062)
);

OR2x2_ASAP7_75t_L g3063 ( 
.A(n_2957),
.B(n_379),
.Y(n_3063)
);

XOR2xp5_ASAP7_75t_L g3064 ( 
.A(n_2891),
.B(n_380),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2887),
.B(n_380),
.Y(n_3065)
);

OR2x2_ASAP7_75t_L g3066 ( 
.A(n_2965),
.B(n_381),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_2924),
.B(n_2979),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2930),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2871),
.B(n_381),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2969),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2893),
.Y(n_3071)
);

AND2x4_ASAP7_75t_L g3072 ( 
.A(n_2878),
.B(n_382),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2933),
.Y(n_3073)
);

OR2x2_ASAP7_75t_L g3074 ( 
.A(n_2985),
.B(n_383),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2986),
.B(n_384),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2987),
.B(n_384),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2948),
.Y(n_3077)
);

OAI21xp5_ASAP7_75t_SL g3078 ( 
.A1(n_2995),
.A2(n_385),
.B(n_386),
.Y(n_3078)
);

NAND2xp33_ASAP7_75t_L g3079 ( 
.A(n_2873),
.B(n_385),
.Y(n_3079)
);

INVx1_ASAP7_75t_SL g3080 ( 
.A(n_2923),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2951),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2953),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2998),
.B(n_386),
.Y(n_3083)
);

OR2x2_ASAP7_75t_L g3084 ( 
.A(n_2877),
.B(n_387),
.Y(n_3084)
);

OAI21xp5_ASAP7_75t_SL g3085 ( 
.A1(n_3017),
.A2(n_3047),
.B(n_3078),
.Y(n_3085)
);

INVx2_ASAP7_75t_SL g3086 ( 
.A(n_3016),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_3016),
.Y(n_3087)
);

OAI21xp33_ASAP7_75t_L g3088 ( 
.A1(n_3055),
.A2(n_2898),
.B(n_2874),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3023),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_3004),
.B(n_2882),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3056),
.Y(n_3091)
);

OR2x2_ASAP7_75t_L g3092 ( 
.A(n_3062),
.B(n_2888),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_3080),
.B(n_2937),
.Y(n_3093)
);

OAI211xp5_ASAP7_75t_SL g3094 ( 
.A1(n_3009),
.A2(n_2983),
.B(n_2935),
.C(n_2972),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_3060),
.Y(n_3095)
);

NOR2xp67_ASAP7_75t_L g3096 ( 
.A(n_3045),
.B(n_2926),
.Y(n_3096)
);

INVx1_ASAP7_75t_SL g3097 ( 
.A(n_3036),
.Y(n_3097)
);

INVxp67_ASAP7_75t_L g3098 ( 
.A(n_3012),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3011),
.Y(n_3099)
);

AOI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_3067),
.A2(n_2955),
.B1(n_2936),
.B2(n_2984),
.Y(n_3100)
);

AOI222xp33_ASAP7_75t_L g3101 ( 
.A1(n_3030),
.A2(n_2885),
.B1(n_2875),
.B2(n_2920),
.C1(n_2870),
.C2(n_2913),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_3008),
.B(n_2881),
.Y(n_3102)
);

AOI21xp33_ASAP7_75t_SL g3103 ( 
.A1(n_3041),
.A2(n_2947),
.B(n_2946),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_3054),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3058),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_3063),
.Y(n_3106)
);

NOR2x1_ASAP7_75t_L g3107 ( 
.A(n_3075),
.B(n_2962),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_3059),
.A2(n_3031),
.B1(n_3006),
.B2(n_3065),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_3070),
.A2(n_2973),
.B1(n_2905),
.B2(n_2908),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_3044),
.A2(n_2890),
.B1(n_2922),
.B2(n_2897),
.Y(n_3110)
);

OAI221xp5_ASAP7_75t_L g3111 ( 
.A1(n_3052),
.A2(n_2996),
.B1(n_2917),
.B2(n_2909),
.C(n_2941),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3066),
.Y(n_3112)
);

HB1xp67_ASAP7_75t_L g3113 ( 
.A(n_3026),
.Y(n_3113)
);

AOI222xp33_ASAP7_75t_L g3114 ( 
.A1(n_3035),
.A2(n_2914),
.B1(n_2889),
.B2(n_2980),
.C1(n_2872),
.C2(n_2867),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_3053),
.B(n_2988),
.Y(n_3115)
);

O2A1O1Ixp33_ASAP7_75t_L g3116 ( 
.A1(n_3043),
.A2(n_2966),
.B(n_2975),
.C(n_2932),
.Y(n_3116)
);

OAI21xp33_ASAP7_75t_SL g3117 ( 
.A1(n_3019),
.A2(n_2954),
.B(n_2942),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3074),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3018),
.Y(n_3119)
);

INVxp67_ASAP7_75t_L g3120 ( 
.A(n_3015),
.Y(n_3120)
);

OAI221xp5_ASAP7_75t_L g3121 ( 
.A1(n_3079),
.A2(n_2916),
.B1(n_2964),
.B2(n_2934),
.C(n_2961),
.Y(n_3121)
);

AND2x4_ASAP7_75t_L g3122 ( 
.A(n_3038),
.B(n_2981),
.Y(n_3122)
);

OAI221xp5_ASAP7_75t_L g3123 ( 
.A1(n_3046),
.A2(n_2971),
.B1(n_2992),
.B2(n_3000),
.C(n_2989),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_3022),
.Y(n_3124)
);

AOI211xp5_ASAP7_75t_L g3125 ( 
.A1(n_3034),
.A2(n_2931),
.B(n_2991),
.C(n_389),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_3007),
.A2(n_390),
.B1(n_387),
.B2(n_388),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3020),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3021),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_SL g3129 ( 
.A1(n_3040),
.A2(n_391),
.B1(n_388),
.B2(n_390),
.Y(n_3129)
);

AOI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_3037),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_3057),
.Y(n_3131)
);

AOI211x1_ASAP7_75t_L g3132 ( 
.A1(n_3013),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_3132)
);

NOR3xp33_ASAP7_75t_L g3133 ( 
.A(n_3076),
.B(n_394),
.C(n_395),
.Y(n_3133)
);

INVxp67_ASAP7_75t_L g3134 ( 
.A(n_3005),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_3010),
.B(n_395),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_3072),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3024),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_3083),
.A2(n_396),
.B(n_397),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_3084),
.Y(n_3139)
);

NOR2x1_ASAP7_75t_L g3140 ( 
.A(n_3064),
.B(n_397),
.Y(n_3140)
);

AOI22xp33_ASAP7_75t_L g3141 ( 
.A1(n_3071),
.A2(n_399),
.B1(n_396),
.B2(n_398),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_3049),
.B(n_398),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3025),
.Y(n_3143)
);

AOI222xp33_ASAP7_75t_L g3144 ( 
.A1(n_3014),
.A2(n_401),
.B1(n_403),
.B2(n_399),
.C1(n_400),
.C2(n_402),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3113),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_SL g3146 ( 
.A1(n_3090),
.A2(n_3028),
.B1(n_3039),
.B2(n_3027),
.Y(n_3146)
);

OAI222xp33_ASAP7_75t_L g3147 ( 
.A1(n_3116),
.A2(n_3051),
.B1(n_3032),
.B2(n_3033),
.C1(n_3029),
.C2(n_3048),
.Y(n_3147)
);

AOI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_3085),
.A2(n_3069),
.B1(n_3050),
.B2(n_3061),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_3122),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3135),
.Y(n_3150)
);

AND3x2_ASAP7_75t_L g3151 ( 
.A(n_3125),
.B(n_3068),
.C(n_3042),
.Y(n_3151)
);

OAI221xp5_ASAP7_75t_L g3152 ( 
.A1(n_3100),
.A2(n_3081),
.B1(n_3082),
.B2(n_3077),
.C(n_3073),
.Y(n_3152)
);

NOR3xp33_ASAP7_75t_L g3153 ( 
.A(n_3098),
.B(n_402),
.C(n_403),
.Y(n_3153)
);

INVx2_ASAP7_75t_SL g3154 ( 
.A(n_3102),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3089),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3092),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_3129),
.B(n_404),
.Y(n_3157)
);

INVxp67_ASAP7_75t_L g3158 ( 
.A(n_3140),
.Y(n_3158)
);

AOI222xp33_ASAP7_75t_L g3159 ( 
.A1(n_3094),
.A2(n_407),
.B1(n_409),
.B2(n_405),
.C1(n_406),
.C2(n_408),
.Y(n_3159)
);

OAI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_3131),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_3160)
);

OAI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_3097),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_3161)
);

NAND3xp33_ASAP7_75t_L g3162 ( 
.A(n_3108),
.B(n_410),
.C(n_412),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3105),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3086),
.B(n_413),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_3087),
.B(n_413),
.Y(n_3165)
);

AOI22xp5_ASAP7_75t_SL g3166 ( 
.A1(n_3120),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_3138),
.A2(n_416),
.B(n_417),
.Y(n_3167)
);

INVx2_ASAP7_75t_SL g3168 ( 
.A(n_3124),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_3117),
.B(n_417),
.Y(n_3169)
);

OAI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_3111),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3104),
.B(n_418),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_3107),
.A2(n_3139),
.B1(n_3101),
.B2(n_3112),
.Y(n_3172)
);

AOI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_3133),
.A2(n_422),
.B1(n_419),
.B2(n_421),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_3132),
.B(n_3115),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_3099),
.B(n_421),
.Y(n_3175)
);

OAI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_3110),
.A2(n_488),
.B(n_489),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3106),
.B(n_490),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3118),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3088),
.B(n_3126),
.Y(n_3179)
);

OR2x2_ASAP7_75t_L g3180 ( 
.A(n_3093),
.B(n_491),
.Y(n_3180)
);

OAI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_3096),
.A2(n_493),
.B(n_494),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3142),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_3147),
.A2(n_3121),
.B(n_3123),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_3158),
.B(n_3103),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_3146),
.A2(n_3114),
.B(n_3134),
.Y(n_3185)
);

AOI21xp33_ASAP7_75t_L g3186 ( 
.A1(n_3174),
.A2(n_3095),
.B(n_3091),
.Y(n_3186)
);

AOI221xp5_ASAP7_75t_L g3187 ( 
.A1(n_3152),
.A2(n_3109),
.B1(n_3127),
.B2(n_3128),
.C(n_3119),
.Y(n_3187)
);

INVx2_ASAP7_75t_SL g3188 ( 
.A(n_3149),
.Y(n_3188)
);

OAI221xp5_ASAP7_75t_L g3189 ( 
.A1(n_3172),
.A2(n_3144),
.B1(n_3141),
.B2(n_3130),
.C(n_3136),
.Y(n_3189)
);

OAI221xp5_ASAP7_75t_L g3190 ( 
.A1(n_3169),
.A2(n_3143),
.B1(n_3137),
.B2(n_498),
.C(n_496),
.Y(n_3190)
);

INVxp67_ASAP7_75t_SL g3191 ( 
.A(n_3166),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3145),
.Y(n_3192)
);

OAI21xp33_ASAP7_75t_L g3193 ( 
.A1(n_3148),
.A2(n_497),
.B(n_500),
.Y(n_3193)
);

NAND3xp33_ASAP7_75t_L g3194 ( 
.A(n_3151),
.B(n_503),
.C(n_504),
.Y(n_3194)
);

OAI221xp5_ASAP7_75t_L g3195 ( 
.A1(n_3167),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.C(n_508),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3175),
.Y(n_3196)
);

AOI22xp5_ASAP7_75t_L g3197 ( 
.A1(n_3150),
.A2(n_512),
.B1(n_509),
.B2(n_511),
.Y(n_3197)
);

AOI222xp33_ASAP7_75t_L g3198 ( 
.A1(n_3156),
.A2(n_519),
.B1(n_522),
.B2(n_514),
.C1(n_515),
.C2(n_520),
.Y(n_3198)
);

NAND3xp33_ASAP7_75t_L g3199 ( 
.A(n_3159),
.B(n_524),
.C(n_525),
.Y(n_3199)
);

XNOR2xp5_ASAP7_75t_L g3200 ( 
.A(n_3154),
.B(n_526),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3180),
.Y(n_3201)
);

AOI221xp5_ASAP7_75t_L g3202 ( 
.A1(n_3179),
.A2(n_531),
.B1(n_527),
.B2(n_529),
.C(n_532),
.Y(n_3202)
);

OAI21xp33_ASAP7_75t_L g3203 ( 
.A1(n_3168),
.A2(n_534),
.B(n_535),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_3165),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3171),
.B(n_537),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_3164),
.Y(n_3206)
);

OAI21xp5_ASAP7_75t_L g3207 ( 
.A1(n_3162),
.A2(n_538),
.B(n_541),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3153),
.B(n_844),
.Y(n_3208)
);

AOI322xp5_ASAP7_75t_L g3209 ( 
.A1(n_3182),
.A2(n_3163),
.A3(n_3178),
.B1(n_3157),
.B2(n_3173),
.C1(n_3155),
.C2(n_3177),
.Y(n_3209)
);

OAI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_3170),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_3210)
);

AOI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_3176),
.A2(n_549),
.B1(n_546),
.B2(n_547),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_3161),
.A2(n_551),
.B(n_554),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3160),
.B(n_560),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3181),
.Y(n_3214)
);

OAI311xp33_ASAP7_75t_L g3215 ( 
.A1(n_3172),
.A2(n_564),
.A3(n_562),
.B1(n_563),
.C1(n_565),
.Y(n_3215)
);

OR2x2_ASAP7_75t_L g3216 ( 
.A(n_3145),
.B(n_566),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3145),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3145),
.B(n_567),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_3149),
.Y(n_3219)
);

NAND3xp33_ASAP7_75t_L g3220 ( 
.A(n_3185),
.B(n_568),
.C(n_569),
.Y(n_3220)
);

NOR3xp33_ASAP7_75t_L g3221 ( 
.A(n_3194),
.B(n_572),
.C(n_574),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3219),
.Y(n_3222)
);

AO22x2_ASAP7_75t_L g3223 ( 
.A1(n_3183),
.A2(n_579),
.B1(n_576),
.B2(n_577),
.Y(n_3223)
);

OAI211xp5_ASAP7_75t_SL g3224 ( 
.A1(n_3187),
.A2(n_3209),
.B(n_3186),
.C(n_3188),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_3191),
.A2(n_580),
.B(n_584),
.Y(n_3225)
);

AOI211x1_ASAP7_75t_L g3226 ( 
.A1(n_3189),
.A2(n_589),
.B(n_585),
.C(n_588),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3196),
.Y(n_3227)
);

NOR3xp33_ASAP7_75t_L g3228 ( 
.A(n_3184),
.B(n_591),
.C(n_592),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3204),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3206),
.B(n_593),
.Y(n_3230)
);

AOI211xp5_ASAP7_75t_L g3231 ( 
.A1(n_3190),
.A2(n_596),
.B(n_594),
.C(n_595),
.Y(n_3231)
);

OAI222xp33_ASAP7_75t_L g3232 ( 
.A1(n_3214),
.A2(n_599),
.B1(n_602),
.B2(n_597),
.C1(n_598),
.C2(n_600),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3213),
.B(n_604),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3192),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3217),
.Y(n_3235)
);

AOI22xp5_ASAP7_75t_L g3236 ( 
.A1(n_3201),
.A2(n_611),
.B1(n_608),
.B2(n_609),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3216),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3193),
.A2(n_612),
.B(n_613),
.Y(n_3238)
);

NOR3xp33_ASAP7_75t_L g3239 ( 
.A(n_3218),
.B(n_614),
.C(n_615),
.Y(n_3239)
);

AO22x2_ASAP7_75t_L g3240 ( 
.A1(n_3199),
.A2(n_619),
.B1(n_616),
.B2(n_617),
.Y(n_3240)
);

AOI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_3203),
.A2(n_623),
.B1(n_620),
.B2(n_622),
.Y(n_3241)
);

AOI22xp5_ASAP7_75t_L g3242 ( 
.A1(n_3200),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_3242)
);

AO22x2_ASAP7_75t_L g3243 ( 
.A1(n_3210),
.A2(n_631),
.B1(n_627),
.B2(n_630),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3224),
.A2(n_3222),
.B(n_3223),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3229),
.Y(n_3245)
);

OAI211xp5_ASAP7_75t_L g3246 ( 
.A1(n_3227),
.A2(n_3207),
.B(n_3202),
.C(n_3212),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3237),
.B(n_3205),
.Y(n_3247)
);

NOR3xp33_ASAP7_75t_L g3248 ( 
.A(n_3220),
.B(n_3208),
.C(n_3195),
.Y(n_3248)
);

NAND4xp25_ASAP7_75t_L g3249 ( 
.A(n_3234),
.B(n_3211),
.C(n_3198),
.D(n_3197),
.Y(n_3249)
);

NOR2xp67_ASAP7_75t_SL g3250 ( 
.A(n_3233),
.B(n_3215),
.Y(n_3250)
);

OAI221xp5_ASAP7_75t_L g3251 ( 
.A1(n_3225),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.C(n_636),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_3235),
.B(n_637),
.Y(n_3252)
);

OAI211xp5_ASAP7_75t_L g3253 ( 
.A1(n_3226),
.A2(n_642),
.B(n_640),
.C(n_641),
.Y(n_3253)
);

NAND3xp33_ASAP7_75t_SL g3254 ( 
.A(n_3231),
.B(n_644),
.C(n_648),
.Y(n_3254)
);

NOR3xp33_ASAP7_75t_L g3255 ( 
.A(n_3230),
.B(n_649),
.C(n_652),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3247),
.Y(n_3256)
);

CKINVDCx16_ASAP7_75t_R g3257 ( 
.A(n_3245),
.Y(n_3257)
);

NOR2x1_ASAP7_75t_L g3258 ( 
.A(n_3244),
.B(n_3232),
.Y(n_3258)
);

OAI22xp5_ASAP7_75t_L g3259 ( 
.A1(n_3252),
.A2(n_3246),
.B1(n_3240),
.B2(n_3253),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3250),
.B(n_3221),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_3257),
.B(n_3248),
.Y(n_3261)
);

AOI22xp5_ASAP7_75t_L g3262 ( 
.A1(n_3260),
.A2(n_3249),
.B1(n_3255),
.B2(n_3254),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3262),
.B(n_3256),
.Y(n_3263)
);

OR2x2_ASAP7_75t_L g3264 ( 
.A(n_3261),
.B(n_3259),
.Y(n_3264)
);

INVx1_ASAP7_75t_SL g3265 ( 
.A(n_3264),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_3263),
.Y(n_3266)
);

AOI221x1_ASAP7_75t_L g3267 ( 
.A1(n_3263),
.A2(n_3228),
.B1(n_3258),
.B2(n_3239),
.C(n_3238),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3265),
.B(n_3242),
.Y(n_3268)
);

NAND4xp25_ASAP7_75t_SL g3269 ( 
.A(n_3267),
.B(n_3266),
.C(n_3251),
.D(n_3241),
.Y(n_3269)
);

CKINVDCx5p33_ASAP7_75t_R g3270 ( 
.A(n_3266),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3270),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3268),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3272),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3273),
.B(n_3271),
.Y(n_3274)
);

OR3x2_ASAP7_75t_L g3275 ( 
.A(n_3274),
.B(n_3269),
.C(n_3236),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3275),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_3276),
.A2(n_3243),
.B(n_653),
.Y(n_3277)
);

AOI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3277),
.A2(n_841),
.B1(n_658),
.B2(n_655),
.Y(n_3278)
);

AOI221xp5_ASAP7_75t_L g3279 ( 
.A1(n_3278),
.A2(n_660),
.B1(n_657),
.B2(n_659),
.C(n_662),
.Y(n_3279)
);

AOI211xp5_ASAP7_75t_L g3280 ( 
.A1(n_3279),
.A2(n_671),
.B(n_667),
.C(n_669),
.Y(n_3280)
);


endmodule