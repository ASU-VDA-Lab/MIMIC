module fake_jpeg_25883_n_311 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_24),
.B1(n_14),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_51),
.B1(n_22),
.B2(n_19),
.Y(n_95)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_60),
.Y(n_93)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_30),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_68),
.C(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_38),
.B1(n_24),
.B2(n_33),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_73),
.B1(n_46),
.B2(n_49),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_24),
.B1(n_38),
.B2(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_90),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_73),
.Y(n_104)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_89),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_20),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_35),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_68),
.C(n_61),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_102),
.Y(n_132)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_111),
.B(n_117),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_59),
.B1(n_68),
.B2(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_119),
.B1(n_70),
.B2(n_48),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_112),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_68),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_82),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_69),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_58),
.B1(n_47),
.B2(n_66),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_121),
.B1(n_27),
.B2(n_29),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_55),
.B1(n_66),
.B2(n_40),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_58),
.B1(n_70),
.B2(n_42),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_78),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_64),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_84),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_147),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_82),
.C(n_94),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_139),
.C(n_26),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_120),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_131),
.B1(n_138),
.B2(n_145),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_71),
.B1(n_88),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_130),
.B1(n_151),
.B2(n_52),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_88),
.B1(n_96),
.B2(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_96),
.B1(n_70),
.B2(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_98),
.B1(n_107),
.B2(n_122),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_70),
.B1(n_64),
.B2(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_146),
.Y(n_177)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_25),
.B1(n_19),
.B2(n_14),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_114),
.C(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_142),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_97),
.B(n_16),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_148),
.B(n_98),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_25),
.B1(n_64),
.B2(n_16),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_35),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_20),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_25),
.B1(n_16),
.B2(n_39),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_107),
.B1(n_102),
.B2(n_100),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_15),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_15),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_169),
.B(n_176),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_184),
.B1(n_176),
.B2(n_135),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_11),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_160),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_186),
.C(n_148),
.Y(n_202)
);

XOR2x2_ASAP7_75t_SL g162 ( 
.A(n_150),
.B(n_15),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_182),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_102),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_168),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_21),
.B1(n_20),
.B2(n_26),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_26),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_132),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_15),
.B(n_13),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_18),
.B(n_17),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_18),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_39),
.B1(n_17),
.B2(n_18),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_181),
.B1(n_145),
.B2(n_148),
.Y(n_203)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_178),
.Y(n_204)
);

AOI22x1_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_13),
.B1(n_27),
.B2(n_35),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_129),
.A2(n_39),
.B1(n_21),
.B2(n_26),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_124),
.B(n_140),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_139),
.C(n_147),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_199),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_194),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_141),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_174),
.Y(n_214)
);

AO221x1_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_142),
.B1(n_149),
.B2(n_10),
.C(n_11),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g225 ( 
.A(n_198),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_161),
.C(n_186),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_156),
.B1(n_13),
.B2(n_21),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_212),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_182),
.B1(n_162),
.B2(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_21),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_231),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_211),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_221),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_157),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_216),
.B(n_233),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_189),
.C(n_227),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_181),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_207),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_159),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_164),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_214),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_156),
.B(n_173),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_194),
.B1(n_212),
.B2(n_210),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_243),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_203),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.C(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_225),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_1),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_197),
.C(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_199),
.B1(n_197),
.B2(n_188),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_217),
.B1(n_208),
.B2(n_195),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_213),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_222),
.B(n_215),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_258),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_216),
.B(n_218),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_267),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_234),
.B(n_231),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_217),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_265),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_261),
.B1(n_260),
.B2(n_258),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_242),
.C(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_245),
.C(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_237),
.C(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_243),
.C(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.C(n_279),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_1),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_3),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_4),
.C(n_5),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_255),
.B1(n_266),
.B2(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_283),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_255),
.B(n_6),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_4),
.B(n_6),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_4),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_6),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_274),
.B(n_272),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_284),
.B(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_269),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_7),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_7),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_297),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_9),
.C(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_295),
.C(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_303),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_302),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_306),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_304),
.B1(n_301),
.B2(n_9),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_9),
.B(n_192),
.Y(n_311)
);


endmodule