module fake_jpeg_20460_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_68),
.Y(n_110)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_43),
.B(n_42),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_35),
.B1(n_23),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_69),
.B1(n_71),
.B2(n_39),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_35),
.B1(n_23),
.B2(n_28),
.Y(n_69)
);

AO22x2_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g128 ( 
.A(n_73),
.Y(n_128)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_83),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_39),
.B1(n_37),
.B2(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_37),
.B1(n_40),
.B2(n_36),
.Y(n_108)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_84),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_40),
.B(n_36),
.C(n_41),
.Y(n_120)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_17),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_98),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_48),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_35),
.B1(n_40),
.B2(n_36),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_62),
.B1(n_92),
.B2(n_20),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_117),
.B(n_120),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_38),
.C(n_18),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_129),
.C(n_131),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_64),
.A2(n_28),
.B(n_15),
.C(n_23),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_33),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_18),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_131),
.B1(n_84),
.B2(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_66),
.A2(n_39),
.B1(n_36),
.B2(n_41),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_162),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_76),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_143),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_142),
.B(n_146),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_145),
.B1(n_108),
.B2(n_122),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_72),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_151),
.B1(n_133),
.B2(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_77),
.B1(n_78),
.B2(n_70),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_73),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_152),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_41),
.C(n_63),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_75),
.C(n_26),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_20),
.B(n_16),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_107),
.B(n_16),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_18),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_33),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_30),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_32),
.B1(n_15),
.B2(n_16),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_161),
.B1(n_106),
.B2(n_133),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_30),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_30),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_30),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_102),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_132),
.B(n_121),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_164),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_167),
.B1(n_172),
.B2(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_132),
.B1(n_112),
.B2(n_119),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_179),
.B(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_193),
.B1(n_156),
.B2(n_149),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_109),
.B1(n_112),
.B2(n_106),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_109),
.B1(n_123),
.B2(n_119),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_148),
.B1(n_152),
.B2(n_163),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_20),
.B(n_24),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_17),
.B(n_22),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_124),
.B1(n_111),
.B2(n_32),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_186),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_111),
.B1(n_32),
.B2(n_15),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_134),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_192),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_138),
.B1(n_149),
.B2(n_137),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_25),
.B1(n_22),
.B2(n_26),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_27),
.B1(n_24),
.B2(n_17),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_151),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_75),
.C(n_26),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_148),
.C(n_146),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_202),
.B1(n_216),
.B2(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_205),
.C(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_158),
.B1(n_153),
.B2(n_151),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_208),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_175),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

OA21x2_ASAP7_75t_SL g210 ( 
.A1(n_170),
.A2(n_155),
.B(n_143),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_29),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_136),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_217),
.B(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_183),
.B(n_142),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_159),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_219),
.B1(n_221),
.B2(n_181),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_160),
.C(n_94),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_160),
.B1(n_96),
.B2(n_90),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_173),
.A2(n_90),
.B1(n_25),
.B2(n_31),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_179),
.B(n_195),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_224),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_164),
.A3(n_176),
.B1(n_169),
.B2(n_165),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_25),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_188),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_168),
.A2(n_164),
.B(n_196),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_174),
.A2(n_172),
.B1(n_176),
.B2(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_200),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_185),
.B1(n_166),
.B2(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_231),
.A2(n_244),
.B(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_166),
.C(n_31),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_242),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_205),
.C(n_224),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_245),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_7),
.B(n_14),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_203),
.B(n_7),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_31),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_204),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_258),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_206),
.B1(n_214),
.B2(n_200),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_263),
.B1(n_209),
.B2(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_226),
.B1(n_199),
.B2(n_202),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_259),
.B1(n_232),
.B2(n_231),
.Y(n_272)
);

OA22x2_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_206),
.B1(n_210),
.B2(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_265),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_232),
.B1(n_238),
.B2(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_203),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_247),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_267),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_218),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_229),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_229),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_242),
.C(n_233),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_286),
.C(n_258),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_234),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_244),
.B1(n_197),
.B2(n_248),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_217),
.B1(n_8),
.B2(n_9),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_243),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_245),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_6),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_257),
.B1(n_253),
.B2(n_258),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_264),
.B(n_256),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_237),
.C(n_217),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_286),
.B1(n_280),
.B2(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_293),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_264),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_263),
.C(n_268),
.Y(n_293)
);

XOR2x2_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_298),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_249),
.B(n_217),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_6),
.C(n_12),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_281),
.B1(n_279),
.B2(n_273),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_308),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_306),
.B1(n_294),
.B2(n_290),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_282),
.B1(n_275),
.B2(n_3),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_282),
.B1(n_2),
.B2(n_3),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_289),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_314),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_293),
.B(n_298),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_315),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_292),
.B(n_287),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_311),
.Y(n_320)
);

NAND4xp25_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.C(n_317),
.D(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_309),
.C(n_302),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_316),
.C(n_302),
.Y(n_323)
);

AOI321xp33_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_308),
.A3(n_287),
.B1(n_299),
.B2(n_9),
.C(n_11),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_14),
.B(n_10),
.Y(n_325)
);

OAI31xp33_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_8),
.A3(n_10),
.B(n_4),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_1),
.Y(n_327)
);


endmodule