module fake_jpeg_18581_n_37 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx13_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_2),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_2),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

A2O1A1Ixp33_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_1),
.B(n_0),
.C(n_3),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.C(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_3),
.B1(n_13),
.B2(n_10),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_3),
.B1(n_9),
.B2(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_13),
.B(n_8),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_14),
.B(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_19),
.B1(n_7),
.B2(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_23),
.B1(n_28),
.B2(n_30),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_31),
.B(n_23),
.Y(n_36)
);

OAI321xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_26),
.A3(n_22),
.B1(n_27),
.B2(n_28),
.C(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_25),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B1(n_31),
.B2(n_34),
.Y(n_37)
);


endmodule