module fake_jpeg_669_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_62),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_1),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_64),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_54),
.C(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_100),
.Y(n_110)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_71),
.B(n_53),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_70),
.B(n_69),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_68),
.B1(n_72),
.B2(n_57),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_96),
.B1(n_99),
.B2(n_50),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_72),
.B1(n_57),
.B2(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_59),
.B1(n_66),
.B2(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_66),
.B1(n_51),
.B2(n_69),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_70),
.B1(n_65),
.B2(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_50),
.Y(n_112)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_93),
.B1(n_96),
.B2(n_26),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_67),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_109),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_65),
.B1(n_60),
.B2(n_55),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_55),
.B(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_2),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_3),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_3),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_4),
.B(n_6),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_145),
.B1(n_131),
.B2(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_22),
.C(n_43),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_136),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_7),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_21),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_137),
.B1(n_11),
.B2(n_12),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_119),
.C(n_114),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_29),
.B1(n_40),
.B2(n_39),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_10),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_139),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_24),
.C(n_37),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_10),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_159),
.B1(n_128),
.B2(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_153),
.B(n_154),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_30),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_31),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_132),
.B(n_137),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_155),
.B(n_159),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_152),
.B1(n_161),
.B2(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_33),
.C(n_36),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_167),
.C(n_169),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_19),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_32),
.C(n_34),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_167),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_158),
.C(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_166),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_165),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_169),
.Y(n_178)
);

OAI21x1_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_179),
.B(n_175),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_178),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_171),
.B1(n_146),
.B2(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_171),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_47),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_17),
.B(n_18),
.Y(n_186)
);


endmodule