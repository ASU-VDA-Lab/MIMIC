module fake_netlist_6_1867_n_1695 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1695);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1695;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_111),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_36),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_104),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_9),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_39),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_75),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_45),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_69),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_72),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_40),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_85),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_37),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_36),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_5),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_28),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_31),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_67),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_62),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_40),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_38),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_38),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_12),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_17),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_66),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_128),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_102),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_15),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_64),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_9),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_56),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_61),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_132),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_148),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_79),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_115),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_101),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_145),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_120),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_105),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_142),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_71),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_18),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_113),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_8),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_91),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_19),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_114),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_138),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_59),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_19),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_89),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_58),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_65),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_80),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_156),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_25),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_10),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_63),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_29),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_35),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_46),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_86),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_76),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_51),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_153),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_55),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_96),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_134),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_103),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_33),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_108),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_121),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_42),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_13),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_4),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_29),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_146),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_41),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_119),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_39),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_28),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_7),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_0),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_112),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_31),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_51),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_129),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_42),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_55),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_78),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_0),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_161),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_20),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_127),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_54),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_21),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_97),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_53),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_57),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_20),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_160),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_14),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_43),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_25),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_99),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_94),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_151),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_83),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_33),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_11),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_159),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_16),
.Y(n_326)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_47),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_100),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_41),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_207),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_242),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_182),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_210),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_216),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_194),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_218),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_258),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_235),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_221),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_228),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_242),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_229),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_242),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_259),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_217),
.B(n_1),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_230),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_251),
.B(n_2),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_240),
.B(n_3),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_183),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_215),
.B(n_3),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_166),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_168),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_231),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_168),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_232),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_242),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_215),
.B(n_4),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_166),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_236),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_239),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_265),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_243),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_170),
.B(n_6),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_242),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_260),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_189),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_245),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_247),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_189),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_248),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_170),
.B(n_6),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_263),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_320),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_328),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_202),
.B(n_8),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_263),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_263),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_177),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_265),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_263),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_263),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_322),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_172),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_289),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_289),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_325),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_289),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_212),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_328),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_250),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_289),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_289),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_187),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_171),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_265),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_202),
.B(n_219),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_187),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_254),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_166),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_281),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_261),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_191),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_268),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_166),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_224),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_219),
.B(n_256),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_224),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_244),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_244),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_273),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_177),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_209),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_279),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_209),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_341),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_407),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_380),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_167),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_332),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_343),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_343),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_264),
.B1(n_293),
.B2(n_275),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_333),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_359),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

CKINVDCx11_ASAP7_75t_R g437 ( 
.A(n_335),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_334),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_389),
.Y(n_441)
);

BUFx4f_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_390),
.B(n_167),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_373),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_336),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_373),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_338),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_339),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_340),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_401),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_342),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_347),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_354),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_380),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_356),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_351),
.B(n_358),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_345),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_385),
.B(n_169),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_360),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_366),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_355),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_386),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_361),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_363),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_412),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_368),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_371),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_391),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_399),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_402),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_411),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_468),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_452),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_441),
.B(n_350),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_414),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_421),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_441),
.B(n_350),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_459),
.B(n_369),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_468),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_362),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_471),
.B(n_369),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_427),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_452),
.B(n_367),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_461),
.B(n_256),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_461),
.B(n_393),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_432),
.A2(n_257),
.B1(n_277),
.B2(n_270),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_432),
.A2(n_396),
.B1(n_195),
.B2(n_205),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_424),
.B(n_466),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_426),
.B(n_319),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_426),
.B(n_353),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_444),
.B(n_370),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_477),
.Y(n_526)
);

AND2x2_ASAP7_75t_SL g527 ( 
.A(n_424),
.B(n_346),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_477),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_444),
.B(n_319),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_466),
.B(n_396),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_473),
.B(n_166),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_473),
.B(n_393),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_420),
.B(n_197),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_478),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_379),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_440),
.B(n_404),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_450),
.B(n_374),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_428),
.B(n_395),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_476),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_431),
.B(n_370),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_476),
.A2(n_372),
.B1(n_364),
.B2(n_376),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_447),
.B(n_337),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_431),
.B(n_395),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_472),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_435),
.B(n_395),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_478),
.Y(n_551)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_486),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_425),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_435),
.B(n_370),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_438),
.B(n_204),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_456),
.B(n_415),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_475),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_445),
.B(n_288),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_458),
.B(n_415),
.Y(n_561)
);

INVx4_ASAP7_75t_SL g562 ( 
.A(n_425),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_446),
.B(n_276),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_460),
.Y(n_564)
);

OAI21xp33_ASAP7_75t_SL g565 ( 
.A1(n_449),
.A2(n_348),
.B(n_349),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_449),
.B(n_283),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_469),
.B(n_344),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_486),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_474),
.B(n_197),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_479),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_451),
.B(n_173),
.Y(n_574)
);

NAND3x1_ASAP7_75t_L g575 ( 
.A(n_451),
.B(n_246),
.C(n_203),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_436),
.B(n_197),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_480),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_436),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_484),
.B(n_413),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_454),
.B(n_176),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_454),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_485),
.B(n_197),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_436),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_487),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_457),
.B(n_413),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_463),
.Y(n_587)
);

BUFx4f_ASAP7_75t_L g588 ( 
.A(n_436),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_464),
.B(n_410),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_489),
.B(n_197),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_464),
.B(n_394),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_490),
.A2(n_383),
.B1(n_387),
.B2(n_199),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_470),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_483),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_491),
.B(n_384),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_483),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_442),
.A2(n_227),
.B1(n_291),
.B2(n_329),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_436),
.Y(n_598)
);

AND2x4_ASAP7_75t_SL g599 ( 
.A(n_488),
.B(n_206),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_488),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_467),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_467),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_467),
.B(n_394),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_467),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_482),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_482),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_482),
.B(n_200),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_419),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_419),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_419),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_419),
.B(n_208),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_443),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_443),
.B(n_211),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_443),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_443),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_453),
.B(n_403),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_416),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_416),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_429),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_429),
.A2(n_270),
.B1(n_277),
.B2(n_257),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_429),
.B(n_410),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_434),
.B(n_169),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_434),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_453),
.B(n_222),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_434),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_439),
.B(n_398),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_501),
.B(n_223),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_522),
.A2(n_274),
.B1(n_271),
.B2(n_310),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_565),
.A2(n_272),
.B(n_233),
.C(n_234),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_515),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_524),
.B(n_174),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_506),
.B(n_398),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_507),
.B(n_174),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_525),
.B(n_237),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_510),
.B(n_175),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_496),
.B(n_175),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_626),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_626),
.Y(n_641)
);

BUFx4_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_591),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g644 ( 
.A1(n_546),
.A2(n_284),
.B(n_298),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_591),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_513),
.B(n_522),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_525),
.B(n_238),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_534),
.B(n_278),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_510),
.B(n_178),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_618),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_589),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_613),
.B(n_280),
.Y(n_652)
);

AOI221xp5_ASAP7_75t_L g653 ( 
.A1(n_516),
.A2(n_198),
.B1(n_196),
.B2(n_190),
.C(n_188),
.Y(n_653)
);

AND2x6_ASAP7_75t_SL g654 ( 
.A(n_547),
.B(n_285),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_512),
.B(n_262),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_512),
.B(n_282),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_580),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_543),
.B(n_595),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_492),
.B(n_290),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_493),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_603),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_494),
.B(n_296),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_495),
.B(n_301),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_558),
.B(n_297),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_570),
.B(n_180),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_497),
.B(n_304),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_518),
.A2(n_302),
.B1(n_196),
.B2(n_190),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_564),
.B(n_180),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_603),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_499),
.B(n_306),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_498),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_537),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_559),
.A2(n_305),
.B1(n_303),
.B2(n_309),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_500),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_498),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_572),
.B(n_185),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_505),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_572),
.B(n_185),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_502),
.B(n_439),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_583),
.B(n_186),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_500),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_509),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_186),
.Y(n_683)
);

AND2x6_ASAP7_75t_SL g684 ( 
.A(n_538),
.B(n_557),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_603),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_590),
.B(n_192),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_509),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_SL g688 ( 
.A(n_592),
.B(n_198),
.C(n_188),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g689 ( 
.A(n_585),
.B(n_193),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_573),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_586),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_602),
.B(n_262),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_508),
.B(n_523),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_602),
.B(n_262),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_559),
.A2(n_299),
.B1(n_316),
.B2(n_179),
.Y(n_696)
);

AND2x6_ASAP7_75t_SL g697 ( 
.A(n_540),
.B(n_406),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_617),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_617),
.Y(n_699)
);

BUFx12f_ASAP7_75t_L g700 ( 
.A(n_529),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_561),
.B(n_199),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_602),
.B(n_266),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_582),
.B(n_448),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_529),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_619),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_559),
.A2(n_181),
.B1(n_184),
.B2(n_179),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_505),
.Y(n_707)
);

AND2x6_ASAP7_75t_SL g708 ( 
.A(n_559),
.B(n_406),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_503),
.B(n_286),
.C(n_213),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_520),
.A2(n_249),
.B1(n_201),
.B2(n_308),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_517),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_593),
.B(n_266),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_578),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_578),
.B(n_249),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_503),
.B(n_181),
.Y(n_715)
);

OAI221xp5_ASAP7_75t_L g716 ( 
.A1(n_621),
.A2(n_214),
.B1(n_220),
.B2(n_225),
.C(n_226),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_600),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_504),
.B(n_184),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_590),
.B(n_308),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_556),
.B(n_311),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_604),
.B(n_266),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_568),
.B(n_315),
.Y(n_722)
);

AND2x6_ASAP7_75t_L g723 ( 
.A(n_520),
.B(n_266),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_522),
.A2(n_315),
.B1(n_321),
.B2(n_241),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_587),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_527),
.A2(n_295),
.B1(n_292),
.B2(n_326),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_522),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_517),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_563),
.B(n_267),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_587),
.B(n_269),
.Y(n_730)
);

AND2x6_ASAP7_75t_SL g731 ( 
.A(n_541),
.B(n_409),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_619),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_599),
.B(n_287),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_504),
.B(n_314),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_594),
.B(n_409),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_526),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_526),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_604),
.B(n_313),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_599),
.B(n_408),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_513),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_596),
.B(n_408),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_532),
.A2(n_313),
.B(n_324),
.C(n_323),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_326),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_569),
.B(n_324),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_555),
.B(n_323),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_605),
.B(n_606),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_522),
.A2(n_318),
.B1(n_317),
.B2(n_314),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_596),
.B(n_318),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_622),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_601),
.B(n_317),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_623),
.B(n_312),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_527),
.B(n_542),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_530),
.B(n_307),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_548),
.B(n_300),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_575),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_530),
.B(n_550),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_561),
.B(n_295),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_605),
.A2(n_607),
.B(n_606),
.C(n_574),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_607),
.A2(n_294),
.B(n_292),
.C(n_16),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_530),
.B(n_294),
.Y(n_760)
);

INVx5_ASAP7_75t_L g761 ( 
.A(n_530),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_530),
.B(n_163),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_511),
.Y(n_763)
);

AND2x6_ASAP7_75t_SL g764 ( 
.A(n_552),
.B(n_10),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_581),
.A2(n_13),
.B(n_21),
.C(n_22),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_610),
.B(n_60),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_752),
.A2(n_519),
.B1(n_531),
.B2(n_608),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_624),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_758),
.A2(n_521),
.B(n_588),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_763),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_632),
.A2(n_608),
.B1(n_516),
.B2(n_610),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_752),
.A2(n_567),
.B1(n_529),
.B2(n_627),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_SL g773 ( 
.A(n_660),
.B(n_528),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_661),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_640),
.B(n_549),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_632),
.A2(n_516),
.B1(n_610),
.B2(n_624),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_669),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_658),
.B(n_567),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_700),
.Y(n_779)
);

AO21x2_ASAP7_75t_L g780 ( 
.A1(n_756),
.A2(n_612),
.B(n_614),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_628),
.A2(n_567),
.B1(n_627),
.B2(n_516),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_740),
.A2(n_598),
.B(n_521),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_685),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_665),
.A2(n_552),
.B(n_625),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_630),
.A2(n_576),
.B(n_535),
.C(n_551),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_705),
.B(n_619),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_725),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_641),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_705),
.B(n_560),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_674),
.A2(n_575),
.B1(n_616),
.B2(n_615),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_722),
.B(n_514),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_681),
.A2(n_611),
.B1(n_514),
.B2(n_533),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_636),
.B(n_536),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_672),
.Y(n_795)
);

BUFx8_ASAP7_75t_L g796 ( 
.A(n_704),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_657),
.B(n_584),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_634),
.Y(n_798)
);

BUFx2_ASAP7_75t_SL g799 ( 
.A(n_690),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_676),
.A2(n_514),
.B(n_533),
.C(n_579),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_676),
.A2(n_533),
.B(n_579),
.C(n_536),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_SL g802 ( 
.A(n_713),
.B(n_554),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_643),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_732),
.A2(n_646),
.B(n_647),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_749),
.B(n_528),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_633),
.B(n_544),
.Y(n_806)
);

AOI21x1_ASAP7_75t_L g807 ( 
.A1(n_746),
.A2(n_551),
.B(n_553),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_746),
.A2(n_579),
.B(n_571),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_645),
.A2(n_571),
.B1(n_544),
.B2(n_577),
.Y(n_809)
);

AO32x2_ASAP7_75t_L g810 ( 
.A1(n_667),
.A2(n_535),
.A3(n_576),
.B1(n_24),
.B2(n_26),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_739),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_640),
.B(n_562),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_651),
.B(n_577),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_698),
.B(n_22),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_693),
.A2(n_766),
.B(n_656),
.Y(n_815)
);

OAI321xp33_ASAP7_75t_L g816 ( 
.A1(n_743),
.A2(n_23),
.A3(n_24),
.B1(n_26),
.B2(n_27),
.C(n_30),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_671),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_722),
.B(n_566),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_682),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_699),
.B(n_34),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_738),
.A2(n_35),
.B(n_43),
.C(n_44),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_SL g822 ( 
.A1(n_762),
.A2(n_562),
.B(n_47),
.C(n_48),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_717),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_735),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_694),
.B(n_562),
.Y(n_825)
);

NAND2x1p5_ASAP7_75t_L g826 ( 
.A(n_682),
.B(n_609),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_691),
.B(n_609),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_675),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_741),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_715),
.B(n_46),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_664),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_677),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_668),
.B(n_620),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_744),
.B(n_48),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_678),
.A2(n_620),
.B1(n_88),
.B2(n_106),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_678),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_664),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_635),
.B(n_49),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_707),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_718),
.B(n_52),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_753),
.A2(n_107),
.B(n_154),
.Y(n_841)
);

AO32x2_ASAP7_75t_L g842 ( 
.A1(n_710),
.A2(n_54),
.A3(n_56),
.B1(n_59),
.B2(n_68),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_648),
.B(n_74),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_711),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_635),
.B(n_77),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_703),
.A2(n_81),
.B(n_82),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_738),
.A2(n_87),
.B(n_109),
.C(n_110),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_754),
.B(n_133),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_637),
.B(n_140),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_754),
.B(n_147),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_728),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_755),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_757),
.B(n_637),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_745),
.B(n_751),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_682),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_689),
.B(n_682),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_745),
.B(n_736),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_757),
.B(n_649),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_680),
.A2(n_686),
.B1(n_719),
.B2(n_683),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_649),
.A2(n_719),
.B1(n_686),
.B2(n_683),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_650),
.A2(n_737),
.B(n_712),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_760),
.A2(n_750),
.B(n_680),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_759),
.A2(n_765),
.B(n_743),
.C(n_742),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_687),
.B(n_747),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_644),
.A2(n_747),
.B(n_652),
.C(n_733),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_687),
.B(n_706),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_687),
.B(n_670),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_688),
.B(n_748),
.Y(n_868)
);

NAND2x1p5_ASAP7_75t_L g869 ( 
.A(n_761),
.B(n_702),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_655),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_638),
.B(n_733),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_629),
.A2(n_761),
.B1(n_663),
.B2(n_734),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_726),
.A2(n_714),
.B(n_653),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_696),
.A2(n_662),
.B(n_666),
.C(n_659),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_731),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_692),
.A2(n_702),
.B(n_695),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_730),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_SL g878 ( 
.A1(n_692),
.A2(n_695),
.B(n_721),
.C(n_696),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_663),
.A2(n_729),
.B(n_720),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_673),
.B(n_706),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_709),
.A2(n_701),
.B1(n_727),
.B2(n_724),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_755),
.A2(n_673),
.B1(n_716),
.B2(n_664),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_723),
.A2(n_655),
.B(n_708),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_684),
.B(n_697),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_723),
.A2(n_655),
.B(n_714),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_723),
.B(n_655),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_655),
.Y(n_887)
);

NAND2x1p5_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_642),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_654),
.A2(n_746),
.B(n_756),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_764),
.B(n_501),
.Y(n_890)
);

AO21x1_ASAP7_75t_L g891 ( 
.A1(n_628),
.A2(n_632),
.B(n_637),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_746),
.A2(n_756),
.B(n_679),
.Y(n_892)
);

NOR2x1_ASAP7_75t_L g893 ( 
.A(n_704),
.B(n_573),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_632),
.B(n_506),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_632),
.A2(n_501),
.B(n_565),
.C(n_628),
.Y(n_895)
);

AND2x6_ASAP7_75t_L g896 ( 
.A(n_756),
.B(n_631),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_632),
.A2(n_501),
.B(n_565),
.C(n_628),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_633),
.Y(n_898)
);

NOR2xp67_ASAP7_75t_SL g899 ( 
.A(n_705),
.B(n_732),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_658),
.B(n_506),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_682),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_630),
.A2(n_471),
.B(n_510),
.C(n_565),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_661),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_763),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_631),
.B(n_501),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_631),
.B(n_501),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_713),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_628),
.A2(n_501),
.B1(n_632),
.B2(n_752),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_661),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_658),
.B(n_506),
.Y(n_910)
);

AND2x6_ASAP7_75t_L g911 ( 
.A(n_756),
.B(n_631),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_658),
.B(n_506),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_661),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_631),
.B(n_501),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_631),
.B(n_501),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_713),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_682),
.Y(n_917)
);

AO31x2_ASAP7_75t_L g918 ( 
.A1(n_891),
.A2(n_859),
.A3(n_801),
.B(n_897),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_823),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_895),
.A2(n_860),
.B(n_905),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_818),
.A2(n_792),
.B(n_892),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_904),
.B(n_905),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_908),
.B(n_854),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_854),
.B(n_853),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_770),
.Y(n_925)
);

AOI221xp5_ASAP7_75t_L g926 ( 
.A1(n_873),
.A2(n_858),
.B1(n_838),
.B2(n_816),
.C(n_880),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_906),
.B(n_914),
.Y(n_927)
);

AOI21xp33_ASAP7_75t_L g928 ( 
.A1(n_849),
.A2(n_863),
.B(n_894),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_805),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_778),
.B(n_799),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_877),
.B(n_870),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_906),
.B(n_914),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_812),
.B(n_901),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_901),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_769),
.A2(n_804),
.B(n_867),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_795),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_915),
.B(n_824),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_915),
.A2(n_862),
.B(n_865),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_805),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_867),
.A2(n_768),
.B(n_794),
.Y(n_940)
);

NOR2x1_ASAP7_75t_SL g941 ( 
.A(n_901),
.B(n_790),
.Y(n_941)
);

AOI21xp33_ASAP7_75t_L g942 ( 
.A1(n_848),
.A2(n_850),
.B(n_845),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_777),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_829),
.B(n_806),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_871),
.B(n_767),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_812),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_857),
.B(n_896),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_825),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_845),
.A2(n_848),
.B(n_850),
.C(n_874),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_898),
.B(n_775),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_857),
.B(n_896),
.Y(n_951)
);

AOI211x1_ASAP7_75t_L g952 ( 
.A1(n_880),
.A2(n_882),
.B(n_866),
.C(n_864),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_900),
.A2(n_912),
.B(n_910),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_896),
.B(n_911),
.Y(n_954)
);

OAI21x1_ASAP7_75t_SL g955 ( 
.A1(n_883),
.A2(n_847),
.B(n_821),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_852),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_784),
.Y(n_957)
);

AO31x2_ASAP7_75t_L g958 ( 
.A1(n_800),
.A2(n_776),
.A3(n_771),
.B(n_809),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_864),
.A2(n_782),
.B1(n_881),
.B2(n_840),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_896),
.B(n_911),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_899),
.A2(n_843),
.B(n_876),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_907),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_780),
.A2(n_843),
.B(n_878),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_916),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_787),
.A2(n_780),
.B(n_872),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_889),
.A2(n_896),
.B(n_911),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_811),
.B(n_834),
.Y(n_967)
);

AND2x2_ASAP7_75t_SL g968 ( 
.A(n_884),
.B(n_802),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_797),
.A2(n_813),
.B(n_827),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_830),
.A2(n_868),
.B1(n_813),
.B2(n_803),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_772),
.B(n_775),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_911),
.A2(n_827),
.B(n_793),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_911),
.B(n_788),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_SL g974 ( 
.A1(n_786),
.A2(n_835),
.B(n_885),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_869),
.A2(n_826),
.B(n_879),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_903),
.A2(n_913),
.B(n_909),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_814),
.B(n_820),
.Y(n_977)
);

INVx6_ASAP7_75t_SL g978 ( 
.A(n_825),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_826),
.A2(n_846),
.B(n_870),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_785),
.A2(n_798),
.B(n_856),
.C(n_781),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_796),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_890),
.B(n_893),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_796),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_789),
.B(n_832),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_890),
.A2(n_791),
.B1(n_833),
.B2(n_917),
.Y(n_985)
);

NAND2x1_ASAP7_75t_L g986 ( 
.A(n_819),
.B(n_917),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_817),
.A2(n_839),
.B(n_844),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_828),
.B(n_851),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_819),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_822),
.A2(n_887),
.B(n_886),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_855),
.B(n_837),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_855),
.B(n_831),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_836),
.A2(n_773),
.B(n_887),
.C(n_886),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_888),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_888),
.B(n_779),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_810),
.A2(n_842),
.B(n_875),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_810),
.A2(n_897),
.B(n_895),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_810),
.A2(n_807),
.B(n_861),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_842),
.B(n_506),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_842),
.B(n_908),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_908),
.B(n_854),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_815),
.A2(n_539),
.B(n_520),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_818),
.A2(n_792),
.B(n_892),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_818),
.A2(n_792),
.B(n_892),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_894),
.B(n_441),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_894),
.B(n_506),
.Y(n_1006)
);

CKINVDCx16_ASAP7_75t_R g1007 ( 
.A(n_779),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_815),
.A2(n_539),
.B(n_520),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_859),
.A2(n_849),
.B(n_860),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_894),
.B(n_441),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_774),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_441),
.Y(n_1012)
);

OA21x2_ASAP7_75t_L g1013 ( 
.A1(n_769),
.A2(n_801),
.B(n_800),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_815),
.A2(n_539),
.B(n_520),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_907),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_SL g1016 ( 
.A(n_901),
.B(n_761),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_799),
.B(n_700),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_774),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_L g1019 ( 
.A1(n_859),
.A2(n_849),
.B(n_897),
.C(n_895),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_812),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_770),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_895),
.A2(n_897),
.B(n_859),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_908),
.B(n_854),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_895),
.A2(n_897),
.B(n_859),
.Y(n_1024)
);

BUFx10_ASAP7_75t_L g1025 ( 
.A(n_884),
.Y(n_1025)
);

AOI221x1_ASAP7_75t_L g1026 ( 
.A1(n_859),
.A2(n_895),
.B1(n_897),
.B2(n_838),
.C(n_849),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_818),
.A2(n_792),
.B(n_892),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_908),
.B(n_854),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_818),
.A2(n_792),
.B(n_892),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_895),
.A2(n_897),
.B(n_859),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_770),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_901),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_815),
.A2(n_539),
.B(n_520),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_908),
.B(n_854),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_807),
.A2(n_861),
.B(n_808),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_894),
.B(n_506),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_860),
.A2(n_897),
.B(n_895),
.C(n_859),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_907),
.B(n_506),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_908),
.B(n_854),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_908),
.B(n_854),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_SL g1041 ( 
.A1(n_841),
.A2(n_902),
.B(n_783),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_1009),
.A2(n_928),
.B1(n_926),
.B2(n_945),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_936),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_919),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_1021),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_922),
.B(n_1005),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_924),
.B(n_927),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_925),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_928),
.A2(n_1019),
.B(n_938),
.C(n_1037),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_927),
.A2(n_932),
.B1(n_937),
.B2(n_924),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_932),
.B(n_937),
.Y(n_1051)
);

NOR2x1_ASAP7_75t_L g1052 ( 
.A(n_920),
.B(n_947),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_956),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_1017),
.B(n_994),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_SL g1055 ( 
.A(n_1006),
.B(n_1036),
.C(n_953),
.Y(n_1055)
);

BUFx4_ASAP7_75t_SL g1056 ( 
.A(n_981),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_982),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_926),
.A2(n_1023),
.B1(n_1040),
.B2(n_1039),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_962),
.B(n_946),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_934),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_944),
.B(n_923),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_944),
.B(n_923),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_949),
.A2(n_1028),
.B(n_1040),
.C(n_1023),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_SL g1065 ( 
.A(n_964),
.B(n_1015),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_992),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_L g1067 ( 
.A(n_946),
.B(n_1020),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_992),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_934),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1001),
.B(n_1028),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1002),
.A2(n_1008),
.B(n_1014),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_959),
.A2(n_1039),
.B1(n_1034),
.B2(n_1001),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_977),
.B(n_967),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_943),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_1020),
.B(n_948),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_934),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_989),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_1007),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1034),
.B(n_1031),
.Y(n_1079)
);

AND2x6_ASAP7_75t_L g1080 ( 
.A(n_948),
.B(n_929),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1038),
.B(n_950),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_1022),
.A2(n_1030),
.B(n_1024),
.C(n_942),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_950),
.B(n_994),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_SL g1084 ( 
.A1(n_942),
.A2(n_997),
.B(n_966),
.C(n_972),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_930),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_968),
.B(n_971),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_957),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_959),
.A2(n_980),
.B(n_985),
.C(n_965),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_939),
.B(n_952),
.Y(n_1089)
);

OR2x2_ASAP7_75t_SL g1090 ( 
.A(n_994),
.B(n_999),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1025),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1011),
.B(n_1018),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1017),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_970),
.A2(n_976),
.B1(n_1000),
.B2(n_951),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_988),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_940),
.B(n_1026),
.Y(n_1096)
);

NAND2xp33_ASAP7_75t_L g1097 ( 
.A(n_931),
.B(n_933),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_1000),
.A2(n_996),
.B(n_947),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_988),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_991),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_991),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_984),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_1017),
.B(n_995),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_995),
.B(n_1025),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1032),
.B(n_987),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_951),
.B(n_918),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_983),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_969),
.B(n_918),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_918),
.B(n_973),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_973),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_986),
.Y(n_1111)
);

NAND2x1_ASAP7_75t_L g1112 ( 
.A(n_1032),
.B(n_989),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_933),
.A2(n_993),
.B1(n_974),
.B2(n_954),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_L g1114 ( 
.A(n_931),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_941),
.B(n_1016),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_954),
.A2(n_960),
.B(n_990),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_998),
.A2(n_935),
.B(n_1035),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_978),
.B(n_960),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_990),
.B(n_958),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_963),
.B(n_1013),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_935),
.A2(n_1033),
.B1(n_1013),
.B2(n_978),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_931),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_958),
.B(n_963),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_975),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_931),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_921),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_958),
.B(n_979),
.Y(n_1127)
);

INVx6_ASAP7_75t_L g1128 ( 
.A(n_931),
.Y(n_1128)
);

OAI321xp33_ASAP7_75t_L g1129 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_1029),
.B1(n_1027),
.B2(n_961),
.C(n_1041),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_955),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_925),
.Y(n_1131)
);

BUFx4_ASAP7_75t_SL g1132 ( 
.A(n_981),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_1017),
.B(n_799),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_925),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_964),
.Y(n_1136)
);

BUFx2_ASAP7_75t_SL g1137 ( 
.A(n_1038),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_924),
.B(n_927),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_927),
.A2(n_860),
.B1(n_908),
.B2(n_859),
.Y(n_1140)
);

BUFx2_ASAP7_75t_SL g1141 ( 
.A(n_1038),
.Y(n_1141)
);

NAND2x1_ASAP7_75t_L g1142 ( 
.A(n_1032),
.B(n_901),
.Y(n_1142)
);

NAND2x1p5_ASAP7_75t_L g1143 ( 
.A(n_962),
.B(n_925),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_992),
.B(n_950),
.Y(n_1144)
);

BUFx12f_ASAP7_75t_L g1145 ( 
.A(n_964),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_934),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_998),
.A2(n_966),
.B(n_1022),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_934),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_928),
.A2(n_860),
.B(n_849),
.C(n_859),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1009),
.A2(n_859),
.B1(n_860),
.B2(n_858),
.Y(n_1151)
);

AOI222xp33_ASAP7_75t_SL g1152 ( 
.A1(n_996),
.A2(n_667),
.B1(n_432),
.B2(n_459),
.C1(n_441),
.C2(n_337),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1037),
.A2(n_1026),
.B(n_949),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1021),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_L g1155 ( 
.A(n_927),
.B(n_860),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_992),
.B(n_950),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_934),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_992),
.B(n_950),
.Y(n_1158)
);

CKINVDCx11_ASAP7_75t_R g1159 ( 
.A(n_981),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_964),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1017),
.B(n_799),
.Y(n_1162)
);

OR2x6_ASAP7_75t_SL g1163 ( 
.A(n_964),
.B(n_713),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1009),
.A2(n_853),
.B1(n_858),
.B2(n_859),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_992),
.B(n_950),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_928),
.A2(n_859),
.B(n_632),
.C(n_894),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_927),
.A2(n_860),
.B1(n_908),
.B2(n_859),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_992),
.B(n_950),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_928),
.A2(n_859),
.B(n_632),
.C(n_894),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1021),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_919),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_922),
.B(n_506),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_946),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_946),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_924),
.B(n_927),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1099),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1126),
.Y(n_1177)
);

BUFx2_ASAP7_75t_SL g1178 ( 
.A(n_1067),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1109),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1154),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1047),
.B(n_1175),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1119),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1133),
.B(n_1139),
.Y(n_1183)
);

OAI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1151),
.A2(n_1057),
.B1(n_1086),
.B2(n_1046),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1150),
.A2(n_1051),
.B1(n_1055),
.B2(n_1042),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1044),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1128),
.Y(n_1187)
);

NAND2x1p5_ASAP7_75t_L g1188 ( 
.A(n_1052),
.B(n_1130),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1138),
.B(n_1164),
.Y(n_1189)
);

INVx6_ASAP7_75t_L g1190 ( 
.A(n_1114),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1140),
.A2(n_1167),
.B1(n_1155),
.B2(n_1151),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1106),
.B(n_1070),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1043),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1148),
.A2(n_1161),
.B1(n_1052),
.B2(n_1059),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1043),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1056),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1053),
.Y(n_1197)
);

INVx8_ASAP7_75t_L g1198 ( 
.A(n_1080),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1050),
.B(n_1062),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1143),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1172),
.A2(n_1058),
.B1(n_1072),
.B2(n_1079),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1159),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1063),
.B(n_1072),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1127),
.B(n_1105),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1152),
.A2(n_1141),
.B1(n_1137),
.B2(n_1085),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1105),
.B(n_1122),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1045),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1110),
.B(n_1095),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1116),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1116),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1152),
.A2(n_1113),
.B1(n_1073),
.B2(n_1134),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1094),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1082),
.A2(n_1166),
.B1(n_1169),
.B2(n_1090),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1061),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1102),
.B(n_1089),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1171),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1098),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1098),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1049),
.A2(n_1088),
.B1(n_1170),
.B2(n_1153),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1048),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1147),
.B(n_1123),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1080),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1074),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1131),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1087),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1144),
.A2(n_1168),
.B1(n_1165),
.B2(n_1158),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1125),
.A2(n_1101),
.B1(n_1081),
.B2(n_1054),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1101),
.A2(n_1054),
.B1(n_1092),
.B2(n_1118),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1144),
.A2(n_1156),
.B1(n_1158),
.B2(n_1168),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1054),
.A2(n_1092),
.B1(n_1091),
.B2(n_1135),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1080),
.Y(n_1231)
);

NAND2x1p5_ASAP7_75t_L g1232 ( 
.A(n_1147),
.B(n_1124),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_SL g1233 ( 
.A(n_1145),
.Y(n_1233)
);

BUFx10_ASAP7_75t_L g1234 ( 
.A(n_1136),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1128),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1104),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1071),
.A2(n_1096),
.B(n_1108),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1064),
.B(n_1156),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1100),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1117),
.B(n_1115),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1117),
.B(n_1115),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1111),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1066),
.A2(n_1093),
.B1(n_1103),
.B2(n_1162),
.Y(n_1243)
);

INVx6_ASAP7_75t_L g1244 ( 
.A(n_1165),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1068),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1134),
.A2(n_1162),
.B1(n_1103),
.B2(n_1163),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1120),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1173),
.B(n_1174),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1174),
.B(n_1067),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1080),
.A2(n_1083),
.B1(n_1103),
.B2(n_1134),
.Y(n_1250)
);

AND2x2_ASAP7_75t_SL g1251 ( 
.A(n_1097),
.B(n_1084),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1083),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1121),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1060),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1075),
.B(n_1077),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1160),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1132),
.Y(n_1257)
);

INVx6_ASAP7_75t_L g1258 ( 
.A(n_1146),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1112),
.A2(n_1142),
.B(n_1129),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1162),
.A2(n_1075),
.B1(n_1065),
.B2(n_1107),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1069),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1069),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1078),
.A2(n_1146),
.B1(n_1076),
.B2(n_1149),
.Y(n_1263)
);

BUFx4f_ASAP7_75t_L g1264 ( 
.A(n_1076),
.Y(n_1264)
);

CKINVDCx8_ASAP7_75t_R g1265 ( 
.A(n_1076),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1149),
.B(n_1157),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1149),
.B(n_1129),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1114),
.Y(n_1268)
);

AO21x1_ASAP7_75t_L g1269 ( 
.A1(n_1166),
.A2(n_1169),
.B(n_928),
.Y(n_1269)
);

BUFx2_ASAP7_75t_R g1270 ( 
.A(n_1078),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_L g1271 ( 
.A(n_1114),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1043),
.Y(n_1272)
);

BUFx4f_ASAP7_75t_SL g1273 ( 
.A(n_1145),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1086),
.A2(n_858),
.B1(n_853),
.B2(n_459),
.Y(n_1274)
);

BUFx2_ASAP7_75t_R g1275 ( 
.A(n_1078),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1150),
.A2(n_860),
.B(n_894),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1154),
.Y(n_1277)
);

BUFx2_ASAP7_75t_SL g1278 ( 
.A(n_1067),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1175),
.B(n_1047),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1056),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1044),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1043),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1043),
.Y(n_1283)
);

AO21x1_ASAP7_75t_L g1284 ( 
.A1(n_1166),
.A2(n_1169),
.B(n_928),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1143),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1044),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1130),
.Y(n_1287)
);

INVx4_ASAP7_75t_SL g1288 ( 
.A(n_1190),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1247),
.B(n_1179),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1247),
.B(n_1179),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1193),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1287),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1240),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1182),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1276),
.A2(n_1185),
.B1(n_1211),
.B2(n_1191),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1177),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1287),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1199),
.B(n_1203),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1198),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1195),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1203),
.B(n_1192),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1199),
.B(n_1181),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1196),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1181),
.B(n_1279),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1232),
.Y(n_1305)
);

AO21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1212),
.A2(n_1253),
.B(n_1218),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1232),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1192),
.B(n_1217),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1272),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1237),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1217),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1256),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1218),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1269),
.A2(n_1284),
.B(n_1253),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1213),
.A2(n_1212),
.A3(n_1209),
.B(n_1210),
.Y(n_1315)
);

BUFx2_ASAP7_75t_SL g1316 ( 
.A(n_1265),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1204),
.B(n_1279),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1241),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1241),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1189),
.B(n_1215),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1188),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1188),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1221),
.B(n_1184),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1189),
.B(n_1215),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1283),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1208),
.B(n_1219),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1243),
.A2(n_1259),
.B(n_1238),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1198),
.B(n_1206),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1259),
.A2(n_1242),
.B(n_1267),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1249),
.B(n_1222),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1208),
.B(n_1201),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1221),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1206),
.A2(n_1216),
.B(n_1223),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1197),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1249),
.B(n_1231),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1251),
.B(n_1176),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1267),
.A2(n_1286),
.B(n_1281),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1194),
.A2(n_1267),
.B(n_1186),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1251),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1274),
.A2(n_1205),
.B1(n_1246),
.B2(n_1183),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1231),
.B(n_1178),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1239),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1225),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1236),
.B(n_1282),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1190),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1220),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_R g1347 ( 
.A(n_1339),
.B(n_1190),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1332),
.B(n_1248),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1306),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1337),
.B(n_1228),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1337),
.B(n_1230),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1332),
.B(n_1248),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1298),
.B(n_1308),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1337),
.B(n_1227),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1306),
.Y(n_1355)
);

NOR4xp25_ASAP7_75t_SL g1356 ( 
.A(n_1339),
.B(n_1280),
.C(n_1196),
.D(n_1252),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1295),
.A2(n_1244),
.B1(n_1207),
.B2(n_1271),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1337),
.B(n_1207),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1292),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1318),
.B(n_1255),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1318),
.B(n_1255),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1298),
.B(n_1260),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1318),
.B(n_1266),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1308),
.B(n_1301),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1294),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1319),
.B(n_1266),
.Y(n_1366)
);

NOR2x1_ASAP7_75t_R g1367 ( 
.A(n_1303),
.B(n_1280),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1310),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1292),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1293),
.B(n_1268),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1309),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1305),
.B(n_1250),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1329),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1301),
.B(n_1278),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1296),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1329),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1312),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1329),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1315),
.B(n_1278),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1293),
.B(n_1268),
.Y(n_1380)
);

INVx5_ASAP7_75t_L g1381 ( 
.A(n_1328),
.Y(n_1381)
);

INVxp67_ASAP7_75t_R g1382 ( 
.A(n_1333),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1315),
.B(n_1263),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1375),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1371),
.B(n_1320),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1371),
.B(n_1320),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1360),
.B(n_1317),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1340),
.C(n_1344),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1324),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1360),
.B(n_1317),
.Y(n_1390)
);

AND2x2_ASAP7_75t_SL g1391 ( 
.A(n_1349),
.B(n_1338),
.Y(n_1391)
);

AND2x2_ASAP7_75t_SL g1392 ( 
.A(n_1349),
.B(n_1338),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1368),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1360),
.B(n_1329),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1362),
.A2(n_1323),
.B1(n_1326),
.B2(n_1316),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1357),
.A2(n_1331),
.B1(n_1326),
.B2(n_1302),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1353),
.B(n_1324),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1362),
.A2(n_1331),
.B1(n_1302),
.B2(n_1316),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1374),
.B(n_1309),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1374),
.B(n_1291),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1364),
.B(n_1300),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1364),
.B(n_1325),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1372),
.A2(n_1323),
.B1(n_1335),
.B2(n_1330),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1307),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1375),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1361),
.B(n_1334),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1356),
.A2(n_1271),
.B1(n_1341),
.B2(n_1304),
.Y(n_1407)
);

NAND4xp25_ASAP7_75t_L g1408 ( 
.A(n_1383),
.B(n_1336),
.C(n_1342),
.D(n_1304),
.Y(n_1408)
);

NAND4xp25_ASAP7_75t_L g1409 ( 
.A(n_1383),
.B(n_1342),
.C(n_1313),
.D(n_1311),
.Y(n_1409)
);

OAI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1351),
.A2(n_1229),
.B1(n_1226),
.B2(n_1271),
.C(n_1257),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_L g1411 ( 
.A(n_1377),
.B(n_1299),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1348),
.B(n_1346),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1348),
.B(n_1315),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1359),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1363),
.B(n_1307),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1351),
.A2(n_1190),
.B1(n_1345),
.B2(n_1180),
.C(n_1277),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1348),
.B(n_1315),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1352),
.B(n_1315),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1354),
.B(n_1314),
.C(n_1343),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1352),
.B(n_1315),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1352),
.B(n_1343),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1363),
.B(n_1297),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1363),
.B(n_1297),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1354),
.B(n_1379),
.C(n_1314),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1379),
.B(n_1345),
.C(n_1327),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1354),
.B(n_1314),
.C(n_1313),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1350),
.A2(n_1268),
.B(n_1299),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_SL g1428 ( 
.A(n_1369),
.B(n_1322),
.C(n_1321),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1366),
.B(n_1289),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1367),
.B(n_1303),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1366),
.B(n_1289),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1366),
.B(n_1290),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1387),
.B(n_1381),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1430),
.B(n_1367),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1387),
.B(n_1381),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1384),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1384),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1405),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1405),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1390),
.B(n_1381),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1414),
.B(n_1359),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1393),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1393),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1421),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1413),
.B(n_1369),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1390),
.B(n_1381),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1409),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1417),
.B(n_1358),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1394),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1418),
.B(n_1358),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1420),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1391),
.B(n_1392),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1391),
.B(n_1373),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1400),
.B(n_1303),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1391),
.B(n_1392),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1358),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1419),
.B(n_1381),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1389),
.B(n_1314),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1397),
.B(n_1314),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1424),
.B(n_1351),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1424),
.B(n_1365),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1404),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1385),
.B(n_1365),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1398),
.B(n_1345),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1392),
.B(n_1415),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1423),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1386),
.B(n_1401),
.Y(n_1468)
);

AND2x4_ASAP7_75t_SL g1469 ( 
.A(n_1428),
.B(n_1349),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1406),
.B(n_1350),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1429),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1431),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1412),
.B(n_1381),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1449),
.B(n_1419),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1453),
.B(n_1381),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1458),
.B(n_1381),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1436),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1436),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1437),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1442),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1448),
.B(n_1399),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1453),
.B(n_1427),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1434),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1382),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1455),
.B(n_1202),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1437),
.Y(n_1486)
);

OAI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1461),
.A2(n_1408),
.B(n_1395),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1464),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1456),
.B(n_1382),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1442),
.Y(n_1490)
);

INVxp33_ASAP7_75t_SL g1491 ( 
.A(n_1465),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1448),
.B(n_1202),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1438),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1438),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1439),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1445),
.B(n_1402),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1458),
.B(n_1425),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1464),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1439),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1441),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1441),
.Y(n_1501)
);

NAND2x1_ASAP7_75t_L g1502 ( 
.A(n_1454),
.B(n_1349),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1466),
.B(n_1382),
.Y(n_1503)
);

NOR3xp33_ASAP7_75t_L g1504 ( 
.A(n_1461),
.B(n_1388),
.C(n_1416),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1462),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1468),
.B(n_1234),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1449),
.B(n_1426),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1445),
.B(n_1432),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1462),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1433),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1466),
.B(n_1349),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1442),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1467),
.B(n_1396),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1483),
.B(n_1233),
.Y(n_1514)
);

OAI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1504),
.A2(n_1454),
.B(n_1388),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1477),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1483),
.B(n_1273),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1491),
.Y(n_1518)
);

AOI322xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1482),
.A2(n_1454),
.A3(n_1463),
.B1(n_1440),
.B2(n_1447),
.C1(n_1435),
.C2(n_1433),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1513),
.B(n_1487),
.Y(n_1520)
);

INVxp33_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1482),
.B(n_1435),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_SL g1523 ( 
.A(n_1491),
.B(n_1270),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1507),
.B(n_1451),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1495),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1477),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1475),
.B(n_1469),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1511),
.B(n_1440),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1511),
.B(n_1447),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1478),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1507),
.B(n_1451),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1495),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1488),
.B(n_1452),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1478),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1498),
.B(n_1471),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1500),
.B(n_1471),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1501),
.B(n_1472),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1472),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1480),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1475),
.A2(n_1411),
.B1(n_1407),
.B2(n_1469),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1480),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1496),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1510),
.B(n_1444),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1476),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1509),
.B(n_1468),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1485),
.B(n_1234),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1479),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1509),
.B(n_1470),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1508),
.B(n_1470),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1474),
.B(n_1459),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1490),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1502),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1515),
.B(n_1510),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1518),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1523),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1529),
.B(n_1497),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1528),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1527),
.Y(n_1562)
);

NOR2x1_ASAP7_75t_L g1563 ( 
.A(n_1514),
.B(n_1502),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1522),
.B(n_1484),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1522),
.B(n_1484),
.Y(n_1565)
);

NOR2x1_ASAP7_75t_L g1566 ( 
.A(n_1517),
.B(n_1497),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1520),
.A2(n_1497),
.B1(n_1489),
.B2(n_1410),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1521),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1530),
.B(n_1489),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1544),
.B(n_1474),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1521),
.A2(n_1529),
.B1(n_1540),
.B2(n_1542),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1528),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1551),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1534),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1516),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1532),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1525),
.A2(n_1503),
.B1(n_1476),
.B2(n_1469),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1536),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.B(n_1459),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1525),
.Y(n_1582)
);

AOI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1547),
.A2(n_1549),
.B1(n_1524),
.B2(n_1552),
.C(n_1537),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1527),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1535),
.A2(n_1426),
.B1(n_1460),
.B2(n_1499),
.C(n_1493),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1530),
.A2(n_1411),
.B1(n_1503),
.B2(n_1473),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1548),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1548),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1550),
.B(n_1256),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1538),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1568),
.A2(n_1519),
.B1(n_1554),
.B2(n_1533),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1531),
.Y(n_1594)
);

AOI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1566),
.A2(n_1556),
.B(n_1533),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1531),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1557),
.A2(n_1519),
.B1(n_1554),
.B2(n_1556),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1572),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1573),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1574),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1580),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1563),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1585),
.A2(n_1546),
.B1(n_1539),
.B2(n_1553),
.C(n_1555),
.Y(n_1605)
);

XOR2x2_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1275),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1571),
.A2(n_1534),
.B(n_1350),
.C(n_1200),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1583),
.B(n_1543),
.C(n_1541),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1570),
.A2(n_1579),
.B(n_1582),
.Y(n_1609)
);

OAI222xp33_ASAP7_75t_L g1610 ( 
.A1(n_1587),
.A2(n_1545),
.B1(n_1555),
.B2(n_1543),
.C1(n_1473),
.C2(n_1446),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1545),
.C(n_1356),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1589),
.B(n_1479),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1560),
.B(n_1564),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1560),
.A2(n_1380),
.B1(n_1370),
.B2(n_1355),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1592),
.B(n_1486),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1577),
.Y(n_1617)
);

OAI211xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1578),
.A2(n_1224),
.B(n_1446),
.C(n_1180),
.Y(n_1618)
);

NOR2x1_ASAP7_75t_L g1619 ( 
.A(n_1615),
.B(n_1560),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1594),
.B(n_1591),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1602),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1603),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1597),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1596),
.B(n_1564),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1615),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1599),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1613),
.B(n_1565),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1604),
.B(n_1565),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1609),
.B(n_1569),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1617),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1616),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1593),
.B(n_1575),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1618),
.B(n_1591),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1593),
.B(n_1576),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1612),
.Y(n_1638)
);

AOI21xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1637),
.A2(n_1598),
.B(n_1611),
.Y(n_1639)
);

OAI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1635),
.A2(n_1598),
.B1(n_1607),
.B2(n_1605),
.C(n_1608),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1619),
.B(n_1607),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1637),
.A2(n_1576),
.B1(n_1562),
.B2(n_1584),
.Y(n_1642)
);

NAND4xp75_ASAP7_75t_L g1643 ( 
.A(n_1635),
.B(n_1590),
.C(n_1614),
.D(n_1586),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1630),
.A2(n_1610),
.B1(n_1576),
.B2(n_1588),
.C(n_1581),
.Y(n_1644)
);

AOI32xp33_ASAP7_75t_L g1645 ( 
.A1(n_1630),
.A2(n_1588),
.A3(n_1581),
.B1(n_1606),
.B2(n_1512),
.Y(n_1645)
);

OAI211xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1624),
.A2(n_1606),
.B(n_1277),
.C(n_1494),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1620),
.A2(n_1486),
.B1(n_1494),
.B2(n_1512),
.C(n_1376),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1631),
.A2(n_1347),
.B1(n_1376),
.B2(n_1373),
.C1(n_1378),
.C2(n_1450),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1638),
.B(n_1627),
.C(n_1629),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1625),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1650),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1641),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1640),
.A2(n_1631),
.B(n_1636),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1639),
.B(n_1628),
.C(n_1638),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1643),
.Y(n_1655)
);

NAND2x1_ASAP7_75t_SL g1656 ( 
.A(n_1645),
.B(n_1628),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1642),
.B(n_1632),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1649),
.B(n_1633),
.C(n_1621),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1644),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1646),
.B(n_1633),
.C(n_1626),
.Y(n_1660)
);

NOR4xp25_ASAP7_75t_L g1661 ( 
.A(n_1647),
.B(n_1622),
.C(n_1623),
.D(n_1626),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1648),
.B(n_1634),
.Y(n_1662)
);

NAND4xp25_ASAP7_75t_SL g1663 ( 
.A(n_1659),
.B(n_1623),
.C(n_1622),
.D(n_1632),
.Y(n_1663)
);

NAND2x1_ASAP7_75t_L g1664 ( 
.A(n_1651),
.B(n_1268),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1656),
.A2(n_1265),
.B(n_1268),
.C(n_1285),
.Y(n_1665)
);

NOR3x1_ASAP7_75t_SL g1666 ( 
.A(n_1655),
.B(n_1234),
.C(n_1463),
.Y(n_1666)
);

NOR3x1_ASAP7_75t_L g1667 ( 
.A(n_1654),
.B(n_1245),
.C(n_1457),
.Y(n_1667)
);

NAND4xp25_ASAP7_75t_SL g1668 ( 
.A(n_1653),
.B(n_1450),
.C(n_1444),
.D(n_1403),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1657),
.A2(n_1347),
.B(n_1285),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1666),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1664),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1667),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1668),
.Y(n_1675)
);

NAND4xp75_ASAP7_75t_L g1676 ( 
.A(n_1670),
.B(n_1653),
.C(n_1662),
.D(n_1669),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1675),
.Y(n_1677)
);

NAND4xp75_ASAP7_75t_L g1678 ( 
.A(n_1671),
.B(n_1652),
.C(n_1658),
.D(n_1660),
.Y(n_1678)
);

OAI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1674),
.A2(n_1200),
.B(n_1245),
.C(n_1214),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1674),
.B(n_1457),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1678),
.B(n_1672),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1680),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_SL g1683 ( 
.A(n_1679),
.B(n_1673),
.C(n_1214),
.Y(n_1683)
);

INVxp33_ASAP7_75t_SL g1684 ( 
.A(n_1682),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1681),
.B1(n_1677),
.B2(n_1683),
.C(n_1676),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1264),
.B(n_1254),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1685),
.A2(n_1235),
.B(n_1187),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1444),
.B1(n_1450),
.B2(n_1288),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1686),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1688),
.A2(n_1262),
.B1(n_1258),
.B2(n_1264),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1690),
.B(n_1254),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1691),
.B1(n_1262),
.B2(n_1264),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1214),
.B1(n_1261),
.B2(n_1443),
.C(n_1370),
.Y(n_1694)
);

AOI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1261),
.B(n_1299),
.C(n_1235),
.Y(n_1695)
);


endmodule