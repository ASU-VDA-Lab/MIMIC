module fake_ariane_417_n_1686 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1686);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1686;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g153 ( 
.A(n_48),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_21),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_21),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_60),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_20),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_84),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_52),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_82),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_77),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_63),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_56),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_3),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_137),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_58),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_81),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_32),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_53),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_23),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_23),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_116),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_104),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_95),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_37),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_83),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_69),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_10),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_42),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_49),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_44),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_103),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_121),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_98),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_86),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_25),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_50),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_85),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_79),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_78),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_129),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_134),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_87),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_48),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_62),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_9),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_1),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_52),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_132),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_41),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_17),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_133),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_102),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_59),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_109),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_34),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_67),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_7),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_16),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_71),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_33),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_6),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_90),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_100),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_19),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_146),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_41),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_143),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_142),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_35),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_4),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_17),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_118),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_110),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_4),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_27),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_22),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_147),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_47),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_45),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_135),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_105),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_29),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_36),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_20),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_89),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_70),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_10),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_112),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_12),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_53),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_50),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_145),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_7),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_22),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_68),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_29),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_55),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_57),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_66),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_91),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_33),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_75),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_15),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_122),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_5),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_5),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_61),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_73),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_31),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_34),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_8),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_181),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_185),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_246),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_263),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_178),
.B(n_1),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_200),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_233),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_212),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_185),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_204),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_265),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_185),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_216),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_224),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_226),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_307),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_227),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_201),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_248),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_228),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_185),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_203),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_240),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_253),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_308),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_158),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_203),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_R g342 ( 
.A(n_197),
.B(n_101),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_203),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_203),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_158),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_165),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_203),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_277),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_R g350 ( 
.A(n_198),
.B(n_126),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_154),
.B(n_2),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_165),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_228),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_160),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_169),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_242),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_247),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_286),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_169),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_174),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_264),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_286),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_286),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_201),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_175),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_264),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_175),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_247),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_285),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_179),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_189),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_247),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_189),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_179),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_187),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_258),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_258),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_187),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_258),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_231),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_231),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_311),
.B(n_161),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_287),
.B1(n_274),
.B2(n_281),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_318),
.B(n_258),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_321),
.B(n_162),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_164),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_309),
.B(n_333),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_255),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_333),
.B(n_353),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_353),
.B(n_258),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_168),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_347),
.B(n_348),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_173),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_176),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_205),
.B(n_199),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_357),
.A2(n_257),
.B1(n_300),
.B2(n_272),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_322),
.A2(n_257),
.B1(n_266),
.B2(n_272),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_351),
.B(n_317),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_374),
.B(n_255),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_285),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_206),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_369),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_319),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_314),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_192),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_331),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_210),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_366),
.B(n_220),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_342),
.B(n_222),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_350),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_345),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_326),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_328),
.C(n_327),
.Y(n_463)
);

NAND2x1p5_ASAP7_75t_L g464 ( 
.A(n_423),
.B(n_213),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_444),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_402),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_385),
.B1(n_384),
.B2(n_382),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_423),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_330),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_332),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_418),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

AND2x2_ASAP7_75t_SL g474 ( 
.A(n_451),
.B(n_209),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_418),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_403),
.B(n_413),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_451),
.A2(n_431),
.B1(n_402),
.B2(n_394),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_428),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_418),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_426),
.B(n_338),
.C(n_337),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_423),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_445),
.B(n_315),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_423),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

NAND3xp33_ASAP7_75t_L g492 ( 
.A(n_426),
.B(n_456),
.C(n_408),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_413),
.B(n_408),
.Y(n_493)
);

CKINVDCx11_ASAP7_75t_R g494 ( 
.A(n_457),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_392),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_392),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_423),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_432),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_402),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_431),
.B(n_346),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_413),
.B(n_352),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_399),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_394),
.B(n_355),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_442),
.B(n_360),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_423),
.B(n_361),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_404),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_404),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_423),
.B(n_367),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_370),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_442),
.B(n_379),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_451),
.B(n_377),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_451),
.B(n_375),
.Y(n_521)
);

OAI22xp33_ASAP7_75t_L g522 ( 
.A1(n_389),
.A2(n_320),
.B1(n_310),
.B2(n_324),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_423),
.B(n_313),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_439),
.B(n_167),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_409),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_456),
.B(n_320),
.C(n_279),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_439),
.B(n_207),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_452),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_447),
.B(n_155),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_452),
.B(n_188),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_452),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_443),
.B(n_312),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_448),
.A2(n_251),
.B1(n_230),
.B2(n_236),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_448),
.A2(n_202),
.B1(n_273),
.B2(n_275),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_415),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_447),
.B(n_155),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_458),
.A2(n_232),
.B(n_225),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_454),
.B(n_188),
.Y(n_548)
);

INVx8_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_454),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_437),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_415),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_410),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_410),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_407),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_447),
.B(n_458),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_454),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_439),
.B(n_448),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_447),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_407),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_445),
.B(n_188),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_407),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_407),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_448),
.B(n_160),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_457),
.A2(n_266),
.B1(n_279),
.B2(n_280),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_441),
.B(n_270),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_457),
.A2(n_293),
.B1(n_280),
.B2(n_281),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_445),
.B(n_289),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_411),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_448),
.B(n_160),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_411),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_425),
.Y(n_577)
);

INVx4_ASAP7_75t_SL g578 ( 
.A(n_393),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_453),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_411),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_446),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_448),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_421),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_446),
.B(n_450),
.C(n_449),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_393),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_441),
.B(n_453),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_428),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_411),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_449),
.B(n_450),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_411),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_424),
.B(n_255),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_389),
.A2(n_183),
.B1(n_190),
.B2(n_214),
.Y(n_594)
);

AO22x2_ASAP7_75t_L g595 ( 
.A1(n_455),
.A2(n_192),
.B1(n_235),
.B2(n_299),
.Y(n_595)
);

INVx6_ASAP7_75t_L g596 ( 
.A(n_411),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_424),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_427),
.B(n_209),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_455),
.B(n_340),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_438),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_387),
.B(n_159),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_387),
.B(n_159),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_427),
.B(n_252),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_429),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_395),
.B(n_349),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_587),
.B(n_356),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_471),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_549),
.B(n_163),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_579),
.B(n_359),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_600),
.B(n_363),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_520),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_475),
.Y(n_614)
);

BUFx6f_ASAP7_75t_SL g615 ( 
.A(n_474),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_492),
.A2(n_256),
.B(n_284),
.C(n_292),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_474),
.A2(n_579),
.B1(n_503),
.B2(n_549),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_534),
.B(n_365),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_549),
.B(n_163),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_549),
.A2(n_303),
.B1(n_299),
.B2(n_235),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_562),
.B(n_484),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_562),
.B(n_166),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_484),
.B(n_166),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_470),
.B(n_323),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_475),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_534),
.B(n_395),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_484),
.B(n_170),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_487),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_493),
.B(n_170),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_605),
.B(n_171),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_520),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_566),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_606),
.B(n_329),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_487),
.B(n_196),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_507),
.A2(n_561),
.B1(n_460),
.B2(n_478),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_539),
.B(n_397),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_561),
.A2(n_302),
.B1(n_195),
.B2(n_194),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_595),
.A2(n_425),
.B1(n_436),
.B2(n_435),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_482),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_605),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_561),
.A2(n_302),
.B1(n_195),
.B2(n_194),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_469),
.B(n_444),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_482),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_528),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_539),
.B(n_397),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_527),
.A2(n_425),
.B(n_414),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_605),
.B(n_171),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_564),
.B(n_196),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_528),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_550),
.B(n_414),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_538),
.B(n_238),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_564),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_486),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_550),
.B(n_417),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_486),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_538),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_560),
.B(n_417),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_490),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_548),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_551),
.B(n_444),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_477),
.B(n_172),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_490),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_560),
.B(n_422),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_593),
.B(n_289),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_462),
.B(n_444),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_548),
.B(n_466),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_571),
.B(n_422),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_460),
.B(n_172),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_488),
.B(n_291),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_581),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_533),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_488),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_559),
.A2(n_396),
.B(n_391),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_497),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_466),
.B(n_196),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_497),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_498),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_508),
.A2(n_276),
.B1(n_193),
.B2(n_191),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_533),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_518),
.B(n_429),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_552),
.B(n_430),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_535),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_502),
.B(n_177),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_535),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_552),
.B(n_430),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_502),
.B(n_177),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_498),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_467),
.B(n_291),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_526),
.B(n_433),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_499),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_532),
.B(n_433),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_581),
.B(n_243),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_595),
.A2(n_425),
.B1(n_436),
.B2(n_435),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_537),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_499),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_505),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_593),
.B(n_293),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_504),
.A2(n_300),
.B1(n_298),
.B2(n_306),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_519),
.B(n_244),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_505),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_602),
.A2(n_391),
.B(n_396),
.C(n_250),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_471),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_481),
.B(n_245),
.C(n_259),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_590),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_496),
.B(n_180),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_537),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_566),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_517),
.A2(n_182),
.B1(n_184),
.B2(n_186),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_547),
.B(n_182),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_496),
.B(n_184),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_540),
.B(n_269),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_543),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_521),
.B(n_416),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_585),
.B(n_213),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_SL g715 ( 
.A1(n_479),
.A2(n_260),
.B1(n_193),
.B2(n_191),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_543),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_509),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_573),
.A2(n_416),
.B(n_295),
.C(n_290),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_461),
.B(n_260),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_547),
.B(n_261),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_465),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_545),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_547),
.B(n_261),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_573),
.B(n_262),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_509),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_SL g726 ( 
.A(n_465),
.B(n_269),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_461),
.B(n_262),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_463),
.B(n_269),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_472),
.B(n_271),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_596),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_511),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_545),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_483),
.B(n_271),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_593),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_483),
.B(n_276),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_494),
.B(n_278),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_595),
.A2(n_249),
.B1(n_239),
.B2(n_297),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_572),
.B(n_278),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_472),
.B(n_288),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_468),
.B(n_485),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_511),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_513),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_491),
.B(n_288),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_536),
.B(n_294),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_566),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_491),
.B(n_294),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_541),
.B(n_239),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_553),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_553),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_495),
.B(n_305),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_495),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_501),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_546),
.B(n_305),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_594),
.A2(n_267),
.B1(n_252),
.B2(n_282),
.C(n_249),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_501),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_506),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_512),
.B(n_208),
.Y(n_757)
);

AOI22x1_ASAP7_75t_L g758 ( 
.A1(n_473),
.A2(n_396),
.B1(n_391),
.B2(n_388),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_512),
.B(n_211),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_473),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_476),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_603),
.B(n_217),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_476),
.B(n_218),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_513),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_480),
.B(n_282),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_593),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_480),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_514),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_522),
.B(n_219),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_588),
.B(n_438),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_632),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_672),
.B(n_479),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_648),
.B(n_569),
.Y(n_773)
);

AOI21x1_ASAP7_75t_L g774 ( 
.A1(n_765),
.A2(n_556),
.B(n_557),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_726),
.Y(n_775)
);

INVx5_ASAP7_75t_L g776 ( 
.A(n_740),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_608),
.B(n_529),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_613),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_660),
.B(n_542),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_615),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_613),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_667),
.B(n_582),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_760),
.A2(n_489),
.B(n_510),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_760),
.A2(n_767),
.B(n_761),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_642),
.B(n_524),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_628),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_761),
.A2(n_489),
.B(n_516),
.Y(n_787)
);

AOI33xp33_ASAP7_75t_L g788 ( 
.A1(n_704),
.A2(n_523),
.A3(n_525),
.B1(n_530),
.B2(n_544),
.B3(n_555),
.Y(n_788)
);

AO21x1_ASAP7_75t_L g789 ( 
.A1(n_709),
.A2(n_464),
.B(n_523),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_666),
.B(n_525),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_615),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_617),
.B(n_566),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_631),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_767),
.A2(n_489),
.B(n_500),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_751),
.A2(n_468),
.B(n_485),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_666),
.B(n_530),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_666),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_751),
.A2(n_500),
.B(n_592),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_752),
.A2(n_756),
.B(n_755),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_659),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_752),
.A2(n_557),
.B(n_584),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_668),
.A2(n_556),
.B(n_598),
.C(n_555),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_755),
.A2(n_544),
.B(n_568),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_631),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_659),
.B(n_568),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_756),
.A2(n_598),
.B(n_592),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_635),
.A2(n_567),
.B(n_575),
.C(n_531),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_632),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_640),
.B(n_566),
.Y(n_810)
);

AO21x1_ASAP7_75t_L g811 ( 
.A1(n_720),
.A2(n_464),
.B(n_567),
.Y(n_811)
);

AO22x1_ASAP7_75t_L g812 ( 
.A1(n_612),
.A2(n_593),
.B1(n_599),
.B2(n_604),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_615),
.A2(n_604),
.B1(n_599),
.B2(n_527),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_668),
.A2(n_601),
.B(n_597),
.C(n_583),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_770),
.B(n_593),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_765),
.A2(n_673),
.B(n_625),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_614),
.A2(n_575),
.B(n_601),
.C(n_531),
.Y(n_817)
);

AND2x4_ASAP7_75t_SL g818 ( 
.A(n_640),
.B(n_527),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_639),
.A2(n_531),
.B(n_601),
.C(n_583),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_768),
.A2(n_464),
.B1(n_597),
.B2(n_583),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_SL g821 ( 
.A(n_633),
.B(n_223),
.C(n_221),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_721),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_632),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_670),
.B(n_599),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_680),
.A2(n_636),
.B(n_626),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_644),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_643),
.Y(n_827)
);

AO22x1_ASAP7_75t_L g828 ( 
.A1(n_721),
.A2(n_769),
.B1(n_665),
.B2(n_624),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_656),
.B(n_599),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_652),
.B(n_651),
.Y(n_830)
);

AOI21x1_ASAP7_75t_L g831 ( 
.A1(n_653),
.A2(n_565),
.B(n_554),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_651),
.B(n_599),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_651),
.B(n_599),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_655),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_658),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_662),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_713),
.B(n_599),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_621),
.B(n_577),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_621),
.B(n_577),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_646),
.A2(n_563),
.B(n_554),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_711),
.B(n_604),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_632),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_675),
.B(n_604),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_645),
.B(n_604),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_650),
.A2(n_597),
.B(n_558),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_654),
.A2(n_558),
.B(n_591),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_734),
.B(n_570),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_657),
.A2(n_574),
.B(n_563),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_663),
.B(n_565),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_692),
.B(n_574),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_674),
.A2(n_596),
.B1(n_576),
.B2(n_580),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_611),
.B(n_576),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_692),
.B(n_580),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_630),
.A2(n_596),
.B1(n_589),
.B2(n_570),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_622),
.B(n_596),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_707),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_692),
.B(n_570),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_676),
.A2(n_589),
.B(n_570),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_724),
.B(n_570),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_734),
.B(n_589),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_677),
.A2(n_589),
.B(n_586),
.Y(n_861)
);

AO21x1_ASAP7_75t_L g862 ( 
.A1(n_723),
.A2(n_388),
.B(n_401),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_687),
.A2(n_695),
.B(n_690),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_696),
.A2(n_717),
.B(n_700),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_707),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_725),
.Y(n_866)
);

CKINVDCx10_ASAP7_75t_R g867 ( 
.A(n_715),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_731),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_622),
.B(n_589),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_741),
.A2(n_586),
.B(n_515),
.Y(n_870)
);

AOI21x1_ASAP7_75t_L g871 ( 
.A1(n_742),
.A2(n_388),
.B(n_401),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_707),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_766),
.B(n_586),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_618),
.B(n_2),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_707),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_764),
.A2(n_586),
.B1(n_515),
.B2(n_391),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_649),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_607),
.A2(n_515),
.B(n_396),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_766),
.B(n_515),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_634),
.B(n_438),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_669),
.B(n_438),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_736),
.B(n_438),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_714),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_758),
.A2(n_578),
.B(n_438),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_607),
.B(n_578),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_689),
.B(n_578),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_691),
.B(n_578),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_698),
.B(n_297),
.C(n_254),
.Y(n_888)
);

OR2x6_ASAP7_75t_SL g889 ( 
.A(n_699),
.B(n_241),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_681),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_623),
.B(n_3),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_745),
.Y(n_892)
);

O2A1O1Ixp5_ASAP7_75t_L g893 ( 
.A1(n_661),
.A2(n_6),
.B(n_8),
.C(n_11),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_609),
.A2(n_702),
.B(n_763),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_738),
.B(n_11),
.Y(n_895)
);

AOI33xp33_ASAP7_75t_L g896 ( 
.A1(n_678),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.B3(n_19),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_609),
.A2(n_237),
.B(n_234),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_616),
.B(n_229),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_616),
.B(n_630),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_609),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_685),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_SL g902 ( 
.A(n_728),
.B(n_215),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_647),
.B(n_13),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_647),
.B(n_14),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_708),
.B(n_683),
.Y(n_905)
);

O2A1O1Ixp5_ASAP7_75t_L g906 ( 
.A1(n_623),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_745),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_637),
.B(n_26),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_702),
.B(n_398),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_702),
.B(n_30),
.Y(n_910)
);

NAND2x1p5_ASAP7_75t_L g911 ( 
.A(n_745),
.B(n_215),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_714),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_718),
.A2(n_215),
.B(n_160),
.C(n_393),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_629),
.A2(n_31),
.B(n_32),
.C(n_36),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_629),
.B(n_37),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_744),
.A2(n_215),
.B(n_160),
.C(n_393),
.Y(n_916)
);

OAI321xp33_ASAP7_75t_L g917 ( 
.A1(n_737),
.A2(n_215),
.A3(n_398),
.B1(n_393),
.B2(n_42),
.C(n_43),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_627),
.A2(n_683),
.B(n_686),
.C(n_610),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_753),
.B(n_38),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_757),
.A2(n_398),
.B(n_74),
.Y(n_920)
);

AO21x2_ASAP7_75t_L g921 ( 
.A1(n_719),
.A2(n_398),
.B(n_76),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_759),
.A2(n_398),
.B(n_64),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_671),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_610),
.A2(n_398),
.B1(n_39),
.B2(n_40),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_714),
.B(n_38),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_641),
.B(n_39),
.Y(n_926)
);

AND2x6_ASAP7_75t_L g927 ( 
.A(n_747),
.B(n_80),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_L g928 ( 
.A1(n_627),
.A2(n_729),
.B(n_727),
.C(n_719),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_679),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_686),
.B(n_43),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_682),
.A2(n_92),
.B(n_120),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_682),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_703),
.B(n_44),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_705),
.B(n_45),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_710),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_619),
.B(n_46),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_745),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_620),
.B(n_47),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_664),
.A2(n_49),
.B(n_51),
.C(n_54),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_619),
.B(n_51),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_825),
.A2(n_697),
.B(n_664),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_831),
.A2(n_729),
.B(n_727),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_822),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_937),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_828),
.B(n_777),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_780),
.B(n_747),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_772),
.A2(n_747),
.B1(n_754),
.B2(n_739),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_777),
.B(n_773),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_794),
.B(n_722),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_775),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_827),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_786),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_870),
.A2(n_697),
.B(n_762),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_867),
.A2(n_638),
.B1(n_693),
.B2(n_743),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_780),
.B(n_739),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_776),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_776),
.B(n_786),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_794),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_890),
.B(n_722),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_891),
.A2(n_740),
.B1(n_746),
.B2(n_735),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_776),
.B(n_733),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_834),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_905),
.A2(n_919),
.B1(n_797),
.B2(n_790),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_894),
.A2(n_750),
.B(n_730),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_935),
.B(n_730),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_937),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_930),
.A2(n_701),
.B(n_749),
.C(n_712),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_891),
.A2(n_706),
.B1(n_732),
.B2(n_716),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_901),
.B(n_694),
.Y(n_969)
);

OA22x2_ASAP7_75t_L g970 ( 
.A1(n_895),
.A2(n_694),
.B1(n_732),
.B2(n_716),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_889),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_802),
.A2(n_684),
.B(n_712),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_791),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_798),
.B(n_748),
.Y(n_974)
);

AND2x2_ASAP7_75t_SL g975 ( 
.A(n_936),
.B(n_740),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_912),
.B(n_740),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_862),
.A2(n_740),
.B(n_123),
.Y(n_977)
);

OA22x2_ASAP7_75t_L g978 ( 
.A1(n_908),
.A2(n_926),
.B1(n_830),
.B2(n_899),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_801),
.B(n_883),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_804),
.A2(n_807),
.B(n_859),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_930),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_809),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_888),
.A2(n_934),
.B1(n_785),
.B2(n_874),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_927),
.Y(n_984)
);

INVx6_ASAP7_75t_L g985 ( 
.A(n_791),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_832),
.B(n_833),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_874),
.A2(n_933),
.B(n_934),
.C(n_940),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_776),
.B(n_785),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_835),
.A2(n_866),
.B1(n_868),
.B2(n_836),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_801),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_882),
.B(n_806),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_918),
.A2(n_888),
.B(n_803),
.C(n_838),
.Y(n_992)
);

BUFx2_ASAP7_75t_SL g993 ( 
.A(n_927),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_782),
.B(n_788),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_841),
.B(n_910),
.Y(n_995)
);

AND3x1_ASAP7_75t_SL g996 ( 
.A(n_896),
.B(n_939),
.C(n_906),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_838),
.B(n_839),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_910),
.B(n_881),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_858),
.A2(n_864),
.B(n_863),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_845),
.A2(n_846),
.B(n_848),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_909),
.A2(n_787),
.B(n_783),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_909),
.A2(n_849),
.B(n_820),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_923),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_840),
.A2(n_871),
.B(n_884),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_788),
.B(n_923),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_809),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_892),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_880),
.B(n_896),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_927),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_940),
.A2(n_939),
.B(n_938),
.C(n_903),
.Y(n_1010)
);

CKINVDCx14_ASAP7_75t_R g1011 ( 
.A(n_821),
.Y(n_1011)
);

OR2x4_ASAP7_75t_L g1012 ( 
.A(n_855),
.B(n_904),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_809),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_914),
.B(n_924),
.C(n_928),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_892),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_857),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_837),
.B(n_779),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_927),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_809),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_778),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_915),
.A2(n_893),
.B(n_819),
.C(n_900),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_817),
.A2(n_916),
.B(n_808),
.Y(n_1022)
);

OAI22x1_ASAP7_75t_L g1023 ( 
.A1(n_925),
.A2(n_869),
.B1(n_855),
.B2(n_898),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_850),
.B(n_853),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_900),
.A2(n_843),
.B1(n_815),
.B2(n_844),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_781),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_851),
.A2(n_861),
.B(n_810),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_823),
.B(n_856),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_810),
.A2(n_795),
.B(n_799),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_927),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_902),
.B(n_852),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_SL g1032 ( 
.A1(n_813),
.A2(n_829),
.B1(n_917),
.B2(n_931),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_886),
.A2(n_887),
.B(n_819),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_885),
.A2(n_792),
.B(n_878),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_823),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_823),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_817),
.A2(n_814),
.B(n_913),
.C(n_808),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_771),
.B(n_875),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_793),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_784),
.A2(n_800),
.B(n_847),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_816),
.A2(n_774),
.B(n_913),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_823),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_847),
.A2(n_860),
.B(n_879),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_860),
.A2(n_879),
.B(n_873),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_771),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_805),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_842),
.B(n_875),
.Y(n_1047)
);

XNOR2xp5_ASAP7_75t_L g1048 ( 
.A(n_812),
.B(n_813),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_873),
.A2(n_796),
.B(n_876),
.Y(n_1049)
);

AND2x6_ASAP7_75t_L g1050 ( 
.A(n_856),
.B(n_872),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_842),
.B(n_865),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_818),
.A2(n_824),
.B(n_920),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_856),
.B(n_907),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_818),
.A2(n_922),
.B(n_907),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_916),
.A2(n_897),
.B(n_854),
.C(n_826),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_856),
.B(n_907),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_865),
.A2(n_872),
.B1(n_911),
.B2(n_929),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_865),
.A2(n_872),
.B1(n_911),
.B2(n_932),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_811),
.A2(n_789),
.B(n_877),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_921),
.B(n_579),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_921),
.A2(n_612),
.B(n_608),
.C(n_919),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_919),
.A2(n_612),
.B(n_608),
.C(n_688),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_828),
.B(n_612),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_772),
.A2(n_588),
.B1(n_479),
.B2(n_633),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_825),
.A2(n_870),
.B(n_894),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_891),
.A2(n_447),
.B(n_434),
.C(n_469),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_SL g1067 ( 
.A(n_822),
.B(n_487),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_825),
.A2(n_870),
.B(n_894),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_775),
.B(n_617),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_775),
.B(n_617),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_905),
.A2(n_617),
.B1(n_635),
.B2(n_474),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_905),
.A2(n_617),
.B1(n_635),
.B2(n_474),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_827),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_930),
.A2(n_891),
.B(n_934),
.C(n_777),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_905),
.A2(n_635),
.B1(n_617),
.B2(n_474),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_772),
.B(n_672),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_825),
.A2(n_870),
.B(n_894),
.Y(n_1077)
);

BUFx8_ASAP7_75t_L g1078 ( 
.A(n_822),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_780),
.B(n_791),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_772),
.B(n_672),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_825),
.A2(n_870),
.B(n_894),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_919),
.A2(n_612),
.B(n_608),
.C(n_688),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_1074),
.A2(n_1063),
.B1(n_1023),
.B2(n_992),
.C(n_945),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_948),
.B(n_981),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1010),
.A2(n_997),
.B(n_1061),
.C(n_963),
.Y(n_1086)
);

AOI221x1_ASAP7_75t_L g1087 ( 
.A1(n_1014),
.A2(n_1075),
.B1(n_1072),
.B2(n_1071),
.C(n_941),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1000),
.A2(n_999),
.B(n_980),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1052),
.A2(n_1081),
.B(n_1077),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_1025),
.A2(n_1068),
.A3(n_1065),
.B(n_1033),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_953),
.A2(n_1002),
.B(n_988),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1054),
.A2(n_964),
.B(n_1027),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_1041),
.A2(n_1059),
.B(n_1029),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1009),
.A2(n_975),
.B1(n_994),
.B2(n_984),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_1035),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_977),
.A2(n_1041),
.B(n_1049),
.Y(n_1096)
);

NAND3x1_ASAP7_75t_L g1097 ( 
.A(n_971),
.B(n_979),
.C(n_1011),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1024),
.B(n_974),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_951),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_998),
.B(n_959),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1026),
.Y(n_1101)
);

NAND3xp33_ASAP7_75t_L g1102 ( 
.A(n_1066),
.B(n_1037),
.C(n_960),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1034),
.A2(n_1021),
.B(n_967),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_984),
.B(n_1009),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1039),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1044),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1050),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_950),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1055),
.A2(n_995),
.B(n_1032),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1046),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_955),
.A2(n_965),
.B(n_947),
.C(n_976),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_972),
.A2(n_984),
.B(n_961),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_942),
.A2(n_1058),
.B(n_1057),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_973),
.B(n_944),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_969),
.B(n_991),
.Y(n_1115)
);

CKINVDCx6p67_ASAP7_75t_R g1116 ( 
.A(n_943),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_952),
.Y(n_1117)
);

AOI221x1_ASAP7_75t_L g1118 ( 
.A1(n_954),
.A2(n_1057),
.B1(n_1058),
.B2(n_1005),
.C(n_1008),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_1067),
.B(n_1022),
.C(n_989),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1003),
.B(n_978),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1064),
.A2(n_990),
.B1(n_1012),
.B2(n_1080),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1076),
.B(n_958),
.Y(n_1122)
);

AO32x2_ASAP7_75t_L g1123 ( 
.A1(n_978),
.A2(n_996),
.A3(n_1006),
.B1(n_1036),
.B2(n_1012),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1053),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_970),
.A2(n_1056),
.B(n_957),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_958),
.B(n_1073),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1018),
.A2(n_962),
.B(n_949),
.C(n_1030),
.Y(n_1127)
);

CKINVDCx14_ASAP7_75t_R g1128 ( 
.A(n_985),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1069),
.A2(n_1070),
.B(n_1045),
.C(n_966),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_982),
.Y(n_1130)
);

INVx3_ASAP7_75t_SL g1131 ( 
.A(n_985),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1016),
.B(n_944),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1078),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1048),
.A2(n_1051),
.B(n_1047),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_966),
.B(n_1007),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1079),
.B(n_946),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1038),
.A2(n_1007),
.B(n_993),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_956),
.A2(n_1006),
.A3(n_986),
.B(n_946),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_956),
.A2(n_1050),
.B(n_986),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_986),
.A2(n_946),
.A3(n_1050),
.B(n_1013),
.Y(n_1140)
);

CKINVDCx11_ASAP7_75t_R g1141 ( 
.A(n_1079),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1050),
.A2(n_982),
.B(n_1013),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1015),
.B(n_1078),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1042),
.A2(n_982),
.B(n_1013),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1019),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1074),
.A2(n_983),
.B(n_997),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_1023),
.A2(n_862),
.A3(n_789),
.B(n_1060),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1150)
);

AOI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1074),
.A2(n_612),
.B1(n_688),
.B2(n_633),
.C(n_1062),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1154)
);

OAI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_983),
.A2(n_1074),
.B(n_612),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_948),
.B(n_997),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1020),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_951),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_982),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1078),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1074),
.A2(n_612),
.B1(n_688),
.B2(n_633),
.C(n_1062),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1063),
.A2(n_633),
.B1(n_612),
.B2(n_479),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_951),
.Y(n_1170)
);

AO32x2_ASAP7_75t_L g1171 ( 
.A1(n_963),
.A2(n_968),
.A3(n_1075),
.B1(n_1072),
.B2(n_1071),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_951),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_952),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_948),
.B(n_612),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_1078),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1074),
.A2(n_983),
.B(n_997),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1074),
.A2(n_983),
.B(n_997),
.Y(n_1178)
);

OAI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_983),
.A2(n_612),
.B1(n_1074),
.B2(n_688),
.C(n_633),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1041),
.A2(n_1000),
.B(n_1004),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_948),
.B(n_997),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_1075),
.A2(n_1072),
.B1(n_1071),
.B2(n_945),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1078),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1074),
.A2(n_983),
.B(n_997),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1187)
);

AOI31xp67_ASAP7_75t_L g1188 ( 
.A1(n_983),
.A2(n_1060),
.A3(n_792),
.B(n_960),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_948),
.B(n_997),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_990),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1059),
.A2(n_977),
.B(n_1065),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1063),
.A2(n_633),
.B1(n_612),
.B2(n_479),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_948),
.B(n_997),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_985),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_983),
.A2(n_1074),
.B1(n_997),
.B2(n_981),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1197)
);

NOR4xp25_ASAP7_75t_L g1198 ( 
.A(n_1074),
.B(n_987),
.C(n_1082),
.D(n_1062),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1074),
.A2(n_983),
.B(n_997),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_L g1202 ( 
.A1(n_1063),
.A2(n_828),
.B(n_1074),
.C(n_919),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_948),
.B(n_997),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1076),
.B(n_1080),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_952),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_948),
.B(n_672),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1004),
.A2(n_1040),
.B(n_1001),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1023),
.A2(n_862),
.A3(n_789),
.B(n_1060),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1076),
.B(n_772),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1076),
.B(n_772),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_948),
.B(n_997),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1074),
.A2(n_983),
.B(n_997),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_990),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_948),
.B(n_997),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1020),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_941),
.A2(n_1068),
.B(n_1065),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1161),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1174),
.A2(n_1147),
.B1(n_1186),
.B2(n_1178),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1121),
.A2(n_1177),
.B1(n_1186),
.B2(n_1178),
.Y(n_1224)
);

INVx8_ASAP7_75t_L g1225 ( 
.A(n_1175),
.Y(n_1225)
);

BUFx4f_ASAP7_75t_SL g1226 ( 
.A(n_1116),
.Y(n_1226)
);

INVx8_ASAP7_75t_L g1227 ( 
.A(n_1136),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1147),
.A2(n_1200),
.B1(n_1177),
.B2(n_1217),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1200),
.A2(n_1217),
.B1(n_1193),
.B2(n_1167),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1133),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1099),
.Y(n_1231)
);

INVx6_ASAP7_75t_L g1232 ( 
.A(n_1107),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1141),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1196),
.A2(n_1184),
.B1(n_1203),
.B2(n_1156),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1156),
.B(n_1183),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1196),
.A2(n_1184),
.B1(n_1189),
.B2(n_1194),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1194),
.A2(n_1203),
.B1(n_1216),
.B2(n_1219),
.Y(n_1237)
);

BUFx8_ASAP7_75t_L g1238 ( 
.A(n_1191),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1158),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1095),
.Y(n_1240)
);

CKINVDCx8_ASAP7_75t_R g1241 ( 
.A(n_1108),
.Y(n_1241)
);

INVx6_ASAP7_75t_L g1242 ( 
.A(n_1136),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1086),
.A2(n_1221),
.B(n_1212),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1213),
.A2(n_1215),
.B1(n_1085),
.B2(n_1207),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1098),
.B(n_1205),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1117),
.Y(n_1247)
);

INVx8_ASAP7_75t_L g1248 ( 
.A(n_1130),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1172),
.Y(n_1249)
);

BUFx2_ASAP7_75t_R g1250 ( 
.A(n_1185),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1130),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1098),
.A2(n_1120),
.B1(n_1100),
.B2(n_1122),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1126),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1195),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1094),
.A2(n_1119),
.B1(n_1120),
.B2(n_1109),
.Y(n_1255)
);

INVx6_ASAP7_75t_L g1256 ( 
.A(n_1160),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1083),
.A2(n_1118),
.B1(n_1087),
.B2(n_1100),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1140),
.B(n_1138),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1160),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1115),
.A2(n_1134),
.B1(n_1102),
.B2(n_1094),
.Y(n_1260)
);

CKINVDCx6p67_ASAP7_75t_R g1261 ( 
.A(n_1143),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1102),
.A2(n_1171),
.B1(n_1115),
.B2(n_1103),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1145),
.Y(n_1263)
);

BUFx2_ASAP7_75t_SL g1264 ( 
.A(n_1114),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1101),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1104),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1173),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1206),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1218),
.A2(n_1110),
.B1(n_1214),
.B2(n_1105),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1128),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1145),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_1097),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1157),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1111),
.A2(n_1132),
.B1(n_1103),
.B2(n_1129),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1220),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1123),
.B(n_1198),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1123),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1144),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1171),
.A2(n_1202),
.B1(n_1124),
.B2(n_1135),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1142),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1138),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1139),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1106),
.A2(n_1125),
.B1(n_1093),
.B2(n_1091),
.Y(n_1283)
);

BUFx8_ASAP7_75t_SL g1284 ( 
.A(n_1192),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_SL g1285 ( 
.A(n_1188),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1127),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1149),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1150),
.A2(n_1201),
.B(n_1210),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1211),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1112),
.A2(n_1093),
.B1(n_1092),
.B2(n_1204),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1137),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_1211),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1113),
.A2(n_1096),
.B1(n_1199),
.B2(n_1169),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1209),
.A2(n_1164),
.B1(n_1197),
.B2(n_1165),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1089),
.A2(n_1180),
.B1(n_1187),
.B2(n_1159),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1153),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1090),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1154),
.A2(n_1176),
.B1(n_1168),
.B2(n_1180),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1088),
.B(n_1084),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1146),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1148),
.Y(n_1301)
);

BUFx8_ASAP7_75t_SL g1302 ( 
.A(n_1152),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1163),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1181),
.A2(n_1182),
.B1(n_1190),
.B2(n_1208),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1131),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1131),
.Y(n_1307)
);

BUFx12f_ASAP7_75t_L g1308 ( 
.A(n_1133),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_L g1309 ( 
.A(n_1161),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1179),
.A2(n_1155),
.B1(n_1151),
.B2(n_1166),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1099),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1179),
.A2(n_1155),
.B1(n_1151),
.B2(n_1166),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1179),
.A2(n_1155),
.B1(n_1151),
.B2(n_1166),
.Y(n_1313)
);

CKINVDCx6p67_ASAP7_75t_R g1314 ( 
.A(n_1161),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1133),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1099),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1099),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1156),
.B(n_1183),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1179),
.A2(n_1155),
.B1(n_1151),
.B2(n_1166),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1179),
.A2(n_983),
.B1(n_1166),
.B2(n_1151),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1179),
.A2(n_983),
.B1(n_1166),
.B2(n_1151),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1099),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1099),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1320),
.A2(n_1321),
.B1(n_1229),
.B2(n_1224),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1276),
.B(n_1228),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1228),
.B(n_1277),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1231),
.B(n_1239),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1223),
.A2(n_1229),
.B1(n_1312),
.B2(n_1319),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1247),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1303),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1273),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1303),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1302),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1282),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1267),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1237),
.B(n_1223),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1287),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1289),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1237),
.B(n_1234),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1291),
.B(n_1258),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1243),
.A2(n_1299),
.B(n_1293),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1234),
.B(n_1236),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1293),
.A2(n_1298),
.B(n_1305),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1282),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1298),
.A2(n_1305),
.B(n_1283),
.Y(n_1346)
);

BUFx4f_ASAP7_75t_SL g1347 ( 
.A(n_1230),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1273),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1323),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1246),
.B(n_1236),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1302),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1283),
.A2(n_1288),
.B(n_1300),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_SL g1353 ( 
.A(n_1241),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1280),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1311),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1322),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1316),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1222),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1317),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1290),
.A2(n_1257),
.B(n_1294),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1268),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1296),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1292),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1278),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1292),
.Y(n_1365)
);

BUFx12f_ASAP7_75t_L g1366 ( 
.A(n_1222),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1286),
.A2(n_1274),
.B(n_1253),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1271),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1262),
.B(n_1297),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1281),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1284),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1235),
.A2(n_1318),
.B1(n_1285),
.B2(n_1240),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_1270),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1245),
.B(n_1252),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1297),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1245),
.B(n_1252),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1265),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1284),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1285),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1304),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1255),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1301),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1330),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1349),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1349),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1324),
.A2(n_1313),
.B(n_1310),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1329),
.A2(n_1260),
.B(n_1295),
.Y(n_1387)
);

AO21x1_ASAP7_75t_L g1388 ( 
.A1(n_1337),
.A2(n_1263),
.B(n_1259),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1324),
.A2(n_1260),
.B(n_1279),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1334),
.B(n_1307),
.Y(n_1390)
);

AO21x1_ASAP7_75t_L g1391 ( 
.A1(n_1381),
.A2(n_1263),
.B(n_1259),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1352),
.A2(n_1269),
.B(n_1306),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_R g1393 ( 
.A(n_1358),
.B(n_1233),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1325),
.B(n_1254),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1364),
.B(n_1326),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1334),
.B(n_1227),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1351),
.B(n_1233),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1361),
.B(n_1238),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1340),
.A2(n_1266),
.B(n_1264),
.C(n_1226),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1336),
.B(n_1238),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1362),
.B(n_1261),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1343),
.A2(n_1309),
.B(n_1227),
.C(n_1225),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_R g1403 ( 
.A(n_1351),
.B(n_1371),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1362),
.B(n_1275),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1327),
.B(n_1250),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1355),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1355),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1366),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1369),
.A2(n_1272),
.B1(n_1232),
.B2(n_1242),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1351),
.B(n_1272),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1327),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1331),
.B(n_1272),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1328),
.B(n_1251),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1329),
.A2(n_1242),
.B1(n_1314),
.B2(n_1225),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1369),
.A2(n_1242),
.B1(n_1225),
.B2(n_1230),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1328),
.B(n_1256),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1356),
.Y(n_1417)
);

BUFx2_ASAP7_75t_SL g1418 ( 
.A(n_1332),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1374),
.A2(n_1248),
.B(n_1226),
.C(n_1308),
.Y(n_1419)
);

BUFx2_ASAP7_75t_SL g1420 ( 
.A(n_1348),
.Y(n_1420)
);

AO32x2_ASAP7_75t_L g1421 ( 
.A1(n_1335),
.A2(n_1308),
.A3(n_1315),
.B1(n_1345),
.B2(n_1368),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1378),
.B(n_1326),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1331),
.B(n_1333),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1380),
.B(n_1375),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1353),
.B(n_1347),
.Y(n_1425)
);

AOI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1372),
.A2(n_1367),
.B1(n_1376),
.B2(n_1374),
.C(n_1357),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1359),
.B(n_1350),
.Y(n_1427)
);

OAI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1379),
.A2(n_1333),
.B1(n_1331),
.B2(n_1365),
.C(n_1363),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1366),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1375),
.B(n_1377),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1383),
.B(n_1411),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1395),
.B(n_1367),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1423),
.B(n_1331),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1428),
.B(n_1360),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1384),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1385),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1406),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1422),
.B(n_1354),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1386),
.A2(n_1387),
.B1(n_1389),
.B2(n_1414),
.Y(n_1439)
);

AND2x2_ASAP7_75t_SL g1440 ( 
.A(n_1426),
.B(n_1341),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1407),
.Y(n_1441)
);

INVxp67_ASAP7_75t_SL g1442 ( 
.A(n_1395),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1389),
.A2(n_1360),
.B1(n_1370),
.B2(n_1341),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1417),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1430),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1427),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1424),
.B(n_1382),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1394),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1413),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1392),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1392),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1416),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1421),
.B(n_1382),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_L g1454 ( 
.A(n_1396),
.B(n_1410),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1421),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1421),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1393),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1448),
.B(n_1346),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1439),
.A2(n_1405),
.B1(n_1414),
.B2(n_1404),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1432),
.B(n_1342),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1442),
.B(n_1344),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1446),
.B(n_1342),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1435),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1440),
.A2(n_1408),
.B1(n_1415),
.B2(n_1401),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1457),
.B(n_1418),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1440),
.A2(n_1415),
.B1(n_1403),
.B2(n_1402),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1443),
.A2(n_1399),
.B1(n_1419),
.B2(n_1388),
.C(n_1420),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1449),
.B(n_1344),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1435),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1454),
.B(n_1433),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1454),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1453),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1455),
.A2(n_1410),
.B(n_1396),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1434),
.B(n_1436),
.Y(n_1474)
);

INVx5_ASAP7_75t_L g1475 ( 
.A(n_1453),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1440),
.A2(n_1409),
.B1(n_1412),
.B2(n_1397),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1450),
.A2(n_1338),
.B(n_1339),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1434),
.A2(n_1412),
.B1(n_1365),
.B2(n_1391),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1437),
.B(n_1441),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1456),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1472),
.B(n_1438),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1472),
.B(n_1438),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1477),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1477),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1486)
);

NAND2xp33_ASAP7_75t_R g1487 ( 
.A(n_1470),
.B(n_1429),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1477),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1472),
.B(n_1452),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1463),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1473),
.B(n_1450),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1474),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1480),
.B(n_1446),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1463),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1463),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1477),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1480),
.B(n_1431),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1468),
.B(n_1444),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1462),
.B(n_1474),
.Y(n_1501)
);

NAND2xp33_ASAP7_75t_R g1502 ( 
.A(n_1470),
.B(n_1451),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1469),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1477),
.Y(n_1504)
);

NOR3xp33_ASAP7_75t_SL g1505 ( 
.A(n_1465),
.B(n_1425),
.C(n_1400),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1475),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1469),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1475),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1462),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1475),
.B(n_1433),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1475),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1492),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1483),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1492),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1505),
.A2(n_1478),
.B(n_1467),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1492),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1483),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1496),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1505),
.Y(n_1520)
);

NOR2x1_ASAP7_75t_L g1521 ( 
.A(n_1506),
.B(n_1465),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1496),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1499),
.B(n_1474),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1483),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1494),
.B(n_1468),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1499),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1470),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1481),
.B(n_1470),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1482),
.B(n_1470),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1494),
.B(n_1468),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1482),
.B(n_1485),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1483),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1495),
.B(n_1462),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1500),
.B(n_1468),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1500),
.B(n_1461),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_SL g1537 ( 
.A(n_1508),
.B(n_1471),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1510),
.A2(n_1461),
.B(n_1467),
.C(n_1478),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1495),
.B(n_1460),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1501),
.B(n_1373),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1484),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1495),
.B(n_1460),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1510),
.B(n_1461),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1487),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1501),
.B(n_1461),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1501),
.B(n_1458),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1497),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1484),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1491),
.B(n_1458),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1503),
.B(n_1460),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1503),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1526),
.B(n_1503),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1516),
.B(n_1507),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1538),
.B(n_1507),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_1540),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1521),
.B(n_1482),
.Y(n_1556)
);

AND3x1_ASAP7_75t_L g1557 ( 
.A(n_1512),
.B(n_1506),
.C(n_1508),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1544),
.B(n_1485),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1532),
.B(n_1485),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1507),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1532),
.B(n_1486),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1523),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1525),
.A2(n_1459),
.B(n_1466),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1527),
.B(n_1486),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1460),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1527),
.B(n_1486),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1528),
.B(n_1491),
.Y(n_1567)
);

AND2x4_ASAP7_75t_SL g1568 ( 
.A(n_1512),
.B(n_1506),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1539),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1515),
.Y(n_1570)
);

INVxp33_ASAP7_75t_L g1571 ( 
.A(n_1545),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1542),
.B(n_1509),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1515),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1550),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1509),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1528),
.B(n_1491),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1514),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1529),
.B(n_1508),
.Y(n_1578)
);

NOR3xp33_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1467),
.C(n_1484),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1513),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1519),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1517),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1550),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1546),
.B(n_1509),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1517),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1529),
.B(n_1488),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1562),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1580),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1530),
.C(n_1531),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1553),
.A2(n_1498),
.B1(n_1484),
.B2(n_1504),
.C(n_1490),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1570),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1570),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1562),
.B(n_1549),
.Y(n_1594)
);

AOI322xp5_ASAP7_75t_L g1595 ( 
.A1(n_1554),
.A2(n_1536),
.A3(n_1498),
.B1(n_1504),
.B2(n_1490),
.C1(n_1459),
.C2(n_1535),
.Y(n_1595)
);

NAND4xp75_ASAP7_75t_L g1596 ( 
.A(n_1557),
.B(n_1466),
.C(n_1508),
.D(n_1498),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1583),
.B(n_1458),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1574),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_1555),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1573),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1557),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1604)
);

NAND2x1_ASAP7_75t_L g1605 ( 
.A(n_1556),
.B(n_1578),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1511),
.Y(n_1606)
);

AOI322xp5_ASAP7_75t_L g1607 ( 
.A1(n_1579),
.A2(n_1490),
.A3(n_1498),
.B1(n_1504),
.B2(n_1464),
.C1(n_1476),
.C2(n_1458),
.Y(n_1607)
);

INVxp33_ASAP7_75t_L g1608 ( 
.A(n_1563),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1573),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1583),
.B(n_1534),
.Y(n_1610)
);

OAI32xp33_ASAP7_75t_L g1611 ( 
.A1(n_1563),
.A2(n_1502),
.A3(n_1487),
.B1(n_1534),
.B2(n_1506),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1574),
.B(n_1488),
.Y(n_1612)
);

OAI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1571),
.A2(n_1489),
.B(n_1488),
.Y(n_1613)
);

AOI221x1_ASAP7_75t_L g1614 ( 
.A1(n_1589),
.A2(n_1552),
.B1(n_1537),
.B2(n_1585),
.C(n_1582),
.Y(n_1614)
);

AOI221x1_ASAP7_75t_L g1615 ( 
.A1(n_1598),
.A2(n_1552),
.B1(n_1537),
.B2(n_1585),
.C(n_1582),
.Y(n_1615)
);

AOI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1608),
.A2(n_1569),
.B(n_1577),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1602),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1605),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1592),
.Y(n_1620)
);

OAI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1599),
.A2(n_1556),
.B(n_1584),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_SL g1622 ( 
.A1(n_1588),
.A2(n_1581),
.B(n_1560),
.C(n_1575),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1593),
.Y(n_1623)
);

OAI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1602),
.A2(n_1502),
.B1(n_1504),
.B2(n_1490),
.C(n_1493),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1608),
.A2(n_1577),
.B1(n_1548),
.B2(n_1518),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1600),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1596),
.A2(n_1565),
.B(n_1493),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1609),
.Y(n_1628)
);

OAI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1604),
.A2(n_1584),
.B(n_1565),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1598),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1561),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1603),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1590),
.B1(n_1601),
.B2(n_1594),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1633),
.B(n_1610),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1618),
.B(n_1606),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1633),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1633),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1631),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1631),
.B(n_1606),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1622),
.A2(n_1611),
.B1(n_1617),
.B2(n_1627),
.C(n_1624),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1632),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_L g1644 ( 
.A(n_1621),
.B(n_1612),
.Y(n_1644)
);

AOI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1642),
.A2(n_1622),
.B(n_1617),
.C(n_1630),
.Y(n_1645)
);

NOR3xp33_ASAP7_75t_L g1646 ( 
.A(n_1643),
.B(n_1623),
.C(n_1620),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1636),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1635),
.A2(n_1614),
.B(n_1615),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1638),
.Y(n_1649)
);

NOR2xp67_ASAP7_75t_L g1650 ( 
.A(n_1640),
.B(n_1619),
.Y(n_1650)
);

NOR4xp25_ASAP7_75t_L g1651 ( 
.A(n_1639),
.B(n_1628),
.C(n_1626),
.D(n_1625),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1641),
.B(n_1629),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1634),
.B(n_1597),
.Y(n_1653)
);

INVxp67_ASAP7_75t_SL g1654 ( 
.A(n_1637),
.Y(n_1654)
);

AOI222xp33_ASAP7_75t_L g1655 ( 
.A1(n_1648),
.A2(n_1591),
.B1(n_1644),
.B2(n_1577),
.C1(n_1614),
.C2(n_1615),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1645),
.A2(n_1634),
.B(n_1619),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1651),
.A2(n_1612),
.B1(n_1595),
.B2(n_1524),
.C(n_1518),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1647),
.B(n_1649),
.Y(n_1658)
);

XOR2xp5_ASAP7_75t_L g1659 ( 
.A(n_1652),
.B(n_1398),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1657),
.A2(n_1651),
.B1(n_1653),
.B2(n_1646),
.C(n_1654),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1656),
.A2(n_1524),
.B1(n_1514),
.B2(n_1533),
.C(n_1541),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1658),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1659),
.Y(n_1663)
);

XOR2x2_ASAP7_75t_L g1664 ( 
.A(n_1655),
.B(n_1650),
.Y(n_1664)
);

O2A1O1Ixp5_ASAP7_75t_L g1665 ( 
.A1(n_1656),
.A2(n_1560),
.B(n_1575),
.C(n_1578),
.Y(n_1665)
);

NAND4xp75_ASAP7_75t_L g1666 ( 
.A(n_1660),
.B(n_1564),
.C(n_1566),
.D(n_1576),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1662),
.B(n_1607),
.Y(n_1667)
);

NAND4xp75_ASAP7_75t_L g1668 ( 
.A(n_1663),
.B(n_1566),
.C(n_1564),
.D(n_1576),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1664),
.B(n_1572),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1665),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1669),
.B(n_1587),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1670),
.B(n_1667),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1671),
.Y(n_1674)
);

AO22x2_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1672),
.B1(n_1666),
.B2(n_1673),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1675),
.B(n_1672),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1675),
.Y(n_1677)
);

OR3x1_ASAP7_75t_L g1678 ( 
.A(n_1677),
.B(n_1672),
.C(n_1373),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1676),
.B(n_1572),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1678),
.A2(n_1661),
.B1(n_1578),
.B2(n_1568),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1679),
.A2(n_1578),
.B1(n_1586),
.B2(n_1522),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1680),
.A2(n_1681),
.B1(n_1568),
.B2(n_1613),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1541),
.B(n_1533),
.Y(n_1683)
);

XNOR2xp5_ASAP7_75t_L g1684 ( 
.A(n_1683),
.B(n_1390),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_R g1685 ( 
.A1(n_1684),
.A2(n_1568),
.B1(n_1586),
.B2(n_1567),
.C(n_1464),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1567),
.B1(n_1551),
.B2(n_1547),
.Y(n_1686)
);


endmodule