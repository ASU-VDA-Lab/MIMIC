module real_aes_867_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g600 ( .A(n_0), .B(n_170), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_1), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g131 ( .A(n_2), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_3), .B(n_537), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g592 ( .A(n_4), .B(n_152), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_5), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g585 ( .A(n_6), .Y(n_585) );
INVx1_ASAP7_75t_L g192 ( .A(n_7), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_8), .Y(n_499) );
AOI22xp5_ASAP7_75t_SL g829 ( .A1(n_9), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_9), .Y(n_830) );
OAI22x1_ASAP7_75t_R g832 ( .A1(n_10), .A2(n_80), .B1(n_833), .B2(n_834), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_10), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_11), .Y(n_208) );
AND2x2_ASAP7_75t_L g534 ( .A(n_12), .B(n_121), .Y(n_534) );
INVx2_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_14), .Y(n_484) );
INVx1_ASAP7_75t_L g171 ( .A(n_15), .Y(n_171) );
AOI221x1_ASAP7_75t_L g588 ( .A1(n_16), .A2(n_154), .B1(n_539), .B2(n_589), .C(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g842 ( .A(n_17), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_18), .B(n_537), .Y(n_572) );
INVx1_ASAP7_75t_L g488 ( .A(n_19), .Y(n_488) );
INVx1_ASAP7_75t_L g168 ( .A(n_20), .Y(n_168) );
INVx1_ASAP7_75t_SL g143 ( .A(n_21), .Y(n_143) );
AND2x2_ASAP7_75t_L g491 ( .A(n_22), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_23), .B(n_146), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_24), .A2(n_31), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_24), .Y(n_478) );
AOI33xp33_ASAP7_75t_L g220 ( .A1(n_25), .A2(n_55), .A3(n_128), .B1(n_139), .B2(n_221), .B3(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_26), .A2(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_27), .B(n_170), .Y(n_541) );
AOI221xp5_ASAP7_75t_SL g564 ( .A1(n_28), .A2(n_46), .B1(n_537), .B2(n_539), .C(n_565), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_29), .A2(n_64), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g201 ( .A(n_30), .Y(n_201) );
INVx1_ASAP7_75t_SL g479 ( .A(n_31), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_31), .B(n_113), .C(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g123 ( .A(n_32), .B(n_92), .Y(n_123) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_32), .A2(n_92), .B(n_122), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_33), .B(n_173), .Y(n_576) );
INVxp67_ASAP7_75t_L g587 ( .A(n_34), .Y(n_587) );
AND2x2_ASAP7_75t_L g560 ( .A(n_35), .B(n_120), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_36), .B(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_37), .A2(n_539), .B(n_599), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_38), .B(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_39), .B(n_173), .Y(n_566) );
AND2x2_ASAP7_75t_L g133 ( .A(n_40), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g138 ( .A(n_40), .Y(n_138) );
AND2x2_ASAP7_75t_L g152 ( .A(n_40), .B(n_131), .Y(n_152) );
OR2x6_ASAP7_75t_L g486 ( .A(n_41), .B(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_42), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_43), .B(n_126), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_44), .A2(n_155), .B1(n_161), .B2(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_45), .B(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_47), .A2(n_84), .B1(n_136), .B2(n_539), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_48), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_49), .B(n_170), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_50), .B(n_189), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_51), .B(n_146), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_52), .Y(n_249) );
AND2x2_ASAP7_75t_L g603 ( .A(n_53), .B(n_120), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_54), .B(n_120), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_56), .B(n_146), .Y(n_232) );
INVx1_ASAP7_75t_L g129 ( .A(n_57), .Y(n_129) );
INVx1_ASAP7_75t_L g148 ( .A(n_57), .Y(n_148) );
AND2x2_ASAP7_75t_L g233 ( .A(n_58), .B(n_120), .Y(n_233) );
AOI221xp5_ASAP7_75t_L g190 ( .A1(n_59), .A2(n_76), .B1(n_126), .B2(n_136), .C(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_60), .B(n_126), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_61), .B(n_537), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_62), .B(n_155), .Y(n_210) );
AOI21xp5_ASAP7_75t_SL g180 ( .A1(n_63), .A2(n_136), .B(n_181), .Y(n_180) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_64), .A2(n_105), .B1(n_494), .B2(n_501), .C(n_510), .Y(n_104) );
INVxp67_ASAP7_75t_L g109 ( .A(n_64), .Y(n_109) );
AND2x2_ASAP7_75t_L g551 ( .A(n_64), .B(n_120), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_65), .B(n_173), .Y(n_601) );
INVx1_ASAP7_75t_L g164 ( .A(n_66), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_67), .B(n_170), .Y(n_549) );
AND2x2_ASAP7_75t_SL g577 ( .A(n_68), .B(n_121), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_69), .A2(n_539), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g231 ( .A(n_70), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_71), .B(n_173), .Y(n_542) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_72), .B(n_189), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_73), .A2(n_136), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g134 ( .A(n_74), .Y(n_134) );
INVx1_ASAP7_75t_L g150 ( .A(n_74), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_75), .B(n_126), .Y(n_223) );
AND2x2_ASAP7_75t_L g153 ( .A(n_77), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g165 ( .A(n_78), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_79), .A2(n_136), .B(n_142), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_80), .Y(n_834) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_81), .A2(n_136), .B(n_215), .C(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_82), .B(n_537), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_83), .A2(n_87), .B1(n_126), .B2(n_537), .Y(n_613) );
INVx1_ASAP7_75t_L g489 ( .A(n_85), .Y(n_489) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_86), .B(n_154), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_88), .A2(n_136), .B1(n_218), .B2(n_219), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_89), .B(n_170), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_90), .B(n_170), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_91), .A2(n_539), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g182 ( .A(n_93), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_94), .B(n_173), .Y(n_548) );
AND2x2_ASAP7_75t_L g224 ( .A(n_95), .B(n_154), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_96), .A2(n_199), .B(n_200), .C(n_202), .Y(n_198) );
INVxp67_ASAP7_75t_L g590 ( .A(n_97), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_98), .B(n_537), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_99), .B(n_173), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_100), .A2(n_539), .B(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g500 ( .A(n_101), .Y(n_500) );
BUFx2_ASAP7_75t_SL g507 ( .A(n_101), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_102), .B(n_146), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_103), .A2(n_476), .B1(n_477), .B2(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_103), .Y(n_476) );
OAI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_481), .B(n_490), .Y(n_105) );
XOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_112), .B1(n_474), .B2(n_475), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR3x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_339), .C(n_410), .Y(n_112) );
INVx1_ASAP7_75t_L g525 ( .A(n_113), .Y(n_525) );
NAND3x1_ASAP7_75t_SL g113 ( .A(n_114), .B(n_266), .C(n_288), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_256), .Y(n_114) );
AOI22xp33_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_185), .B1(n_234), .B2(n_238), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_116), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_441) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_157), .Y(n_116) );
AND2x2_ASAP7_75t_L g257 ( .A(n_117), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_117), .B(n_304), .Y(n_323) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g241 ( .A(n_118), .Y(n_241) );
AND2x2_ASAP7_75t_L g291 ( .A(n_118), .B(n_159), .Y(n_291) );
INVx1_ASAP7_75t_L g330 ( .A(n_118), .Y(n_330) );
OR2x2_ASAP7_75t_L g367 ( .A(n_118), .B(n_177), .Y(n_367) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_118), .Y(n_379) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_118), .Y(n_403) );
AND2x2_ASAP7_75t_L g460 ( .A(n_118), .B(n_287), .Y(n_460) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_153), .Y(n_118) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_119), .A2(n_545), .B(n_551), .Y(n_544) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_119), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x2_ASAP7_75t_L g692 ( .A1(n_119), .A2(n_554), .B(n_560), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
OA21x2_ASAP7_75t_L g563 ( .A1(n_120), .A2(n_564), .B(n_568), .Y(n_563) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x4_ASAP7_75t_L g161 ( .A(n_122), .B(n_123), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_135), .Y(n_124) );
INVx1_ASAP7_75t_L g211 ( .A(n_126), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_126), .A2(n_136), .B1(n_584), .B2(n_586), .Y(n_583) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
INVx1_ASAP7_75t_L g247 ( .A(n_127), .Y(n_247) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
OR2x6_ASAP7_75t_L g144 ( .A(n_128), .B(n_140), .Y(n_144) );
INVxp33_ASAP7_75t_L g221 ( .A(n_128), .Y(n_221) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g141 ( .A(n_129), .B(n_131), .Y(n_141) );
AND2x4_ASAP7_75t_L g173 ( .A(n_129), .B(n_149), .Y(n_173) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g248 ( .A(n_132), .Y(n_248) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_L g539 ( .A(n_133), .B(n_141), .Y(n_539) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
AND2x6_ASAP7_75t_L g170 ( .A(n_134), .B(n_147), .Y(n_170) );
INVxp67_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NOR2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_144), .B(n_145), .C(n_151), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_144), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_144), .A2(n_151), .B(n_182), .C(n_183), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_144), .A2(n_151), .B(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_144), .A2(n_151), .B(n_231), .C(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g254 ( .A(n_144), .Y(n_254) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
AND2x4_ASAP7_75t_L g537 ( .A(n_146), .B(n_152), .Y(n_537) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_151), .B(n_161), .Y(n_174) );
INVx1_ASAP7_75t_L g218 ( .A(n_151), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_151), .A2(n_252), .B(n_253), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_151), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_151), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_151), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_151), .A2(n_566), .B(n_567), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_151), .A2(n_575), .B(n_576), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_151), .A2(n_600), .B(n_601), .Y(n_599) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_154), .A2(n_198), .B1(n_203), .B2(n_204), .Y(n_197) );
INVx3_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_155), .B(n_207), .Y(n_206) );
AOI21x1_ASAP7_75t_L g596 ( .A1(n_155), .A2(n_597), .B(n_603), .Y(n_596) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
NOR2x1_ASAP7_75t_L g157 ( .A(n_158), .B(n_175), .Y(n_157) );
INVx1_ASAP7_75t_L g335 ( .A(n_158), .Y(n_335) );
AND2x2_ASAP7_75t_L g361 ( .A(n_158), .B(n_177), .Y(n_361) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_158), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g258 ( .A(n_159), .B(n_244), .Y(n_258) );
INVx3_ASAP7_75t_L g287 ( .A(n_159), .Y(n_287) );
NOR2x1_ASAP7_75t_SL g406 ( .A(n_159), .B(n_177), .Y(n_406) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_161), .A2(n_180), .B(n_184), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_161), .A2(n_536), .B(n_538), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_161), .B(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_161), .B(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_161), .B(n_590), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_161), .B(n_166), .C(n_592), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_167), .B(n_174), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_166), .B(n_201), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B1(n_171), .B2(n_172), .Y(n_167) );
INVxp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVxp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_175), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g285 ( .A(n_176), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g255 ( .A(n_177), .Y(n_255) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_177), .Y(n_300) );
AND2x2_ASAP7_75t_L g372 ( .A(n_177), .B(n_244), .Y(n_372) );
AND2x4_ASAP7_75t_L g389 ( .A(n_177), .B(n_333), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_177), .B(n_331), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_177), .B(n_240), .Y(n_465) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_185), .A2(n_282), .B1(n_353), .B2(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_212), .Y(n_185) );
INVx2_ASAP7_75t_L g355 ( .A(n_186), .Y(n_355) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_195), .Y(n_186) );
BUFx3_ASAP7_75t_L g345 ( .A(n_187), .Y(n_345) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_188), .B(n_214), .Y(n_237) );
INVx2_ASAP7_75t_L g261 ( .A(n_188), .Y(n_261) );
INVx1_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
AND2x4_ASAP7_75t_L g280 ( .A(n_188), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g297 ( .A(n_188), .B(n_196), .Y(n_297) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_188), .Y(n_311) );
INVxp67_ASAP7_75t_L g319 ( .A(n_188), .Y(n_319) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_194), .Y(n_188) );
INVx2_ASAP7_75t_SL g215 ( .A(n_189), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_189), .A2(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g348 ( .A(n_195), .B(n_264), .Y(n_348) );
AND2x2_ASAP7_75t_L g364 ( .A(n_195), .B(n_265), .Y(n_364) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_195), .B(n_264), .Y(n_451) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x4_ASAP7_75t_L g260 ( .A(n_196), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
INVx1_ASAP7_75t_L g284 ( .A(n_196), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_196), .B(n_226), .Y(n_321) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_205), .Y(n_196) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_204), .A2(n_227), .B(n_233), .Y(n_226) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_204), .A2(n_227), .B(n_233), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g444 ( .A(n_212), .Y(n_444) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_225), .Y(n_212) );
AND2x2_ASAP7_75t_L g318 ( .A(n_213), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g347 ( .A(n_213), .Y(n_347) );
AND2x2_ASAP7_75t_L g449 ( .A(n_213), .B(n_264), .Y(n_449) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_214), .B(n_226), .Y(n_309) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_214) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_265) );
AOI21x1_ASAP7_75t_L g611 ( .A1(n_215), .A2(n_612), .B(n_615), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_217), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g235 ( .A(n_225), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_225), .B(n_345), .Y(n_424) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_226), .Y(n_338) );
AND2x2_ASAP7_75t_L g365 ( .A(n_226), .B(n_311), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g279 ( .A(n_235), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g295 ( .A(n_235), .Y(n_295) );
AND2x2_ASAP7_75t_L g383 ( .A(n_235), .B(n_260), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_235), .B(n_403), .Y(n_408) );
AND2x2_ASAP7_75t_L g418 ( .A(n_235), .B(n_297), .Y(n_418) );
OR2x2_ASAP7_75t_L g455 ( .A(n_235), .B(n_355), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_236), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g415 ( .A(n_236), .B(n_271), .Y(n_415) );
AND2x2_ASAP7_75t_L g431 ( .A(n_236), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g425 ( .A(n_237), .B(n_321), .Y(n_425) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
INVx1_ASAP7_75t_L g307 ( .A(n_239), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_239), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g405 ( .A(n_239), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_239), .B(n_286), .Y(n_430) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_240), .Y(n_277) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_241), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_242), .A2(n_275), .B1(n_293), .B2(n_296), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_242), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g409 ( .A(n_242), .Y(n_409) );
AND2x4_ASAP7_75t_SL g242 ( .A(n_243), .B(n_255), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x4_ASAP7_75t_L g286 ( .A(n_244), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
INVx1_ASAP7_75t_L g333 ( .A(n_244), .Y(n_333) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
NOR3xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .C(n_249), .Y(n_246) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
AND2x4_ASAP7_75t_L g332 ( .A(n_255), .B(n_333), .Y(n_332) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_255), .B(n_362), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
AND2x2_ASAP7_75t_L g357 ( .A(n_257), .B(n_300), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_257), .A2(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_259), .A2(n_369), .B1(n_373), .B2(n_376), .Y(n_368) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_260), .Y(n_326) );
AND2x2_ASAP7_75t_L g336 ( .A(n_260), .B(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g375 ( .A(n_260), .Y(n_375) );
NAND2x1_ASAP7_75t_SL g400 ( .A(n_260), .B(n_269), .Y(n_400) );
AND2x2_ASAP7_75t_L g296 ( .A(n_262), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2x1_ASAP7_75t_L g272 ( .A(n_264), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
INVx2_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
AOI21xp5_ASAP7_75t_SL g266 ( .A1(n_267), .A2(n_274), .B(n_278), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_269), .B(n_463), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_270), .A2(n_359), .B1(n_363), .B2(n_366), .Y(n_358) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
BUFx2_ASAP7_75t_L g463 ( .A(n_271), .Y(n_463) );
INVx1_ASAP7_75t_SL g470 ( .A(n_271), .Y(n_470) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_272), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B(n_285), .Y(n_278) );
AND2x2_ASAP7_75t_L g282 ( .A(n_280), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g324 ( .A(n_280), .B(n_320), .Y(n_324) );
AND2x2_ASAP7_75t_L g439 ( .A(n_280), .B(n_337), .Y(n_439) );
AND2x2_ASAP7_75t_L g442 ( .A(n_280), .B(n_348), .Y(n_442) );
AND2x4_ASAP7_75t_L g450 ( .A(n_280), .B(n_451), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g404 ( .A1(n_282), .A2(n_405), .B(n_407), .Y(n_404) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g432 ( .A(n_284), .Y(n_432) );
AND2x2_ASAP7_75t_L g448 ( .A(n_284), .B(n_449), .Y(n_448) );
INVx4_ASAP7_75t_L g362 ( .A(n_286), .Y(n_362) );
INVx1_ASAP7_75t_L g331 ( .A(n_287), .Y(n_331) );
AND2x2_ASAP7_75t_L g353 ( .A(n_287), .B(n_306), .Y(n_353) );
NOR2x1_ASAP7_75t_L g288 ( .A(n_289), .B(n_312), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .B(n_298), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_291), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_291), .B(n_304), .Y(n_452) );
AND2x2_ASAP7_75t_L g473 ( .A(n_291), .B(n_389), .Y(n_473) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g399 ( .A(n_296), .Y(n_399) );
OAI21xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_301), .B(n_308), .Y(n_298) );
OR2x6_ASAP7_75t_L g351 ( .A(n_300), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_307), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OR2x2_ASAP7_75t_L g374 ( .A(n_309), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g471 ( .A(n_309), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_310), .B(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_325), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_322), .B2(n_324), .Y(n_313) );
OR2x2_ASAP7_75t_L g385 ( .A(n_315), .B(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_317), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g391 ( .A(n_320), .Y(n_391) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_334), .B2(n_336), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AND2x4_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g334 ( .A(n_332), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g395 ( .A(n_335), .B(n_389), .Y(n_395) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_340), .B(n_380), .Y(n_339) );
INVx1_ASAP7_75t_L g523 ( .A(n_340), .Y(n_523) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_341), .B(n_354), .Y(n_340) );
AOI21xp33_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_343), .B(n_349), .Y(n_341) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp33_ASAP7_75t_SL g419 ( .A1(n_351), .A2(n_420), .B1(n_422), .B2(n_425), .Y(n_419) );
NOR2x1_ASAP7_75t_L g366 ( .A(n_352), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g402 ( .A(n_353), .B(n_403), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B(n_358), .C(n_368), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVxp33_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g371 ( .A(n_362), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_363), .A2(n_383), .B1(n_384), .B2(n_387), .C(n_390), .Y(n_382) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g423 ( .A(n_364), .Y(n_423) );
INVx2_ASAP7_75t_SL g421 ( .A(n_367), .Y(n_421) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_371), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g417 ( .A(n_377), .Y(n_417) );
INVx1_ASAP7_75t_L g446 ( .A(n_378), .Y(n_446) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g519 ( .A(n_380), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_380), .A2(n_479), .B(n_521), .Y(n_526) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_396), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_394), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g435 ( .A(n_386), .Y(n_435) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g456 ( .A(n_389), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g461 ( .A(n_389), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVxp33_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g414 ( .A(n_393), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_401), .B(n_404), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
AND2x2_ASAP7_75t_L g445 ( .A(n_406), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_R g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g521 ( .A(n_410), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_426), .C(n_453), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_419), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_416), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_440), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_437), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_436), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_441), .B(n_447), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B(n_452), .Y(n_447) );
INVx1_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B(n_458), .C(n_467), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B1(n_464), .B2(n_466), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g480 ( .A(n_477), .Y(n_480) );
AOI21xp5_ASAP7_75t_SL g524 ( .A1(n_479), .A2(n_522), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g493 ( .A(n_483), .Y(n_493) );
BUFx2_ASAP7_75t_L g509 ( .A(n_483), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
AND2x6_ASAP7_75t_SL g516 ( .A(n_484), .B(n_486), .Y(n_516) );
OR2x6_ASAP7_75t_SL g827 ( .A(n_484), .B(n_485), .Y(n_827) );
OR2x2_ASAP7_75t_L g845 ( .A(n_484), .B(n_486), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g847 ( .A(n_493), .B(n_848), .Y(n_847) );
CKINVDCx9p33_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_SL g497 ( .A(n_498), .B(n_500), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_498), .A2(n_505), .B(n_508), .Y(n_504) );
INVx2_ASAP7_75t_L g850 ( .A(n_498), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g849 ( .A(n_500), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
CKINVDCx11_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx8_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_840), .B(n_846), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_828), .B1(n_835), .B2(n_839), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_517), .B1(n_527), .B2(n_825), .Y(n_512) );
CKINVDCx6p67_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
CKINVDCx11_ASAP7_75t_R g838 ( .A(n_514), .Y(n_838) );
INVx3_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
AOI211xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .B(n_524), .C(n_526), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_518), .A2(n_520), .B(n_524), .Y(n_836) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_526), .B(n_838), .Y(n_837) );
AO22x2_ASAP7_75t_L g835 ( .A1(n_527), .A2(n_826), .B1(n_836), .B2(n_837), .Y(n_835) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_736), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_658), .C(n_708), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_625), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_561), .B1(n_578), .B2(n_608), .C(n_617), .Y(n_531) );
INVx1_ASAP7_75t_SL g707 ( .A(n_532), .Y(n_707) );
AND2x4_ASAP7_75t_SL g532 ( .A(n_533), .B(n_543), .Y(n_532) );
INVx2_ASAP7_75t_L g629 ( .A(n_533), .Y(n_629) );
OR2x2_ASAP7_75t_L g651 ( .A(n_533), .B(n_642), .Y(n_651) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_533), .Y(n_666) );
INVx5_ASAP7_75t_L g673 ( .A(n_533), .Y(n_673) );
AND2x4_ASAP7_75t_L g679 ( .A(n_533), .B(n_553), .Y(n_679) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_533), .B(n_610), .Y(n_682) );
OR2x2_ASAP7_75t_L g691 ( .A(n_533), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g698 ( .A(n_533), .B(n_544), .Y(n_698) );
AND2x2_ASAP7_75t_L g799 ( .A(n_533), .B(n_552), .Y(n_799) );
OR2x6_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx3_ASAP7_75t_SL g650 ( .A(n_543), .Y(n_650) );
AND2x2_ASAP7_75t_L g694 ( .A(n_543), .B(n_610), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_543), .A2(n_698), .B(n_699), .Y(n_697) );
AND2x2_ASAP7_75t_L g735 ( .A(n_543), .B(n_673), .Y(n_735) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_552), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_544), .B(n_553), .Y(n_616) );
OR2x2_ASAP7_75t_L g620 ( .A(n_544), .B(n_553), .Y(n_620) );
INVx1_ASAP7_75t_L g628 ( .A(n_544), .Y(n_628) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_544), .Y(n_640) );
INVx2_ASAP7_75t_L g648 ( .A(n_544), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_544), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g757 ( .A(n_544), .B(n_642), .Y(n_757) );
AND2x2_ASAP7_75t_L g772 ( .A(n_544), .B(n_610), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g641 ( .A(n_553), .B(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_553), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_561), .B(n_765), .Y(n_764) );
NOR2x1p5_ASAP7_75t_L g561 ( .A(n_562), .B(n_569), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g594 ( .A(n_563), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_563), .B(n_570), .Y(n_623) );
INVx1_ASAP7_75t_L g633 ( .A(n_563), .Y(n_633) );
INVx2_ASAP7_75t_L g656 ( .A(n_563), .Y(n_656) );
INVx2_ASAP7_75t_L g662 ( .A(n_563), .Y(n_662) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_563), .Y(n_732) );
OR2x2_ASAP7_75t_L g763 ( .A(n_563), .B(n_570), .Y(n_763) );
OR2x2_ASAP7_75t_L g779 ( .A(n_569), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_570), .B(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g606 ( .A(n_570), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g643 ( .A(n_570), .B(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g655 ( .A(n_570), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g668 ( .A(n_570), .B(n_634), .Y(n_668) );
OR2x2_ASAP7_75t_L g676 ( .A(n_570), .B(n_582), .Y(n_676) );
INVx2_ASAP7_75t_L g703 ( .A(n_570), .Y(n_703) );
INVx1_ASAP7_75t_L g721 ( .A(n_570), .Y(n_721) );
NOR2xp33_ASAP7_75t_R g754 ( .A(n_570), .B(n_595), .Y(n_754) );
OR2x6_ASAP7_75t_L g570 ( .A(n_571), .B(n_577), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_604), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_579), .A2(n_646), .B1(n_649), .B2(n_652), .Y(n_645) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_593), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g660 ( .A(n_581), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g695 ( .A(n_581), .B(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g774 ( .A(n_581), .B(n_752), .Y(n_774) );
INVx3_ASAP7_75t_L g607 ( .A(n_582), .Y(n_607) );
AND2x4_ASAP7_75t_L g634 ( .A(n_582), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_582), .B(n_595), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_582), .B(n_656), .Y(n_701) );
AND2x2_ASAP7_75t_L g706 ( .A(n_582), .B(n_703), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_582), .B(n_594), .Y(n_743) );
INVx1_ASAP7_75t_L g813 ( .A(n_582), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_582), .B(n_731), .Y(n_824) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_588), .Y(n_582) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g605 ( .A(n_595), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_595), .B(n_607), .Y(n_624) );
INVx2_ASAP7_75t_L g635 ( .A(n_595), .Y(n_635) );
AND2x2_ASAP7_75t_L g661 ( .A(n_595), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g677 ( .A(n_595), .B(n_656), .Y(n_677) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_595), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_595), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g766 ( .A(n_595), .Y(n_766) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_605), .B(n_633), .Y(n_644) );
AOI221x1_ASAP7_75t_SL g738 ( .A1(n_606), .A2(n_739), .B1(n_742), .B2(n_744), .C(n_748), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_606), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g796 ( .A(n_606), .B(n_661), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_606), .B(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g727 ( .A(n_607), .B(n_655), .Y(n_727) );
AND2x2_ASAP7_75t_L g765 ( .A(n_607), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_616), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_610), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g713 ( .A(n_610), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_610), .B(n_629), .Y(n_718) );
AND2x4_ASAP7_75t_L g747 ( .A(n_610), .B(n_648), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_610), .B(n_679), .Y(n_783) );
OR2x2_ASAP7_75t_L g801 ( .A(n_610), .B(n_732), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_610), .B(n_692), .Y(n_811) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g642 ( .A(n_611), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g667 ( .A(n_616), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_616), .A2(n_675), .B1(n_678), .B2(n_680), .Y(n_674) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
INVx2_ASAP7_75t_L g630 ( .A(n_618), .Y(n_630) );
AND2x2_ASAP7_75t_L g769 ( .A(n_619), .B(n_629), .Y(n_769) );
AND2x2_ASAP7_75t_L g815 ( .A(n_619), .B(n_682), .Y(n_815) );
AND2x2_ASAP7_75t_L g820 ( .A(n_619), .B(n_671), .Y(n_820) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI32xp33_ASAP7_75t_L g789 ( .A1(n_621), .A2(n_691), .A3(n_771), .B1(n_790), .B2(n_792), .Y(n_789) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g657 ( .A(n_624), .Y(n_657) );
AOI211xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_631), .B(n_636), .C(n_645), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_628), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_629), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g809 ( .A(n_629), .Y(n_809) );
AND2x2_ASAP7_75t_L g719 ( .A(n_631), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_632), .B(n_634), .Y(n_631) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_632), .Y(n_819) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_633), .Y(n_688) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_633), .Y(n_788) );
INVx1_ASAP7_75t_L g685 ( .A(n_634), .Y(n_685) );
AND2x2_ASAP7_75t_L g751 ( .A(n_634), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_634), .B(n_762), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_643), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g717 ( .A1(n_638), .A2(n_718), .B(n_719), .Y(n_717) );
AND2x2_ASAP7_75t_SL g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g647 ( .A(n_642), .B(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g671 ( .A(n_642), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_647), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g778 ( .A(n_647), .Y(n_778) );
AND2x2_ASAP7_75t_L g808 ( .A(n_647), .B(n_809), .Y(n_808) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_648), .Y(n_785) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_650), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_SL g725 ( .A(n_651), .Y(n_725) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g684 ( .A(n_655), .B(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_656), .Y(n_752) );
AND2x2_ASAP7_75t_L g761 ( .A(n_657), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_681), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_668), .B2(n_669), .C(n_674), .Y(n_659) );
INVx1_ASAP7_75t_L g780 ( .A(n_661), .Y(n_780) );
INVxp33_ASAP7_75t_SL g812 ( .A(n_661), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_663), .A2(n_759), .B(n_767), .Y(n_758) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_667), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g680 ( .A(n_668), .Y(n_680) );
AND2x2_ASAP7_75t_L g715 ( .A(n_668), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g734 ( .A(n_668), .B(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_668), .A2(n_796), .B1(n_797), .B2(n_800), .Y(n_795) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OR2x2_ASAP7_75t_L g690 ( .A(n_671), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_671), .B(n_679), .Y(n_729) );
AND2x4_ASAP7_75t_L g746 ( .A(n_673), .B(n_692), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_673), .B(n_747), .Y(n_793) );
AND2x2_ASAP7_75t_L g805 ( .A(n_673), .B(n_757), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g790 ( .A(n_675), .B(n_791), .Y(n_790) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_SL g733 ( .A(n_676), .Y(n_733) );
INVx1_ASAP7_75t_L g804 ( .A(n_677), .Y(n_804) );
INVx2_ASAP7_75t_SL g756 ( .A(n_679), .Y(n_756) );
AOI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B(n_686), .C(n_704), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .B(n_693), .C(n_697), .Y(n_686) );
OR2x6_ASAP7_75t_SL g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g716 ( .A(n_688), .Y(n_716) );
INVx1_ASAP7_75t_SL g741 ( .A(n_691), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_691), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_696), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_700), .A2(n_783), .B1(n_784), .B2(n_786), .Y(n_782) );
OR2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_714), .B(n_717), .C(n_722), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_726), .B1(n_728), .B2(n_730), .C(n_734), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI222xp33_ASAP7_75t_L g814 ( .A1(n_733), .A2(n_815), .B1(n_816), .B2(n_820), .C1(n_821), .C2(n_823), .Y(n_814) );
INVx2_ASAP7_75t_L g749 ( .A(n_735), .Y(n_749) );
NOR3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_775), .C(n_794), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_758), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_746), .B(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_747), .B(n_809), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_753), .B2(n_755), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVxp33_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_756), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_764), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_764), .A2(n_768), .B1(n_770), .B2(n_773), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
CKINVDCx16_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
OAI211xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_779), .B(n_781), .C(n_789), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_802), .C(n_814), .Y(n_794) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_806), .B(n_813), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_810), .B(n_812), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
CKINVDCx11_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g839 ( .A(n_828), .Y(n_839) );
INVxp33_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVxp33_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
INVx1_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_SL g846 ( .A(n_847), .Y(n_846) );
INVxp67_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
endmodule