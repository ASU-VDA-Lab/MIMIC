module fake_jpeg_19169_n_164 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_30),
.B(n_24),
.C(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_17),
.B1(n_27),
.B2(n_16),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_27),
.B1(n_16),
.B2(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_59),
.B1(n_56),
.B2(n_45),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_60),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_15),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_31),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_39),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_37),
.C(n_36),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_64),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_57),
.C(n_53),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_39),
.B1(n_37),
.B2(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_28),
.B1(n_21),
.B2(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_74),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_48),
.B(n_44),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_92),
.B(n_98),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_44),
.B(n_45),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_47),
.B(n_4),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_47),
.B(n_3),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_67),
.B1(n_64),
.B2(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_69),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_12),
.Y(n_122)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_73),
.B1(n_85),
.B2(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_123),
.B1(n_89),
.B2(n_99),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_79),
.B1(n_78),
.B2(n_75),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_113),
.B(n_100),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_81),
.B1(n_74),
.B2(n_70),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_6),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_11),
.C(n_12),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_99),
.C(n_106),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_13),
.B1(n_109),
.B2(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_112),
.B(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_108),
.B1(n_103),
.B2(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_114),
.B1(n_117),
.B2(n_93),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_105),
.C(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_128),
.C(n_133),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_102),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_140),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_139),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_117),
.B1(n_93),
.B2(n_102),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_98),
.B1(n_104),
.B2(n_95),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_130),
.C(n_132),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_138),
.C(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_149),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_107),
.C(n_142),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_155),
.Y(n_159)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_144),
.B(n_139),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_150),
.B(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.C(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_153),
.C(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);


endmodule