module fake_jpeg_31256_n_550 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_550);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_29),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_72),
.B(n_98),
.Y(n_146)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_33),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_100),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_102),
.Y(n_169)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_106),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_24),
.A2(n_16),
.B(n_14),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_54),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_18),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_111),
.Y(n_141)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_109),
.Y(n_144)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_50),
.Y(n_151)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_34),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_33),
.B1(n_22),
.B2(n_51),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_115),
.A2(n_136),
.B1(n_160),
.B2(n_179),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_49),
.B1(n_26),
.B2(n_18),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_119),
.B(n_121),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_44),
.B(n_52),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_132),
.B(n_149),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_71),
.A2(n_33),
.B1(n_50),
.B2(n_51),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_134),
.A2(n_113),
.B1(n_111),
.B2(n_85),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_49),
.B1(n_26),
.B2(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_139),
.B(n_157),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_69),
.B(n_32),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_151),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_69),
.B(n_44),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_52),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_174),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_88),
.A2(n_27),
.B1(n_48),
.B2(n_45),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_75),
.B(n_27),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_176),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_89),
.A2(n_30),
.B1(n_39),
.B2(n_54),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_168),
.A2(n_134),
.B1(n_131),
.B2(n_161),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_105),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_90),
.B(n_48),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_96),
.B(n_43),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_97),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_186),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_117),
.A2(n_101),
.B1(n_57),
.B2(n_58),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_182),
.A2(n_184),
.B1(n_187),
.B2(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_124),
.A2(n_62),
.B1(n_68),
.B2(n_70),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_39),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_122),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_188),
.B(n_191),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_42),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_208),
.Y(n_246)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_135),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_202),
.Y(n_257)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_196),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_123),
.B1(n_164),
.B2(n_154),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_83),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_201),
.A2(n_226),
.B(n_231),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_130),
.A2(n_38),
.B(n_64),
.C(n_78),
.D(n_77),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_205),
.B(n_209),
.Y(n_264)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_206),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_131),
.A2(n_38),
.B1(n_82),
.B2(n_80),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_207),
.A2(n_172),
.B1(n_171),
.B2(n_148),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_146),
.B(n_0),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_0),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_163),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_210),
.Y(n_280)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_213),
.Y(n_270)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_142),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_218),
.Y(n_271)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_222),
.Y(n_261)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_115),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_140),
.B1(n_143),
.B2(n_178),
.Y(n_259)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_142),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_236),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_116),
.B(n_2),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_233),
.Y(n_238)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_3),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_165),
.B(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_153),
.B(n_4),
.Y(n_237)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx6_ASAP7_75t_SL g250 ( 
.A(n_210),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_222),
.A2(n_163),
.B1(n_133),
.B2(n_116),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_212),
.B1(n_195),
.B2(n_214),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_266),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_204),
.A2(n_178),
.B1(n_172),
.B2(n_171),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_181),
.B1(n_219),
.B2(n_203),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_259),
.A2(n_281),
.B1(n_215),
.B2(n_228),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_211),
.B(n_175),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_232),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_273),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_288),
.B1(n_301),
.B2(n_239),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_186),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_306),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_256),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_194),
.B(n_201),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_291),
.A2(n_304),
.B(n_248),
.Y(n_325)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_241),
.B(n_208),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_293),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_194),
.C(n_181),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_317),
.C(n_238),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_302),
.Y(n_323)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_259),
.A2(n_204),
.B1(n_200),
.B2(n_184),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_201),
.B(n_231),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_266),
.B1(n_190),
.B2(n_242),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_189),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_246),
.B(n_227),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_237),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_311),
.Y(n_340)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_264),
.A2(n_226),
.B(n_231),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_312),
.A2(n_315),
.B(n_316),
.Y(n_346)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_283),
.Y(n_328)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_205),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_257),
.B(n_235),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_198),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_318),
.A2(n_335),
.B1(n_341),
.B2(n_305),
.Y(n_358)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_275),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_336),
.C(n_339),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_326),
.A2(n_337),
.B1(n_314),
.B2(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_300),
.A2(n_250),
.B1(n_274),
.B2(n_242),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_329),
.A2(n_280),
.B1(n_274),
.B2(n_289),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_254),
.B1(n_229),
.B2(n_220),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_249),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_292),
.A2(n_234),
.B1(n_233),
.B2(n_213),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_288),
.A2(n_296),
.B1(n_315),
.B2(n_316),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_345),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_249),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_317),
.C(n_304),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_243),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_298),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_316),
.Y(n_351)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_350),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_291),
.C(n_293),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_354),
.B(n_361),
.C(n_366),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_299),
.Y(n_355)
);

AO21x1_ASAP7_75t_L g408 ( 
.A1(n_355),
.A2(n_377),
.B(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_358),
.A2(n_378),
.B1(n_333),
.B2(n_327),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_299),
.Y(n_360)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_293),
.C(n_309),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_310),
.Y(n_362)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_332),
.B(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_365),
.Y(n_383)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_364),
.Y(n_398)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_312),
.C(n_311),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_368),
.Y(n_396)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_344),
.B1(n_324),
.B2(n_319),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_345),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_370),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_371),
.A2(n_320),
.B1(n_338),
.B2(n_319),
.Y(n_381)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_374),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_331),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_373),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_332),
.B(n_308),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_341),
.B(n_303),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_325),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_297),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_265),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_290),
.B(n_284),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_318),
.A2(n_285),
.B1(n_287),
.B2(n_302),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_352),
.A2(n_333),
.B(n_338),
.C(n_343),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_380),
.A2(n_399),
.B(n_349),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_381),
.A2(n_245),
.B1(n_280),
.B2(n_240),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_382),
.A2(n_384),
.B1(n_388),
.B2(n_245),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_327),
.B1(n_336),
.B2(n_335),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_355),
.A2(n_337),
.B1(n_346),
.B2(n_343),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_397),
.B1(n_255),
.B2(n_217),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_353),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_392),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_404),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_366),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_393),
.B(n_368),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_364),
.A2(n_334),
.B1(n_344),
.B2(n_324),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_252),
.B(n_244),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_351),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_365),
.C(n_376),
.Y(n_411)
);

AOI21xp33_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_243),
.B(n_269),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_SL g438 ( 
.A(n_401),
.B(n_277),
.C(n_272),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_377),
.A2(n_244),
.B(n_247),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_405),
.A2(n_371),
.B(n_372),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_356),
.B(n_269),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_406),
.B(n_247),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_248),
.Y(n_407)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_378),
.B(n_369),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_412),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_414),
.C(n_427),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_394),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_396),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_413),
.B(n_424),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_355),
.C(n_367),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_416),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_417),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_370),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_423),
.Y(n_460)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_420),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_421),
.A2(n_199),
.B(n_129),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_422),
.B(n_384),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_402),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_359),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_430),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_359),
.B(n_349),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_277),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_390),
.C(n_392),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_428),
.A2(n_438),
.B1(n_381),
.B2(n_405),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_432),
.A2(n_263),
.B1(n_267),
.B2(n_206),
.Y(n_456)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_402),
.Y(n_433)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_434),
.B(n_437),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_436),
.A2(n_398),
.B1(n_395),
.B2(n_397),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_388),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_439),
.A2(n_444),
.B1(n_454),
.B2(n_438),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_409),
.C(n_400),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_448),
.C(n_452),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_453),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_382),
.B1(n_395),
.B2(n_399),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_445),
.A2(n_456),
.B1(n_459),
.B2(n_434),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_407),
.C(n_408),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_380),
.C(n_255),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_436),
.A2(n_272),
.B1(n_263),
.B2(n_267),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_145),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_458),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_415),
.A2(n_225),
.B1(n_148),
.B2(n_129),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_422),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_474),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_420),
.C(n_419),
.Y(n_464)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_457),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_472),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_475),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_411),
.C(n_424),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_470),
.B(n_476),
.C(n_447),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_457),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_473),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_419),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_417),
.C(n_433),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_429),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_478),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_416),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_421),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_458),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_431),
.Y(n_480)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

NOR2x1_ASAP7_75t_R g481 ( 
.A(n_457),
.B(n_413),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_481),
.A2(n_461),
.B(n_440),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_453),
.C(n_450),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_483),
.C(n_493),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_439),
.C(n_444),
.Y(n_483)
);

AO21x1_ASAP7_75t_L g510 ( 
.A1(n_484),
.A2(n_145),
.B(n_9),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_494),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_481),
.Y(n_492)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_492),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_447),
.C(n_449),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_454),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_466),
.Y(n_497)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_497),
.Y(n_509)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_498),
.A2(n_469),
.B1(n_5),
.B2(n_7),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_499),
.B(n_478),
.C(n_479),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_502),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_485),
.A2(n_451),
.B1(n_463),
.B2(n_459),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_469),
.C(n_456),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_504),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_128),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_507),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_487),
.A2(n_170),
.B1(n_7),
.B2(n_8),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_513),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_9),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_145),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_511),
.Y(n_516)
);

NOR2x1p5_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_4),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_512),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_9),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_491),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_487),
.Y(n_521)
);

FAx1_ASAP7_75t_SL g517 ( 
.A(n_514),
.B(n_489),
.CI(n_488),
.CON(n_517),
.SN(n_517)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_488),
.C(n_494),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_520),
.B(n_522),
.Y(n_529)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_521),
.Y(n_534)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_9),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_525),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_515),
.B1(n_506),
.B2(n_509),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_528),
.A2(n_533),
.B1(n_519),
.B2(n_517),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_511),
.C(n_508),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_530),
.B(n_535),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_522),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_520),
.Y(n_535)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_529),
.A2(n_510),
.B(n_516),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_536),
.B(n_537),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_531),
.A2(n_517),
.B(n_527),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_538),
.B(n_539),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_533),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_534),
.C(n_532),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_543),
.A2(n_525),
.B(n_10),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_544),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_541),
.B(n_10),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_545),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_542),
.B(n_10),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_11),
.C(n_403),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_11),
.Y(n_550)
);


endmodule