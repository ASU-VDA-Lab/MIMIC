module fake_jpeg_18879_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_50),
.B1(n_55),
.B2(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_52),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_18),
.B2(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_22),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_33),
.B1(n_21),
.B2(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_42),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_41),
.C(n_39),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_63),
.C(n_35),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_84),
.B1(n_35),
.B2(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_41),
.C(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_38),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_73),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_70),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_38),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_80),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_17),
.B(n_25),
.C(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_21),
.B1(n_39),
.B2(n_34),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_86),
.B1(n_40),
.B2(n_53),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_17),
.B(n_29),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_42),
.B1(n_40),
.B2(n_33),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_42),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_44),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_16),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_21),
.B1(n_40),
.B2(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_76),
.B1(n_74),
.B2(n_62),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_49),
.B(n_25),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_85),
.B(n_68),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_108),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_40),
.B1(n_28),
.B2(n_32),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_32),
.B1(n_31),
.B2(n_28),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_99),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_31),
.B1(n_44),
.B2(n_29),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_35),
.B1(n_24),
.B2(n_22),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_35),
.B1(n_72),
.B2(n_22),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_71),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_113),
.B(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_67),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_0),
.B(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_125),
.B1(n_58),
.B2(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_26),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_73),
.B(n_85),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_130),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_15),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_91),
.B1(n_106),
.B2(n_101),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_109),
.B1(n_90),
.B2(n_103),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_111),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_140),
.B1(n_142),
.B2(n_146),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_91),
.B(n_103),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_144),
.B(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_91),
.B1(n_104),
.B2(n_98),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_108),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_105),
.B1(n_107),
.B2(n_30),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_118),
.B(n_127),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_105),
.B1(n_107),
.B2(n_30),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_117),
.B1(n_128),
.B2(n_5),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_135),
.B1(n_125),
.B2(n_130),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_58),
.B(n_1),
.Y(n_150)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_126),
.A3(n_122),
.B1(n_131),
.B2(n_120),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_117),
.Y(n_161)
);

AO22x1_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_58),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_3),
.B(n_4),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_140),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_149),
.B1(n_147),
.B2(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_14),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_166),
.A2(n_174),
.B(n_163),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_4),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_5),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_152),
.C(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_136),
.C(n_150),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_177),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_191),
.B1(n_153),
.B2(n_190),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_189),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_172),
.B(n_176),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_139),
.C(n_146),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_195),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_172),
.B1(n_177),
.B2(n_162),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_165),
.B(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_162),
.B1(n_153),
.B2(n_158),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_161),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_178),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_192),
.B(n_189),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_174),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_174),
.C(n_148),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_174),
.B(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_193),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_185),
.C(n_180),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_196),
.C(n_194),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_209),
.C(n_9),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_197),
.C(n_147),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_11),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_8),
.B(n_10),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_8),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_10),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_11),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.C(n_215),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.C(n_225),
.Y(n_229)
);

AOI21x1_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_216),
.B(n_12),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_11),
.B(n_13),
.C(n_186),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_13),
.Y(n_232)
);


endmodule