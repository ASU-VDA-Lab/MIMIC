module fake_ibex_175_n_3554 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_898, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_3554);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_3554;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_2017;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_2290;
wire n_957;
wire n_3272;
wire n_3255;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_2918;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_2957;
wire n_2586;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_978;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3510;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_2369;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_1395;
wire n_998;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_1400;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_3495;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1683;
wire n_1185;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_2180;
wire n_1952;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3427;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_3162;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_2272;
wire n_1956;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2675;
wire n_2417;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_956;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_2119;
wire n_1010;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_1762;
wire n_940;
wire n_2534;
wire n_1404;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_2544;
wire n_3193;
wire n_3501;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_SL g907 ( 
.A(n_361),
.Y(n_907)
);

CKINVDCx16_ASAP7_75t_R g908 ( 
.A(n_276),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_539),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_297),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_634),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_106),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_48),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_866),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_290),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_341),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_105),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_20),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_581),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_664),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_675),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_610),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_814),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_246),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_554),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_328),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_287),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_272),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_330),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_166),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_697),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_771),
.Y(n_932)
);

CKINVDCx14_ASAP7_75t_R g933 ( 
.A(n_254),
.Y(n_933)
);

INVxp33_ASAP7_75t_L g934 ( 
.A(n_127),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_551),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_754),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_654),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_633),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_877),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_52),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_122),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_320),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_272),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_75),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_545),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_208),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_867),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_735),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_593),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_500),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_39),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_773),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_437),
.Y(n_953)
);

CKINVDCx16_ASAP7_75t_R g954 ( 
.A(n_324),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_873),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_724),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_371),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_627),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_557),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_485),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_819),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_884),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_218),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_906),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_634),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_338),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_359),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_315),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_757),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_292),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_568),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_11),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_583),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_53),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_758),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_243),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_78),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_821),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_745),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_460),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_258),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_787),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_868),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_489),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_617),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_500),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_850),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_875),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_375),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_63),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_609),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_708),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_879),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_482),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_587),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_91),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_636),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_628),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_905),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_649),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_279),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_462),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_854),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_359),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_846),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_173),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_771),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_490),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_485),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_109),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_593),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_696),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_613),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_6),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_18),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_58),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_350),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_217),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_855),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_876),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_800),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_645),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_570),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_785),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_528),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_587),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_824),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_675),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_706),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_878),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_870),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_68),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_758),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_863),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_717),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_799),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_376),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_25),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_116),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_79),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_29),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_189),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_132),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_269),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_616),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_534),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_48),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_595),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_282),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_376),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_65),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_403),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_357),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_838),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_274),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_204),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_196),
.Y(n_1057)
);

BUFx5_ASAP7_75t_L g1058 ( 
.A(n_391),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_621),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_184),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_457),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_398),
.Y(n_1062)
);

BUFx10_ASAP7_75t_L g1063 ( 
.A(n_826),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_762),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_872),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_741),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_128),
.Y(n_1067)
);

INVxp33_ASAP7_75t_L g1068 ( 
.A(n_525),
.Y(n_1068)
);

BUFx5_ASAP7_75t_L g1069 ( 
.A(n_575),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_400),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_326),
.Y(n_1071)
);

INVx4_ASAP7_75t_R g1072 ( 
.A(n_852),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_793),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_871),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_630),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_904),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_415),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_740),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_433),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_849),
.Y(n_1080)
);

CKINVDCx14_ASAP7_75t_R g1081 ( 
.A(n_148),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_431),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_700),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_559),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_859),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_491),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_470),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_559),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_811),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_897),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_265),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_716),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_614),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_444),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_863),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_722),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_769),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_455),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_551),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_176),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_635),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_232),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_837),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_62),
.Y(n_1104)
);

BUFx5_ASAP7_75t_L g1105 ( 
.A(n_727),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_66),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_436),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_646),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_300),
.Y(n_1109)
);

BUFx10_ASAP7_75t_L g1110 ( 
.A(n_237),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_531),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_425),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_361),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_718),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_619),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_587),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_106),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_568),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_393),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_127),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_683),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_861),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_865),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_141),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_25),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_809),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_848),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_56),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_407),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_246),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_851),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_860),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_853),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_768),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_81),
.Y(n_1135)
);

BUFx10_ASAP7_75t_L g1136 ( 
.A(n_838),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_869),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_67),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_880),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_340),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_537),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_849),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_238),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_456),
.Y(n_1144)
);

CKINVDCx16_ASAP7_75t_R g1145 ( 
.A(n_790),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_45),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_3),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_762),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_417),
.Y(n_1149)
);

BUFx5_ASAP7_75t_L g1150 ( 
.A(n_510),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_584),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_26),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_319),
.Y(n_1153)
);

BUFx5_ASAP7_75t_L g1154 ( 
.A(n_185),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_444),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_200),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_199),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_572),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_737),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_726),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_520),
.Y(n_1161)
);

BUFx10_ASAP7_75t_L g1162 ( 
.A(n_230),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_864),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_503),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_884),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_397),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_722),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_206),
.Y(n_1168)
);

BUFx8_ASAP7_75t_SL g1169 ( 
.A(n_549),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_229),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_861),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_724),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_903),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_473),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_103),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_698),
.Y(n_1176)
);

BUFx10_ASAP7_75t_L g1177 ( 
.A(n_74),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_17),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_406),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_339),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_830),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_729),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_762),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_385),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_711),
.Y(n_1185)
);

CKINVDCx14_ASAP7_75t_R g1186 ( 
.A(n_182),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_24),
.Y(n_1187)
);

BUFx5_ASAP7_75t_L g1188 ( 
.A(n_32),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_741),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_794),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_700),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_269),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_248),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_468),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_403),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_331),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_483),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_874),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_845),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_856),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_857),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_122),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_47),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_858),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_150),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_72),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_86),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_132),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_406),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_280),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_260),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_593),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_676),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_494),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_10),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_672),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_278),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_6),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_696),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_120),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_442),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_727),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_575),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_828),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_49),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_16),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_592),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_738),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_747),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_597),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_761),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_237),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_488),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_557),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_240),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_882),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_129),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_86),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_115),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_134),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_896),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_186),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_413),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_728),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_166),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_881),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_148),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_506),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_370),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_414),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_600),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_644),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_327),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_268),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_237),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_332),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_847),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_528),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_862),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_759),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_625),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_855),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_232),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_329),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_902),
.Y(n_1265)
);

BUFx10_ASAP7_75t_L g1266 ( 
.A(n_864),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_561),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_73),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_545),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_54),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_309),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_776),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_376),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_2),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_428),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_3),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_344),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_883),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_448),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1177),
.Y(n_1280)
);

INVxp33_ASAP7_75t_SL g1281 ( 
.A(n_957),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1225),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1177),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1177),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_972),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1047),
.Y(n_1286)
);

INVxp33_ASAP7_75t_SL g1287 ( 
.A(n_1012),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1215),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1225),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1188),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1225),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_974),
.Y(n_1292)
);

INVxp33_ASAP7_75t_SL g1293 ( 
.A(n_1017),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1106),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_977),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1014),
.Y(n_1296)
);

INVxp67_ASAP7_75t_SL g1297 ( 
.A(n_1106),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1038),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_933),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1081),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_981),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1188),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1040),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1125),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1146),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_973),
.Y(n_1306)
);

INVxp33_ASAP7_75t_L g1307 ( 
.A(n_1133),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1015),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1276),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1186),
.Y(n_1310)
);

INVxp33_ASAP7_75t_SL g1311 ( 
.A(n_1277),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_981),
.Y(n_1312)
);

INVxp67_ASAP7_75t_SL g1313 ( 
.A(n_934),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1088),
.Y(n_1314)
);

INVxp33_ASAP7_75t_SL g1315 ( 
.A(n_913),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1169),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1173),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1199),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1249),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1258),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_965),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_917),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1023),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1191),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1188),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1195),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1169),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1228),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1241),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1188),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_908),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1058),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_990),
.Y(n_1333)
);

INVxp33_ASAP7_75t_SL g1334 ( 
.A(n_940),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_922),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_944),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_951),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1068),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_990),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_923),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_925),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1058),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1058),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1016),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1058),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1041),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1051),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_960),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1058),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_921),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_961),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_962),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_967),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_969),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1058),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_970),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_971),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1068),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1104),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_975),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_976),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_920),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_980),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_982),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1058),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_983),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1135),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1032),
.Y(n_1368)
);

INVxp33_ASAP7_75t_SL g1369 ( 
.A(n_1128),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_918),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1138),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_973),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_987),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_918),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_964),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_991),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_921),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1282),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1307),
.B(n_954),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1368),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1306),
.Y(n_1381)
);

OAI22x1_ASAP7_75t_L g1382 ( 
.A1(n_1368),
.A2(n_1152),
.B1(n_1178),
.B2(n_1147),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1306),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1300),
.B(n_943),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1306),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1372),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1289),
.A2(n_1226),
.B(n_911),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1288),
.A2(n_1203),
.B1(n_1206),
.B2(n_1187),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1291),
.A2(n_1226),
.B(n_911),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1292),
.A2(n_1296),
.B(n_1295),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1338),
.B(n_1207),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1315),
.B(n_1145),
.Y(n_1392)
);

AND2x6_ASAP7_75t_L g1393 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1358),
.A2(n_1238),
.B1(n_1270),
.B2(n_1218),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1308),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1370),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1372),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1370),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1298),
.Y(n_1399)
);

INVx6_ASAP7_75t_L g1400 ( 
.A(n_1331),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1290),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1294),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1297),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1303),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1333),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1304),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1301),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1305),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1329),
.B(n_1321),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1284),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1334),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1332),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1302),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1312),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1367),
.B(n_917),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1369),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1342),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1343),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1345),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1330),
.A2(n_937),
.B(n_910),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1325),
.A2(n_937),
.B(n_910),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1350),
.B(n_912),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1336),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1337),
.B(n_1344),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1349),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1377),
.B(n_914),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1323),
.B(n_943),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1355),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1374),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1339),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1346),
.Y(n_1431)
);

INVx5_ASAP7_75t_L g1432 ( 
.A(n_1365),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1309),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1347),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1314),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1359),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1317),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1318),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1319),
.Y(n_1439)
);

AND2x6_ASAP7_75t_L g1440 ( 
.A(n_1285),
.B(n_966),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1286),
.B(n_966),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1320),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1287),
.A2(n_1002),
.B1(n_1004),
.B2(n_997),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1293),
.A2(n_1004),
.B1(n_1005),
.B2(n_1002),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1371),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1335),
.Y(n_1446)
);

INVx5_ASAP7_75t_L g1447 ( 
.A(n_1311),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1340),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1341),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1376),
.A2(n_992),
.B(n_986),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1324),
.B(n_968),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1348),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1351),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1352),
.Y(n_1455)
);

AND2x6_ASAP7_75t_L g1456 ( 
.A(n_1326),
.B(n_984),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1353),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1354),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1356),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1299),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1328),
.B(n_917),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1357),
.Y(n_1462)
);

AND2x6_ASAP7_75t_L g1463 ( 
.A(n_1360),
.B(n_984),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1375),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1310),
.B(n_927),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1361),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1363),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1364),
.B(n_927),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1366),
.B(n_927),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1373),
.B(n_1037),
.Y(n_1470)
);

BUFx8_ASAP7_75t_L g1471 ( 
.A(n_1362),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1282),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1288),
.A2(n_916),
.B1(n_919),
.B2(n_915),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1307),
.B(n_952),
.Y(n_1474)
);

BUFx8_ASAP7_75t_L g1475 ( 
.A(n_1300),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1282),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1282),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1282),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1282),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1282),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1282),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1282),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1313),
.B(n_924),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1282),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1282),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1313),
.B(n_926),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1282),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1288),
.A2(n_929),
.B1(n_931),
.B2(n_928),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1313),
.B(n_935),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1282),
.Y(n_1490)
);

BUFx8_ASAP7_75t_L g1491 ( 
.A(n_1300),
.Y(n_1491)
);

OAI22x1_ASAP7_75t_L g1492 ( 
.A1(n_1368),
.A2(n_938),
.B1(n_939),
.B2(n_936),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1315),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1282),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1289),
.A2(n_1000),
.B(n_994),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1281),
.A2(n_1060),
.B1(n_1094),
.B2(n_1056),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1313),
.B(n_952),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1282),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1307),
.B(n_952),
.Y(n_1499)
);

INVx5_ASAP7_75t_L g1500 ( 
.A(n_1322),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1289),
.A2(n_1001),
.B(n_1000),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1282),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1313),
.B(n_941),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1313),
.B(n_942),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1282),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1288),
.A2(n_946),
.B1(n_947),
.B2(n_945),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1368),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1313),
.B(n_948),
.Y(n_1508)
);

BUFx12f_ASAP7_75t_L g1509 ( 
.A(n_1316),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1368),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1282),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

BUFx8_ASAP7_75t_L g1513 ( 
.A(n_1300),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1282),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1281),
.A2(n_1117),
.B1(n_1132),
.B2(n_1100),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1368),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1390),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1396),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1501),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1387),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1389),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1398),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1450),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1510),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1405),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1437),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_R g1527 ( 
.A(n_1416),
.B(n_1140),
.Y(n_1527)
);

BUFx10_ASAP7_75t_L g1528 ( 
.A(n_1507),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1395),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1493),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_R g1531 ( 
.A(n_1452),
.B(n_1140),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1430),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1495),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1471),
.Y(n_1534)
);

BUFx10_ASAP7_75t_L g1535 ( 
.A(n_1507),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1464),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1434),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1442),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1461),
.B(n_999),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1421),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1509),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_R g1542 ( 
.A(n_1400),
.B(n_1143),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1429),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1420),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1475),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1379),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1447),
.B(n_0),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1491),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1513),
.Y(n_1549)
);

XNOR2xp5_ASAP7_75t_L g1550 ( 
.A(n_1443),
.B(n_1149),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_L g1551 ( 
.A(n_1447),
.B(n_0),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1404),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1404),
.Y(n_1553)
);

BUFx10_ASAP7_75t_L g1554 ( 
.A(n_1409),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_R g1555 ( 
.A(n_1423),
.B(n_1149),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1458),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1444),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1496),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1435),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1515),
.Y(n_1560)
);

NAND2xp33_ASAP7_75t_SL g1561 ( 
.A(n_1445),
.B(n_950),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1406),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1474),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1388),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1431),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1473),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1488),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1499),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1439),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1506),
.Y(n_1570)
);

AND3x2_ASAP7_75t_L g1571 ( 
.A(n_1436),
.B(n_1192),
.C(n_1176),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1399),
.B(n_1069),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1394),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1382),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1497),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1454),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1454),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1433),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1422),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1433),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1492),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1468),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1460),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1456),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1463),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1415),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_R g1587 ( 
.A(n_1440),
.B(n_1192),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1457),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1463),
.Y(n_1589)
);

INVx11_ASAP7_75t_L g1590 ( 
.A(n_1456),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1469),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1456),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1500),
.B(n_0),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1463),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1424),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1426),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1477),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_R g1598 ( 
.A(n_1465),
.B(n_953),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1408),
.B(n_956),
.Y(n_1599)
);

NOR2xp67_ASAP7_75t_L g1600 ( 
.A(n_1500),
.B(n_0),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1408),
.B(n_956),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_R g1602 ( 
.A(n_1410),
.B(n_1193),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1466),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1407),
.A2(n_1246),
.B1(n_1257),
.B2(n_1244),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1384),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1392),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1391),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1449),
.B(n_956),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1378),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1378),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1438),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1472),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1476),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1479),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1480),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1414),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1483),
.B(n_955),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1481),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1478),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1403),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1481),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1486),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_R g1623 ( 
.A(n_1410),
.B(n_1244),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1489),
.B(n_958),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1484),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1490),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1503),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1504),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1508),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1494),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1505),
.Y(n_1631)
);

BUFx3_ASAP7_75t_SL g1632 ( 
.A(n_1393),
.Y(n_1632)
);

NAND2xp33_ASAP7_75t_R g1633 ( 
.A(n_1427),
.B(n_959),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1498),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1393),
.Y(n_1635)
);

BUFx10_ASAP7_75t_L g1636 ( 
.A(n_1470),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1451),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1502),
.Y(n_1638)
);

BUFx10_ASAP7_75t_L g1639 ( 
.A(n_1402),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1511),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1446),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1448),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1482),
.Y(n_1643)
);

BUFx10_ASAP7_75t_L g1644 ( 
.A(n_1485),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1487),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1453),
.B(n_1069),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1455),
.B(n_1069),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1459),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1462),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1514),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_SL g1651 ( 
.A(n_1467),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1432),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1412),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1441),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1417),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1425),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1418),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1428),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1418),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1401),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1419),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1413),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1381),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1397),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1383),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1383),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1385),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1385),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1386),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1386),
.A2(n_1009),
.B(n_1001),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1380),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1380),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1390),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1380),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1501),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1380),
.B(n_907),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1380),
.Y(n_1677)
);

NAND2xp33_ASAP7_75t_R g1678 ( 
.A(n_1411),
.B(n_963),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1501),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1512),
.B(n_1),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1380),
.Y(n_1681)
);

INVxp33_ASAP7_75t_L g1682 ( 
.A(n_1516),
.Y(n_1682)
);

BUFx10_ASAP7_75t_L g1683 ( 
.A(n_1516),
.Y(n_1683)
);

INVx5_ASAP7_75t_L g1684 ( 
.A(n_1463),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1380),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1555),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1682),
.B(n_909),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1523),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1543),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1676),
.B(n_949),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1607),
.B(n_930),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1683),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1533),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1582),
.B(n_996),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1518),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1522),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1627),
.B(n_1622),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1545),
.Y(n_1698)
);

INVx4_ASAP7_75t_L g1699 ( 
.A(n_1549),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1591),
.B(n_998),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1563),
.B(n_932),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1528),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1671),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1672),
.Y(n_1704)
);

INVx5_ASAP7_75t_L g1705 ( 
.A(n_1535),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1616),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1629),
.B(n_1579),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1517),
.Y(n_1708)
);

INVx8_ASAP7_75t_L g1709 ( 
.A(n_1651),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1620),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1563),
.B(n_1011),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1596),
.B(n_1539),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1542),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1568),
.B(n_1194),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1539),
.B(n_978),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1559),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1534),
.Y(n_1717)
);

INVx4_ASAP7_75t_SL g1718 ( 
.A(n_1651),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1548),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1585),
.B(n_979),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1661),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1673),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1617),
.B(n_1624),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1585),
.B(n_985),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1674),
.B(n_1049),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1569),
.Y(n_1726)
);

BUFx10_ASAP7_75t_L g1727 ( 
.A(n_1525),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1544),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1554),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1589),
.B(n_988),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1609),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1662),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1610),
.Y(n_1733)
);

INVx4_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1520),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1565),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1526),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1589),
.B(n_989),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1521),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1589),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1519),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1681),
.B(n_1141),
.Y(n_1742)
);

INVx5_ASAP7_75t_L g1743 ( 
.A(n_1594),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1604),
.B(n_1021),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1594),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1675),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1602),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1623),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1679),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1642),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1649),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1586),
.A2(n_1028),
.B1(n_1074),
.B2(n_1055),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1594),
.B(n_993),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1540),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1546),
.A2(n_1075),
.B1(n_1092),
.B2(n_1074),
.Y(n_1755)
);

INVx6_ASAP7_75t_L g1756 ( 
.A(n_1631),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1641),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1631),
.Y(n_1758)
);

BUFx4f_ASAP7_75t_L g1759 ( 
.A(n_1637),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1648),
.Y(n_1760)
);

INVx5_ASAP7_75t_L g1761 ( 
.A(n_1631),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1583),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1527),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1599),
.B(n_1024),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1646),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1614),
.Y(n_1766)
);

AND2x6_ASAP7_75t_L g1767 ( 
.A(n_1632),
.B(n_1075),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1601),
.B(n_1025),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1644),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1603),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1647),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1556),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1531),
.Y(n_1773)
);

OR2x2_ASAP7_75t_SL g1774 ( 
.A(n_1587),
.B(n_1072),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1597),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1639),
.B(n_1003),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1608),
.B(n_1027),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1680),
.A2(n_1157),
.B1(n_1168),
.B2(n_1092),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1572),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1572),
.Y(n_1780)
);

AND2x6_ASAP7_75t_L g1781 ( 
.A(n_1529),
.B(n_1157),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1538),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1541),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1547),
.B(n_1168),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1619),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1625),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1644),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1634),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1670),
.A2(n_1034),
.B(n_1031),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1684),
.B(n_1007),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1626),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1640),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1612),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1639),
.B(n_1008),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1630),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1573),
.A2(n_1239),
.B1(n_1235),
.B2(n_995),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1635),
.B(n_1010),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1613),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1638),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1593),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1600),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1656),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1658),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1660),
.Y(n_1804)
);

NOR3xp33_ASAP7_75t_L g1805 ( 
.A(n_1557),
.B(n_1248),
.C(n_1216),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1636),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1551),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1561),
.B(n_1018),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1643),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1584),
.B(n_1019),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1615),
.Y(n_1811)
);

INVx5_ASAP7_75t_L g1812 ( 
.A(n_1636),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1628),
.A2(n_1564),
.B1(n_1567),
.B2(n_1566),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1550),
.B(n_1020),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1654),
.Y(n_1815)
);

INVx5_ASAP7_75t_L g1816 ( 
.A(n_1667),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1552),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1532),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1592),
.B(n_1022),
.Y(n_1819)
);

AND2x6_ASAP7_75t_L g1820 ( 
.A(n_1590),
.B(n_1235),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1618),
.Y(n_1821)
);

NOR3xp33_ASAP7_75t_L g1822 ( 
.A(n_1558),
.B(n_1029),
.C(n_1026),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1578),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1621),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1570),
.A2(n_1033),
.B1(n_1035),
.B2(n_1030),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1553),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1580),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1530),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_SL g1829 ( 
.A(n_1537),
.B(n_1063),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1645),
.B(n_1039),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1605),
.B(n_1063),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1571),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1650),
.B(n_1042),
.Y(n_1833)
);

NAND2x1p5_ASAP7_75t_L g1834 ( 
.A(n_1669),
.B(n_1239),
.Y(n_1834)
);

OR2x6_ASAP7_75t_L g1835 ( 
.A(n_1633),
.B(n_1009),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1560),
.B(n_1070),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1655),
.B(n_1043),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1536),
.B(n_1070),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1606),
.B(n_1595),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1659),
.Y(n_1840)
);

NAND2xp33_ASAP7_75t_L g1841 ( 
.A(n_1562),
.B(n_1069),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1574),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1611),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1652),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1665),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1576),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1577),
.B(n_1044),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1581),
.B(n_1046),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1588),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1666),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1653),
.Y(n_1851)
);

AND2x6_ASAP7_75t_L g1852 ( 
.A(n_1657),
.B(n_973),
.Y(n_1852)
);

CKINVDCx20_ASAP7_75t_R g1853 ( 
.A(n_1678),
.Y(n_1853)
);

AND2x6_ASAP7_75t_L g1854 ( 
.A(n_1598),
.B(n_973),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1663),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1668),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1664),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1543),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1543),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1528),
.Y(n_1860)
);

OR2x6_ASAP7_75t_L g1861 ( 
.A(n_1524),
.B(n_1013),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1543),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1528),
.B(n_1057),
.Y(n_1863)
);

BUFx10_ASAP7_75t_L g1864 ( 
.A(n_1545),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1543),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1543),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1543),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1682),
.B(n_1062),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1528),
.B(n_1064),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1685),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1607),
.A2(n_1066),
.B1(n_1073),
.B2(n_1065),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1682),
.B(n_1076),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1523),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1575),
.A2(n_1110),
.B1(n_1127),
.B2(n_1080),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1685),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1523),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1543),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1682),
.B(n_1077),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1523),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1523),
.Y(n_1880)
);

BUFx4f_ASAP7_75t_L g1881 ( 
.A(n_1524),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1685),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1582),
.B(n_1048),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1528),
.B(n_1079),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1528),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1523),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1627),
.B(n_1082),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1523),
.Y(n_1888)
);

AND2x2_ASAP7_75t_SL g1889 ( 
.A(n_1524),
.B(n_1036),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1716),
.B(n_1084),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1701),
.B(n_1085),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1707),
.B(n_1086),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1697),
.B(n_1087),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1735),
.A2(n_1052),
.B(n_1050),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1695),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1711),
.B(n_1095),
.Y(n_1896)
);

NAND2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1705),
.B(n_1006),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1712),
.B(n_1690),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1714),
.B(n_1097),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1706),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1710),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1705),
.B(n_1702),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1744),
.A2(n_1822),
.B1(n_1805),
.B2(n_1889),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1708),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1726),
.B(n_1102),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1722),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1758),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1696),
.B(n_1108),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1858),
.B(n_1109),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1881),
.B(n_1112),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1859),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1687),
.A2(n_1113),
.B1(n_1116),
.B2(n_1114),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1862),
.B(n_1118),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1865),
.B(n_1119),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1866),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1867),
.B(n_1122),
.Y(n_1916)
);

OR2x6_ASAP7_75t_SL g1917 ( 
.A(n_1713),
.B(n_1124),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_L g1918 ( 
.A(n_1813),
.B(n_1054),
.C(n_1053),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1836),
.B(n_1130),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1877),
.B(n_1131),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1688),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1736),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1779),
.B(n_1137),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1806),
.B(n_1142),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1693),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1812),
.B(n_1144),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1732),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1814),
.B(n_1151),
.Y(n_1928)
);

NAND2xp33_ASAP7_75t_L g1929 ( 
.A(n_1854),
.B(n_1153),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1812),
.B(n_1155),
.Y(n_1930)
);

NAND2x1_ASAP7_75t_L g1931 ( 
.A(n_1756),
.B(n_1006),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1838),
.B(n_1110),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1769),
.B(n_1159),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1723),
.B(n_1160),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1861),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1787),
.B(n_1161),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1860),
.B(n_1163),
.Y(n_1937)
);

OAI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1728),
.A2(n_1129),
.B1(n_1139),
.B2(n_1091),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1709),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1743),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1743),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1754),
.A2(n_1061),
.B(n_1059),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1830),
.A2(n_1136),
.B1(n_1164),
.B2(n_1162),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1873),
.A2(n_1139),
.B1(n_1165),
.B2(n_1129),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1719),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1737),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1757),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1704),
.B(n_1180),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1876),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1879),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1725),
.B(n_1742),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1739),
.A2(n_1071),
.B(n_1067),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1887),
.B(n_1184),
.Y(n_1953)
);

BUFx5_ASAP7_75t_L g1954 ( 
.A(n_1852),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1694),
.B(n_1189),
.Y(n_1955)
);

NOR2xp67_ASAP7_75t_L g1956 ( 
.A(n_1698),
.B(n_90),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1694),
.B(n_1190),
.Y(n_1957)
);

NAND2xp33_ASAP7_75t_L g1958 ( 
.A(n_1740),
.B(n_1197),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1760),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1802),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1747),
.B(n_1748),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1700),
.B(n_1883),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1880),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1886),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1888),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1883),
.B(n_1196),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1804),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1703),
.B(n_1198),
.Y(n_1968)
);

BUFx12f_ASAP7_75t_L g1969 ( 
.A(n_1864),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1803),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1870),
.B(n_1201),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1741),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_SL g1973 ( 
.A(n_1740),
.B(n_1164),
.Y(n_1973)
);

BUFx8_ASAP7_75t_L g1974 ( 
.A(n_1882),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1746),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1743),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1871),
.B(n_1202),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1749),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1750),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1751),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1772),
.Y(n_1981)
);

OAI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1835),
.A2(n_1205),
.B1(n_1208),
.B2(n_1204),
.Y(n_1982)
);

BUFx5_ASAP7_75t_L g1983 ( 
.A(n_1852),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1764),
.B(n_1209),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1782),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1764),
.B(n_1211),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1734),
.B(n_1212),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1775),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1785),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1786),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1768),
.B(n_1213),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1795),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1791),
.Y(n_1993)
);

NOR2xp67_ASAP7_75t_SL g1994 ( 
.A(n_1762),
.B(n_1279),
.Y(n_1994)
);

INVx4_ASAP7_75t_L g1995 ( 
.A(n_1793),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1799),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1809),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1815),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1777),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1745),
.Y(n_2000)
);

BUFx5_ASAP7_75t_L g2001 ( 
.A(n_1852),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1793),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1823),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1868),
.A2(n_1222),
.B1(n_1224),
.B2(n_1221),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1776),
.B(n_1227),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1794),
.B(n_1232),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1715),
.B(n_1233),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1798),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1780),
.B(n_1234),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1872),
.B(n_1243),
.Y(n_2010)
);

AND2x6_ASAP7_75t_SL g2011 ( 
.A(n_1839),
.B(n_1078),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1765),
.B(n_1242),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_SL g2013 ( 
.A(n_1745),
.B(n_1243),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1761),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1847),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1771),
.B(n_1250),
.Y(n_2016)
);

OR2x6_ASAP7_75t_L g2017 ( 
.A(n_1699),
.B(n_1174),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1767),
.B(n_1755),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1827),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1878),
.A2(n_1259),
.B1(n_1260),
.B2(n_1254),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1885),
.B(n_1686),
.Y(n_2021)
);

AND3x1_ASAP7_75t_L g2022 ( 
.A(n_1848),
.B(n_1275),
.C(n_1273),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1752),
.B(n_1261),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1796),
.B(n_1263),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1781),
.B(n_1264),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1770),
.B(n_1265),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1717),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1825),
.B(n_1272),
.Y(n_2028)
);

NAND3xp33_ASAP7_75t_L g2029 ( 
.A(n_1800),
.B(n_1045),
.C(n_1006),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_SL g2030 ( 
.A(n_1761),
.B(n_1266),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1843),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1721),
.B(n_1278),
.Y(n_2032)
);

A2O1A1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1801),
.A2(n_1200),
.B(n_1210),
.C(n_1175),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1756),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1807),
.Y(n_2035)
);

O2A1O1Ixp5_ASAP7_75t_L g2036 ( 
.A1(n_1720),
.A2(n_1200),
.B(n_1210),
.C(n_1175),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1855),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_1840),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_1821),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1831),
.B(n_1083),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1874),
.B(n_1089),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1784),
.B(n_1090),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1817),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1840),
.B(n_1093),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1788),
.Y(n_2045)
);

INVx8_ASAP7_75t_L g2046 ( 
.A(n_1820),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1828),
.B(n_1096),
.Y(n_2047)
);

INVx8_ASAP7_75t_L g2048 ( 
.A(n_1820),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1792),
.B(n_1098),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1884),
.B(n_1101),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1774),
.A2(n_1219),
.B1(n_1236),
.B2(n_1217),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1773),
.A2(n_1107),
.B1(n_1111),
.B2(n_1103),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1761),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1826),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1834),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1863),
.B(n_1115),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1763),
.A2(n_1120),
.B1(n_1126),
.B2(n_1123),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1869),
.B(n_1833),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1842),
.B(n_1134),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1724),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1730),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_1824),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1846),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1837),
.B(n_1148),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1808),
.B(n_1158),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1738),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1849),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1797),
.B(n_1166),
.Y(n_2068)
);

AO22x1_ASAP7_75t_L g2069 ( 
.A1(n_1832),
.A2(n_1818),
.B1(n_1783),
.B2(n_1842),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1851),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1729),
.B(n_1167),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1853),
.A2(n_1171),
.B1(n_1172),
.B2(n_1170),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1753),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1816),
.B(n_1179),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1816),
.B(n_1181),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1810),
.B(n_1182),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1819),
.B(n_1183),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1789),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1856),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1766),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1850),
.B(n_1185),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1857),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1845),
.B(n_1268),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1790),
.Y(n_2084)
);

INVx3_ASAP7_75t_L g2085 ( 
.A(n_1845),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1718),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1718),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1844),
.Y(n_2088)
);

BUFx8_ASAP7_75t_L g2089 ( 
.A(n_1731),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1759),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1733),
.B(n_1214),
.Y(n_2091)
);

INVxp67_ASAP7_75t_L g2092 ( 
.A(n_1811),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1727),
.B(n_1220),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1841),
.B(n_1223),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1744),
.A2(n_1150),
.B1(n_1154),
.B2(n_1105),
.Y(n_2095)
);

NAND3xp33_ASAP7_75t_L g2096 ( 
.A(n_1778),
.B(n_1099),
.C(n_1045),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1707),
.B(n_1229),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1695),
.Y(n_2098)
);

AOI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1691),
.A2(n_1231),
.B1(n_1237),
.B2(n_1230),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1701),
.B(n_1240),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_SL g2101 ( 
.A(n_1719),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1707),
.B(n_1252),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_1691),
.A2(n_1256),
.B1(n_1262),
.B2(n_1253),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1707),
.B(n_1274),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1689),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1707),
.B(n_1271),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1695),
.Y(n_2107)
);

NOR3xp33_ASAP7_75t_L g2108 ( 
.A(n_1691),
.B(n_1247),
.C(n_1245),
.Y(n_2108)
);

INVx4_ASAP7_75t_L g2109 ( 
.A(n_1705),
.Y(n_2109)
);

NOR3xp33_ASAP7_75t_L g2110 ( 
.A(n_1691),
.B(n_1267),
.C(n_1251),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_1744),
.A2(n_1150),
.B1(n_1154),
.B2(n_1105),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1707),
.B(n_1274),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_1744),
.A2(n_1154),
.B1(n_1150),
.B2(n_1099),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1707),
.B(n_1154),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1707),
.B(n_1267),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_1701),
.B(n_1269),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_1875),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1754),
.A2(n_1274),
.B(n_1),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_1707),
.B(n_90),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1707),
.B(n_1274),
.Y(n_2120)
);

AND2x4_ASAP7_75t_SL g2121 ( 
.A(n_1692),
.B(n_1045),
.Y(n_2121)
);

INVx4_ASAP7_75t_L g2122 ( 
.A(n_1705),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1707),
.B(n_1),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1707),
.B(n_898),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1707),
.B(n_1),
.Y(n_2125)
);

OR2x6_ASAP7_75t_L g2126 ( 
.A(n_1709),
.B(n_1099),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1689),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1707),
.B(n_1121),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1695),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1688),
.A2(n_1156),
.B1(n_1255),
.B2(n_1121),
.Y(n_2130)
);

INVx2_ASAP7_75t_SL g2131 ( 
.A(n_1705),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1705),
.Y(n_2132)
);

BUFx10_ASAP7_75t_L g2133 ( 
.A(n_1692),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1705),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1707),
.B(n_901),
.Y(n_2135)
);

INVx4_ASAP7_75t_L g2136 ( 
.A(n_1705),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1691),
.A2(n_1255),
.B1(n_92),
.B2(n_93),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1707),
.B(n_91),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1692),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1707),
.B(n_92),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1707),
.B(n_3),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1707),
.B(n_93),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_1707),
.B(n_94),
.Y(n_2143)
);

O2A1O1Ixp5_ASAP7_75t_L g2144 ( 
.A1(n_1800),
.A2(n_96),
.B(n_97),
.C(n_95),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1754),
.A2(n_4),
.B(n_5),
.Y(n_2145)
);

O2A1O1Ixp5_ASAP7_75t_L g2146 ( 
.A1(n_1800),
.A2(n_98),
.B(n_99),
.C(n_97),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1691),
.A2(n_99),
.B1(n_100),
.B2(n_98),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1707),
.B(n_7),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1689),
.Y(n_2149)
);

OAI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_1829),
.A2(n_102),
.B1(n_103),
.B2(n_101),
.Y(n_2150)
);

AOI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_1691),
.A2(n_102),
.B1(n_103),
.B2(n_101),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1707),
.B(n_7),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1689),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_1705),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1707),
.B(n_8),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_1707),
.B(n_104),
.Y(n_2156)
);

AND2x6_ASAP7_75t_L g2157 ( 
.A(n_1702),
.B(n_104),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1695),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1707),
.B(n_8),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1695),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_SL g2161 ( 
.A(n_1719),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1707),
.B(n_8),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_1707),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1689),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1689),
.Y(n_2165)
);

INVx4_ASAP7_75t_L g2166 ( 
.A(n_1705),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1707),
.B(n_8),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1695),
.Y(n_2168)
);

INVx4_ASAP7_75t_L g2169 ( 
.A(n_1705),
.Y(n_2169)
);

NAND2xp33_ASAP7_75t_L g2170 ( 
.A(n_1702),
.B(n_9),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_1692),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1707),
.B(n_9),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1707),
.B(n_106),
.Y(n_2173)
);

A2O1A1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_1723),
.A2(n_108),
.B(n_109),
.C(n_107),
.Y(n_2174)
);

NOR2xp67_ASAP7_75t_L g2175 ( 
.A(n_1806),
.B(n_108),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1695),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1707),
.B(n_108),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1707),
.B(n_110),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1695),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1707),
.B(n_897),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1695),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1707),
.B(n_110),
.Y(n_2182)
);

INVx8_ASAP7_75t_L g2183 ( 
.A(n_1705),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1689),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1707),
.B(n_111),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1707),
.B(n_111),
.Y(n_2186)
);

AND2x4_ASAP7_75t_L g2187 ( 
.A(n_1705),
.B(n_111),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1758),
.Y(n_2188)
);

BUFx5_ASAP7_75t_L g2189 ( 
.A(n_1852),
.Y(n_2189)
);

NOR2x1p5_ASAP7_75t_L g2190 ( 
.A(n_1719),
.B(n_112),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1689),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1716),
.B(n_11),
.Y(n_2192)
);

OR2x6_ASAP7_75t_L g2193 ( 
.A(n_1709),
.B(n_113),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1716),
.B(n_11),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_1705),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_SL g2196 ( 
.A(n_1719),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1716),
.B(n_11),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1695),
.Y(n_2198)
);

NAND3xp33_ASAP7_75t_L g2199 ( 
.A(n_1778),
.B(n_115),
.C(n_114),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1716),
.B(n_12),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1707),
.B(n_114),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_1754),
.A2(n_12),
.B(n_13),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1707),
.B(n_116),
.Y(n_2203)
);

OAI221xp5_ASAP7_75t_L g2204 ( 
.A1(n_1707),
.A2(n_118),
.B1(n_119),
.B2(n_117),
.C(n_116),
.Y(n_2204)
);

INVx8_ASAP7_75t_L g2205 ( 
.A(n_1705),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1707),
.B(n_117),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1689),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1707),
.B(n_117),
.Y(n_2208)
);

INVx3_ASAP7_75t_L g2209 ( 
.A(n_1705),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1716),
.B(n_12),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1716),
.B(n_13),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1689),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1689),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1716),
.B(n_13),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_2133),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1921),
.Y(n_2216)
);

AO21x1_ASAP7_75t_L g2217 ( 
.A1(n_2051),
.A2(n_123),
.B(n_121),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_SL g2218 ( 
.A(n_1932),
.B(n_123),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2163),
.B(n_124),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2163),
.B(n_125),
.Y(n_2220)
);

INVx1_ASAP7_75t_SL g2221 ( 
.A(n_2038),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1898),
.B(n_126),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2183),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1927),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1951),
.B(n_126),
.Y(n_2225)
);

OR2x6_ASAP7_75t_L g2226 ( 
.A(n_2183),
.B(n_128),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1907),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2044),
.B(n_129),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1997),
.Y(n_2229)
);

OR2x6_ASAP7_75t_L g2230 ( 
.A(n_2205),
.B(n_129),
.Y(n_2230)
);

BUFx12f_ASAP7_75t_L g2231 ( 
.A(n_1969),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_2078),
.A2(n_131),
.B(n_130),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_1923),
.A2(n_131),
.B(n_130),
.Y(n_2233)
);

BUFx12f_ASAP7_75t_L g2234 ( 
.A(n_1974),
.Y(n_2234)
);

AOI21x1_ASAP7_75t_L g2235 ( 
.A1(n_2018),
.A2(n_134),
.B(n_133),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_1962),
.A2(n_134),
.B1(n_135),
.B2(n_133),
.Y(n_2236)
);

CKINVDCx20_ASAP7_75t_R g2237 ( 
.A(n_2117),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2115),
.B(n_135),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2100),
.B(n_136),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2047),
.B(n_137),
.Y(n_2240)
);

BUFx4f_ASAP7_75t_L g2241 ( 
.A(n_2193),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2030),
.B(n_1982),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1907),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2205),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_1928),
.B(n_137),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2040),
.B(n_138),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2124),
.B(n_139),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2009),
.A2(n_2112),
.B(n_2104),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2120),
.A2(n_141),
.B(n_140),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1935),
.B(n_141),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1925),
.Y(n_2251)
);

NOR2x1_ASAP7_75t_L g2252 ( 
.A(n_2109),
.B(n_894),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2135),
.B(n_142),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2128),
.A2(n_144),
.B(n_143),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2012),
.A2(n_144),
.B(n_143),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2016),
.A2(n_144),
.B(n_143),
.Y(n_2256)
);

CKINVDCx11_ASAP7_75t_R g2257 ( 
.A(n_1917),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2180),
.B(n_145),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_1935),
.B(n_146),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_1890),
.A2(n_149),
.B(n_147),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_1891),
.A2(n_150),
.B1(n_151),
.B2(n_149),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2116),
.B(n_152),
.Y(n_2262)
);

OAI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2126),
.A2(n_154),
.B1(n_155),
.B2(n_153),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_1919),
.B(n_155),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1900),
.B(n_1901),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2118),
.A2(n_157),
.B(n_156),
.Y(n_2266)
);

AOI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_1905),
.A2(n_1909),
.B(n_1908),
.Y(n_2267)
);

BUFx4f_ASAP7_75t_L g2268 ( 
.A(n_2193),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1911),
.B(n_1915),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_1907),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_1896),
.A2(n_159),
.B1(n_160),
.B2(n_158),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2188),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_1913),
.A2(n_161),
.B(n_160),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_1913),
.A2(n_162),
.B(n_161),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_1914),
.A2(n_163),
.B(n_162),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_1916),
.A2(n_164),
.B(n_163),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_1920),
.A2(n_165),
.B(n_164),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1949),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_2188),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1950),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1998),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2114),
.A2(n_1975),
.B(n_1972),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2022),
.A2(n_168),
.B1(n_169),
.B2(n_167),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_1978),
.A2(n_169),
.B(n_168),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1963),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_2027),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2105),
.B(n_2127),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_1942),
.A2(n_170),
.B(n_169),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_1942),
.A2(n_171),
.B(n_170),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_1904),
.A2(n_172),
.B(n_171),
.Y(n_2290)
);

AOI21x1_ASAP7_75t_L g2291 ( 
.A1(n_2130),
.A2(n_1944),
.B(n_1938),
.Y(n_2291)
);

NOR2x1p5_ASAP7_75t_SL g2292 ( 
.A(n_1954),
.B(n_173),
.Y(n_2292)
);

OAI21xp33_ASAP7_75t_L g2293 ( 
.A1(n_1899),
.A2(n_14),
.B(n_15),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2149),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2153),
.Y(n_2295)
);

BUFx8_ASAP7_75t_L g2296 ( 
.A(n_2101),
.Y(n_2296)
);

AOI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_1906),
.A2(n_175),
.B(n_174),
.Y(n_2297)
);

AOI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_1964),
.A2(n_175),
.B(n_174),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2164),
.B(n_2165),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2022),
.A2(n_176),
.B1(n_177),
.B2(n_175),
.Y(n_2300)
);

AOI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_1965),
.A2(n_178),
.B(n_177),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2032),
.Y(n_2302)
);

INVx5_ASAP7_75t_L g2303 ( 
.A(n_2157),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_1934),
.A2(n_14),
.B(n_15),
.Y(n_2304)
);

O2A1O1Ixp33_ASAP7_75t_L g2305 ( 
.A1(n_2138),
.A2(n_2142),
.B(n_2143),
.C(n_2140),
.Y(n_2305)
);

INVx4_ASAP7_75t_L g2306 ( 
.A(n_2046),
.Y(n_2306)
);

INVx3_ASAP7_75t_L g2307 ( 
.A(n_2122),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2064),
.A2(n_180),
.B(n_179),
.Y(n_2308)
);

INVx5_ASAP7_75t_L g2309 ( 
.A(n_2157),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2119),
.A2(n_183),
.B1(n_184),
.B2(n_181),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2156),
.A2(n_186),
.B1(n_187),
.B2(n_185),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1895),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2059),
.B(n_188),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2184),
.Y(n_2314)
);

INVxp67_ASAP7_75t_L g2315 ( 
.A(n_2042),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2191),
.B(n_189),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2207),
.B(n_190),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2212),
.B(n_2213),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2053),
.B(n_190),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1999),
.B(n_2097),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2102),
.B(n_191),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_2089),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2053),
.B(n_191),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_1929),
.A2(n_192),
.B(n_191),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2106),
.B(n_192),
.Y(n_2325)
);

AOI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2015),
.A2(n_194),
.B(n_193),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1946),
.B(n_195),
.Y(n_2327)
);

OR2x6_ASAP7_75t_L g2328 ( 
.A(n_2046),
.B(n_195),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_2188),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2094),
.A2(n_197),
.B(n_196),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1947),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_1897),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2122),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2098),
.Y(n_2334)
);

AOI21x1_ASAP7_75t_L g2335 ( 
.A1(n_1938),
.A2(n_198),
.B(n_197),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_1894),
.A2(n_199),
.B(n_198),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1897),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_1952),
.A2(n_200),
.B(n_199),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2036),
.A2(n_202),
.B(n_201),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1959),
.B(n_202),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_1960),
.B(n_1967),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2136),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2091),
.B(n_203),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1970),
.Y(n_2344)
);

AOI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_1979),
.A2(n_205),
.B(n_204),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2107),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_2139),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1981),
.B(n_205),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_1980),
.A2(n_207),
.B(n_206),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1985),
.B(n_206),
.Y(n_2350)
);

NOR2x1_ASAP7_75t_L g2351 ( 
.A(n_2166),
.B(n_895),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2123),
.B(n_208),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2125),
.B(n_208),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_1988),
.A2(n_210),
.B(n_209),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1989),
.Y(n_2355)
);

INVx11_ASAP7_75t_L g2356 ( 
.A(n_1974),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_1990),
.A2(n_210),
.B(n_209),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_1992),
.A2(n_212),
.B(n_211),
.Y(n_2358)
);

AOI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_1996),
.A2(n_213),
.B(n_212),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_1903),
.B(n_212),
.Y(n_2360)
);

BUFx3_ASAP7_75t_L g2361 ( 
.A(n_2171),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_2169),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2141),
.A2(n_215),
.B(n_214),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1993),
.Y(n_2364)
);

BUFx8_ASAP7_75t_L g2365 ( 
.A(n_2161),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2169),
.B(n_216),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2099),
.A2(n_218),
.B1(n_219),
.B2(n_217),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_1893),
.B(n_220),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2148),
.B(n_221),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2152),
.B(n_222),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_1922),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2155),
.A2(n_224),
.B(n_223),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2159),
.A2(n_224),
.B(n_223),
.Y(n_2373)
);

INVx4_ASAP7_75t_L g2374 ( 
.A(n_2048),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2017),
.Y(n_2375)
);

AOI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2162),
.A2(n_226),
.B(n_225),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2167),
.A2(n_226),
.B(n_225),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2014),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_2187),
.B(n_227),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2172),
.A2(n_229),
.B(n_228),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_1973),
.B(n_230),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2192),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2173),
.A2(n_231),
.B(n_230),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1918),
.B(n_231),
.Y(n_2384)
);

AOI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2177),
.A2(n_233),
.B(n_232),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2178),
.A2(n_2208),
.B(n_2185),
.Y(n_2386)
);

OAI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2103),
.A2(n_234),
.B1(n_235),
.B2(n_233),
.Y(n_2387)
);

OAI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_1953),
.A2(n_19),
.B(n_20),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2192),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2010),
.B(n_235),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2182),
.A2(n_238),
.B(n_236),
.Y(n_2391)
);

O2A1O1Ixp33_ASAP7_75t_SL g2392 ( 
.A1(n_2083),
.A2(n_240),
.B(n_241),
.C(n_239),
.Y(n_2392)
);

O2A1O1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2186),
.A2(n_240),
.B(n_241),
.C(n_239),
.Y(n_2393)
);

BUFx2_ASAP7_75t_L g2394 ( 
.A(n_2017),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2201),
.A2(n_2206),
.B(n_2203),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_1984),
.B(n_242),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2005),
.A2(n_243),
.B(n_242),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2129),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_2013),
.B(n_244),
.Y(n_2399)
);

A2O1A1Ixp33_ASAP7_75t_L g2400 ( 
.A1(n_2199),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_2400)
);

INVx4_ASAP7_75t_L g2401 ( 
.A(n_2048),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2006),
.A2(n_245),
.B(n_244),
.Y(n_2402)
);

BUFx12f_ASAP7_75t_L g2403 ( 
.A(n_1939),
.Y(n_2403)
);

INVx1_ASAP7_75t_SL g2404 ( 
.A(n_2008),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2194),
.Y(n_2405)
);

A2O1A1Ixp33_ASAP7_75t_L g2406 ( 
.A1(n_2199),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_2406)
);

AOI21xp5_ASAP7_75t_L g2407 ( 
.A1(n_2197),
.A2(n_248),
.B(n_247),
.Y(n_2407)
);

A2O1A1Ixp33_ASAP7_75t_L g2408 ( 
.A1(n_2145),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2200),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2210),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2134),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_1986),
.B(n_249),
.Y(n_2412)
);

AOI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_1971),
.A2(n_250),
.B1(n_251),
.B2(n_249),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2137),
.A2(n_252),
.B1(n_253),
.B2(n_251),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_L g2415 ( 
.A(n_2108),
.B(n_253),
.C(n_252),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2041),
.B(n_253),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2013),
.B(n_255),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2110),
.B(n_256),
.Y(n_2418)
);

INVxp67_ASAP7_75t_L g2419 ( 
.A(n_1994),
.Y(n_2419)
);

O2A1O1Ixp33_ASAP7_75t_L g2420 ( 
.A1(n_2033),
.A2(n_257),
.B(n_258),
.C(n_256),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2211),
.A2(n_258),
.B(n_257),
.Y(n_2421)
);

AOI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2214),
.A2(n_260),
.B(n_259),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2214),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2043),
.A2(n_261),
.B(n_260),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_1991),
.B(n_261),
.Y(n_2425)
);

OAI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2007),
.A2(n_2023),
.B(n_1944),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2204),
.A2(n_263),
.B1(n_264),
.B2(n_262),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2175),
.B(n_263),
.Y(n_2428)
);

AOI21xp5_ASAP7_75t_L g2429 ( 
.A1(n_2054),
.A2(n_267),
.B(n_266),
.Y(n_2429)
);

BUFx3_ASAP7_75t_L g2430 ( 
.A(n_1945),
.Y(n_2430)
);

BUFx4f_ASAP7_75t_L g2431 ( 
.A(n_2048),
.Y(n_2431)
);

INVx11_ASAP7_75t_L g2432 ( 
.A(n_2196),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2158),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2160),
.B(n_2168),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_1995),
.Y(n_2435)
);

A2O1A1Ixp33_ASAP7_75t_L g2436 ( 
.A1(n_2202),
.A2(n_27),
.B(n_24),
.C(n_26),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2176),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2179),
.B(n_270),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_2195),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2181),
.Y(n_2440)
);

INVxp67_ASAP7_75t_L g2441 ( 
.A(n_2093),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2209),
.B(n_271),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2198),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_2121),
.B(n_273),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2031),
.B(n_275),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_1956),
.B(n_276),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2150),
.B(n_277),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2025),
.B(n_277),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2096),
.A2(n_278),
.B(n_277),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2014),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_1940),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_1955),
.B(n_280),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2003),
.Y(n_2453)
);

AO21x1_ASAP7_75t_L g2454 ( 
.A1(n_2170),
.A2(n_282),
.B(n_281),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_1957),
.B(n_281),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2019),
.Y(n_2456)
);

A2O1A1Ixp33_ASAP7_75t_L g2457 ( 
.A1(n_2174),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_1940),
.Y(n_2458)
);

OAI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2147),
.A2(n_284),
.B1(n_285),
.B2(n_283),
.Y(n_2459)
);

A2O1A1Ixp33_ASAP7_75t_L g2460 ( 
.A1(n_2144),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2037),
.Y(n_2461)
);

BUFx2_ASAP7_75t_L g2462 ( 
.A(n_2039),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1966),
.B(n_283),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2082),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2151),
.A2(n_287),
.B1(n_288),
.B2(n_286),
.Y(n_2465)
);

AOI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2096),
.A2(n_287),
.B(n_286),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2029),
.A2(n_290),
.B(n_289),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2063),
.A2(n_291),
.B(n_290),
.Y(n_2468)
);

AOI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2067),
.A2(n_293),
.B(n_291),
.Y(n_2469)
);

A2O1A1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_2146),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_1941),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2070),
.A2(n_2079),
.B(n_2084),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2074),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_1892),
.A2(n_294),
.B(n_293),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2024),
.B(n_294),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_1977),
.B(n_294),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2058),
.A2(n_296),
.B(n_295),
.Y(n_2477)
);

HB1xp67_ASAP7_75t_L g2478 ( 
.A(n_2062),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2075),
.Y(n_2479)
);

AOI21xp5_ASAP7_75t_L g2480 ( 
.A1(n_2060),
.A2(n_299),
.B(n_298),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_1941),
.Y(n_2481)
);

AOI21xp5_ASAP7_75t_L g2482 ( 
.A1(n_2061),
.A2(n_302),
.B(n_301),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2028),
.B(n_303),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2382),
.B(n_2072),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_2441),
.B(n_2011),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2456),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2332),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2224),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_2241),
.B(n_1954),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2228),
.B(n_2190),
.Y(n_2490)
);

NOR3xp33_ASAP7_75t_SL g2491 ( 
.A(n_2322),
.B(n_1961),
.C(n_2021),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2281),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2389),
.B(n_2057),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2332),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2229),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2294),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2405),
.B(n_2052),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2302),
.B(n_2092),
.Y(n_2498)
);

NOR3xp33_ASAP7_75t_SL g2499 ( 
.A(n_2286),
.B(n_1987),
.C(n_1968),
.Y(n_2499)
);

HB1xp67_ASAP7_75t_L g2500 ( 
.A(n_2221),
.Y(n_2500)
);

OAI22xp5_ASAP7_75t_L g2501 ( 
.A1(n_2268),
.A2(n_2113),
.B1(n_2111),
.B2(n_2095),
.Y(n_2501)
);

AOI21x1_ASAP7_75t_L g2502 ( 
.A1(n_2291),
.A2(n_1931),
.B(n_1902),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2409),
.B(n_2410),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2295),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2303),
.B(n_1954),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_R g2506 ( 
.A(n_2237),
.B(n_2196),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2371),
.B(n_1910),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2303),
.B(n_1983),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2267),
.A2(n_2000),
.B(n_1958),
.Y(n_2509)
);

AOI33xp33_ASAP7_75t_L g2510 ( 
.A1(n_2225),
.A2(n_1943),
.A3(n_2035),
.B1(n_1912),
.B2(n_2020),
.B3(n_2004),
.Y(n_2510)
);

OR2x6_ASAP7_75t_L g2511 ( 
.A(n_2234),
.B(n_2069),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2309),
.B(n_1983),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_2309),
.B(n_1983),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2313),
.B(n_2085),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2332),
.Y(n_2515)
);

OR2x2_ASAP7_75t_L g2516 ( 
.A(n_2315),
.B(n_2085),
.Y(n_2516)
);

BUFx3_ASAP7_75t_L g2517 ( 
.A(n_2215),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2314),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2423),
.B(n_2071),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2240),
.B(n_2343),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_2309),
.B(n_1983),
.Y(n_2521)
);

BUFx12f_ASAP7_75t_L g2522 ( 
.A(n_2231),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2453),
.B(n_2002),
.Y(n_2523)
);

BUFx6f_ASAP7_75t_L g2524 ( 
.A(n_2337),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2218),
.B(n_2001),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2223),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2375),
.B(n_1948),
.Y(n_2527)
);

AOI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2248),
.A2(n_2073),
.B(n_2066),
.Y(n_2528)
);

CKINVDCx6p67_ASAP7_75t_R g2529 ( 
.A(n_2257),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2331),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2461),
.B(n_2219),
.Y(n_2531)
);

AOI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2282),
.A2(n_2034),
.B(n_2049),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2426),
.A2(n_1976),
.B(n_2081),
.Y(n_2533)
);

AO22x1_ASAP7_75t_L g2534 ( 
.A1(n_2296),
.A2(n_2132),
.B1(n_2154),
.B2(n_2131),
.Y(n_2534)
);

AND2x6_ASAP7_75t_SL g2535 ( 
.A(n_2226),
.B(n_2086),
.Y(n_2535)
);

O2A1O1Ixp5_ASAP7_75t_L g2536 ( 
.A1(n_2242),
.A2(n_1926),
.B(n_1930),
.C(n_1924),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2386),
.A2(n_1937),
.B(n_1936),
.Y(n_2537)
);

OR2x6_ASAP7_75t_SL g2538 ( 
.A(n_2356),
.B(n_2087),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2473),
.B(n_2050),
.Y(n_2539)
);

AOI21xp33_ASAP7_75t_L g2540 ( 
.A1(n_2305),
.A2(n_2055),
.B(n_2088),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2337),
.B(n_2001),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2479),
.B(n_2056),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2265),
.B(n_2068),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2269),
.B(n_2065),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2287),
.B(n_2076),
.Y(n_2545)
);

INVxp67_ASAP7_75t_L g2546 ( 
.A(n_2462),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2395),
.A2(n_1933),
.B(n_2080),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2312),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2342),
.B(n_2001),
.Y(n_2549)
);

HB1xp67_ASAP7_75t_L g2550 ( 
.A(n_2230),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2299),
.B(n_2077),
.Y(n_2551)
);

BUFx6f_ASAP7_75t_L g2552 ( 
.A(n_2342),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2318),
.B(n_2341),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2362),
.B(n_2001),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_SL g2555 ( 
.A(n_2431),
.B(n_2090),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2264),
.B(n_2045),
.Y(n_2556)
);

NOR2xp33_ASAP7_75t_L g2557 ( 
.A(n_2394),
.B(n_2026),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2245),
.B(n_2396),
.Y(n_2558)
);

BUFx4f_ASAP7_75t_SL g2559 ( 
.A(n_2296),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2355),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2334),
.Y(n_2561)
);

NAND2x1p5_ASAP7_75t_L g2562 ( 
.A(n_2244),
.B(n_2189),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2362),
.B(n_2189),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2346),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2412),
.B(n_2425),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2307),
.B(n_2189),
.Y(n_2566)
);

OR2x6_ASAP7_75t_L g2567 ( 
.A(n_2328),
.B(n_304),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2472),
.A2(n_306),
.B(n_305),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2364),
.Y(n_2569)
);

AOI21xp33_ASAP7_75t_L g2570 ( 
.A1(n_2262),
.A2(n_308),
.B(n_307),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_R g2571 ( 
.A(n_2365),
.B(n_307),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2435),
.Y(n_2572)
);

OAI21x1_ASAP7_75t_L g2573 ( 
.A1(n_2266),
.A2(n_311),
.B(n_310),
.Y(n_2573)
);

NAND2x1p5_ASAP7_75t_L g2574 ( 
.A(n_2306),
.B(n_314),
.Y(n_2574)
);

A2O1A1Ixp33_ASAP7_75t_L g2575 ( 
.A1(n_2293),
.A2(n_313),
.B(n_314),
.C(n_312),
.Y(n_2575)
);

INVx4_ASAP7_75t_L g2576 ( 
.A(n_2403),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2464),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2333),
.B(n_313),
.Y(n_2578)
);

INVx5_ASAP7_75t_L g2579 ( 
.A(n_2227),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2344),
.Y(n_2580)
);

INVx5_ASAP7_75t_L g2581 ( 
.A(n_2227),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2478),
.Y(n_2582)
);

NOR2xp67_ASAP7_75t_L g2583 ( 
.A(n_2419),
.B(n_316),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2320),
.B(n_317),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2398),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_SL g2586 ( 
.A(n_2430),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2239),
.B(n_318),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2360),
.B(n_319),
.Y(n_2588)
);

OAI21x1_ASAP7_75t_L g2589 ( 
.A1(n_2235),
.A2(n_321),
.B(n_320),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2433),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2227),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2434),
.A2(n_322),
.B(n_321),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2440),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2443),
.Y(n_2594)
);

AOI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2352),
.A2(n_324),
.B(n_323),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2353),
.A2(n_326),
.B(n_325),
.Y(n_2596)
);

OR2x6_ASAP7_75t_L g2597 ( 
.A(n_2374),
.B(n_2401),
.Y(n_2597)
);

CKINVDCx6p67_ASAP7_75t_R g2598 ( 
.A(n_2361),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2220),
.B(n_2246),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2243),
.Y(n_2600)
);

NOR2xp33_ASAP7_75t_L g2601 ( 
.A(n_2404),
.B(n_2384),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2432),
.Y(n_2602)
);

INVx4_ASAP7_75t_L g2603 ( 
.A(n_2378),
.Y(n_2603)
);

O2A1O1Ixp33_ASAP7_75t_L g2604 ( 
.A1(n_2418),
.A2(n_334),
.B(n_335),
.C(n_333),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2368),
.B(n_333),
.Y(n_2605)
);

OAI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2415),
.A2(n_337),
.B(n_336),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2437),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2216),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2243),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2222),
.B(n_341),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_2390),
.B(n_2347),
.Y(n_2611)
);

NOR3xp33_ASAP7_75t_L g2612 ( 
.A(n_2283),
.B(n_343),
.C(n_342),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2321),
.B(n_344),
.Y(n_2613)
);

AOI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2369),
.A2(n_346),
.B(n_345),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2325),
.B(n_346),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_L g2616 ( 
.A(n_2270),
.Y(n_2616)
);

AND2x4_ASAP7_75t_L g2617 ( 
.A(n_2439),
.B(n_347),
.Y(n_2617)
);

AOI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2370),
.A2(n_348),
.B(n_347),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2251),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2460),
.A2(n_351),
.B(n_349),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2450),
.B(n_349),
.Y(n_2621)
);

AOI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2470),
.A2(n_352),
.B(n_351),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2471),
.Y(n_2623)
);

INVx5_ASAP7_75t_L g2624 ( 
.A(n_2270),
.Y(n_2624)
);

BUFx6f_ASAP7_75t_L g2625 ( 
.A(n_2272),
.Y(n_2625)
);

AOI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2475),
.A2(n_354),
.B(n_353),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2471),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2272),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2442),
.Y(n_2629)
);

AOI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2428),
.A2(n_355),
.B(n_354),
.Y(n_2630)
);

NOR3xp33_ASAP7_75t_SL g2631 ( 
.A(n_2300),
.B(n_889),
.C(n_888),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2278),
.Y(n_2632)
);

A2O1A1Ixp33_ASAP7_75t_L g2633 ( 
.A1(n_2420),
.A2(n_356),
.B(n_357),
.C(n_355),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2471),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2238),
.B(n_356),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2442),
.B(n_2250),
.Y(n_2636)
);

A2O1A1Ixp33_ASAP7_75t_L g2637 ( 
.A1(n_2288),
.A2(n_360),
.B(n_361),
.C(n_358),
.Y(n_2637)
);

OAI22xp5_ASAP7_75t_SL g2638 ( 
.A1(n_2259),
.A2(n_362),
.B1(n_363),
.B2(n_360),
.Y(n_2638)
);

INVx3_ASAP7_75t_L g2639 ( 
.A(n_2481),
.Y(n_2639)
);

NOR3xp33_ASAP7_75t_L g2640 ( 
.A(n_2446),
.B(n_363),
.C(n_362),
.Y(n_2640)
);

BUFx6f_ASAP7_75t_L g2641 ( 
.A(n_2279),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2280),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_2481),
.B(n_364),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2451),
.B(n_2458),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2285),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2392),
.A2(n_366),
.B(n_365),
.Y(n_2646)
);

A2O1A1Ixp33_ASAP7_75t_L g2647 ( 
.A1(n_2289),
.A2(n_367),
.B(n_368),
.C(n_366),
.Y(n_2647)
);

OAI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2408),
.A2(n_368),
.B1(n_369),
.B2(n_367),
.Y(n_2648)
);

BUFx4f_ASAP7_75t_L g2649 ( 
.A(n_2411),
.Y(n_2649)
);

OR2x6_ASAP7_75t_L g2650 ( 
.A(n_2379),
.B(n_369),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2436),
.A2(n_372),
.B1(n_373),
.B2(n_371),
.Y(n_2651)
);

A2O1A1Ixp33_ASAP7_75t_L g2652 ( 
.A1(n_2324),
.A2(n_374),
.B(n_375),
.C(n_373),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2452),
.B(n_2455),
.Y(n_2653)
);

OR2x2_ASAP7_75t_L g2654 ( 
.A(n_2247),
.B(n_2253),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2261),
.A2(n_378),
.B1(n_379),
.B2(n_377),
.Y(n_2655)
);

AO32x1_ASAP7_75t_L g2656 ( 
.A1(n_2263),
.A2(n_2414),
.A3(n_2427),
.B1(n_2465),
.B2(n_2459),
.Y(n_2656)
);

OR2x6_ASAP7_75t_L g2657 ( 
.A(n_2252),
.B(n_379),
.Y(n_2657)
);

A2O1A1Ixp33_ASAP7_75t_L g2658 ( 
.A1(n_2304),
.A2(n_381),
.B(n_382),
.C(n_380),
.Y(n_2658)
);

BUFx2_ASAP7_75t_L g2659 ( 
.A(n_2279),
.Y(n_2659)
);

A2O1A1Ixp33_ASAP7_75t_L g2660 ( 
.A1(n_2388),
.A2(n_383),
.B(n_384),
.C(n_382),
.Y(n_2660)
);

OAI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2271),
.A2(n_384),
.B1(n_385),
.B2(n_383),
.Y(n_2661)
);

OR2x6_ASAP7_75t_L g2662 ( 
.A(n_2351),
.B(n_384),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2258),
.B(n_386),
.Y(n_2663)
);

OAI22xp5_ASAP7_75t_SL g2664 ( 
.A1(n_2413),
.A2(n_387),
.B1(n_388),
.B2(n_386),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2279),
.B(n_387),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2329),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2463),
.B(n_388),
.Y(n_2667)
);

NOR2x1_ASAP7_75t_R g2668 ( 
.A(n_2381),
.B(n_389),
.Y(n_2668)
);

OR2x2_ASAP7_75t_L g2669 ( 
.A(n_2316),
.B(n_389),
.Y(n_2669)
);

NOR3xp33_ASAP7_75t_SL g2670 ( 
.A(n_2367),
.B(n_896),
.C(n_895),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2217),
.B(n_390),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2483),
.B(n_392),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_2335),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2317),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2476),
.B(n_392),
.Y(n_2675)
);

INVx1_ASAP7_75t_SL g2676 ( 
.A(n_2444),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_2387),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2438),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2310),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2311),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2327),
.Y(n_2681)
);

AOI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_2416),
.A2(n_2466),
.B(n_2449),
.Y(n_2682)
);

OR2x6_ASAP7_75t_L g2683 ( 
.A(n_2399),
.B(n_394),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2454),
.B(n_394),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2400),
.A2(n_396),
.B(n_395),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2448),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2340),
.B(n_397),
.Y(n_2687)
);

AOI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2406),
.A2(n_400),
.B(n_399),
.Y(n_2688)
);

NAND2x2_ASAP7_75t_L g2689 ( 
.A(n_2348),
.B(n_399),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_2350),
.Y(n_2690)
);

OR2x6_ASAP7_75t_L g2691 ( 
.A(n_2417),
.B(n_400),
.Y(n_2691)
);

AO21x2_ASAP7_75t_L g2692 ( 
.A1(n_2447),
.A2(n_402),
.B(n_401),
.Y(n_2692)
);

OAI22x1_ASAP7_75t_L g2693 ( 
.A1(n_2366),
.A2(n_404),
.B1(n_405),
.B2(n_402),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2457),
.A2(n_2233),
.B1(n_2256),
.B2(n_2255),
.Y(n_2694)
);

AO32x2_ASAP7_75t_L g2695 ( 
.A1(n_2236),
.A2(n_410),
.A3(n_411),
.B1(n_409),
.B2(n_408),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2445),
.B(n_408),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2467),
.A2(n_412),
.B(n_409),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2319),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2323),
.Y(n_2699)
);

INVx4_ASAP7_75t_L g2700 ( 
.A(n_2292),
.Y(n_2700)
);

NAND2x1p5_ASAP7_75t_L g2701 ( 
.A(n_2407),
.B(n_418),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2308),
.B(n_414),
.Y(n_2702)
);

A2O1A1Ixp33_ASAP7_75t_L g2703 ( 
.A1(n_2393),
.A2(n_415),
.B(n_416),
.C(n_414),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2232),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2474),
.Y(n_2705)
);

HB1xp67_ASAP7_75t_L g2706 ( 
.A(n_2421),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2422),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_2249),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2468),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2260),
.A2(n_417),
.B(n_416),
.Y(n_2710)
);

A2O1A1Ixp33_ASAP7_75t_L g2711 ( 
.A1(n_2273),
.A2(n_419),
.B(n_420),
.C(n_418),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2274),
.B(n_418),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2275),
.B(n_419),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2276),
.B(n_420),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2277),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2469),
.Y(n_2716)
);

OAI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2383),
.A2(n_422),
.B1(n_423),
.B2(n_421),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2339),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2284),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2298),
.Y(n_2720)
);

A2O1A1Ixp33_ASAP7_75t_L g2721 ( 
.A1(n_2397),
.A2(n_424),
.B(n_425),
.C(n_423),
.Y(n_2721)
);

BUFx6f_ASAP7_75t_L g2722 ( 
.A(n_2254),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2385),
.A2(n_425),
.B1(n_426),
.B2(n_424),
.Y(n_2723)
);

A2O1A1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_2402),
.A2(n_426),
.B(n_427),
.C(n_424),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2326),
.B(n_427),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2363),
.B(n_427),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2301),
.Y(n_2727)
);

INVx6_ASAP7_75t_L g2728 ( 
.A(n_2477),
.Y(n_2728)
);

AND2x6_ASAP7_75t_L g2729 ( 
.A(n_2391),
.B(n_429),
.Y(n_2729)
);

AOI221xp5_ASAP7_75t_L g2730 ( 
.A1(n_2372),
.A2(n_432),
.B1(n_433),
.B2(n_431),
.C(n_430),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_L g2731 ( 
.A(n_2373),
.B(n_432),
.Y(n_2731)
);

A2O1A1Ixp33_ASAP7_75t_L g2732 ( 
.A1(n_2376),
.A2(n_433),
.B(n_434),
.C(n_432),
.Y(n_2732)
);

NAND3xp33_ASAP7_75t_L g2733 ( 
.A(n_2377),
.B(n_887),
.C(n_886),
.Y(n_2733)
);

OAI22xp5_ASAP7_75t_L g2734 ( 
.A1(n_2380),
.A2(n_436),
.B1(n_437),
.B2(n_435),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2330),
.A2(n_2338),
.B1(n_2336),
.B2(n_2480),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2482),
.B(n_438),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2290),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.Y(n_2737)
);

INVx4_ASAP7_75t_L g2738 ( 
.A(n_2297),
.Y(n_2738)
);

NAND2x1p5_ASAP7_75t_L g2739 ( 
.A(n_2345),
.B(n_443),
.Y(n_2739)
);

AND2x6_ASAP7_75t_L g2740 ( 
.A(n_2349),
.B(n_438),
.Y(n_2740)
);

INVx1_ASAP7_75t_SL g2741 ( 
.A(n_2354),
.Y(n_2741)
);

INVx6_ASAP7_75t_L g2742 ( 
.A(n_2357),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2358),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_L g2744 ( 
.A(n_2359),
.B(n_439),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2424),
.Y(n_2745)
);

O2A1O1Ixp5_ASAP7_75t_L g2746 ( 
.A1(n_2429),
.A2(n_441),
.B(n_442),
.C(n_440),
.Y(n_2746)
);

AO32x2_ASAP7_75t_L g2747 ( 
.A1(n_2700),
.A2(n_444),
.A3(n_445),
.B1(n_443),
.B2(n_441),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2553),
.B(n_441),
.Y(n_2748)
);

INVx5_ASAP7_75t_L g2749 ( 
.A(n_2567),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2503),
.B(n_443),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2486),
.Y(n_2751)
);

OAI21x1_ASAP7_75t_L g2752 ( 
.A1(n_2502),
.A2(n_447),
.B(n_446),
.Y(n_2752)
);

AO32x2_ASAP7_75t_L g2753 ( 
.A1(n_2638),
.A2(n_448),
.A3(n_449),
.B1(n_447),
.B2(n_446),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2520),
.B(n_448),
.Y(n_2754)
);

OAI21x1_ASAP7_75t_L g2755 ( 
.A1(n_2673),
.A2(n_450),
.B(n_449),
.Y(n_2755)
);

AO32x2_ASAP7_75t_L g2756 ( 
.A1(n_2664),
.A2(n_453),
.A3(n_454),
.B1(n_452),
.B2(n_451),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2488),
.B(n_454),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_R g2758 ( 
.A(n_2559),
.B(n_900),
.Y(n_2758)
);

AOI21x1_ASAP7_75t_L g2759 ( 
.A1(n_2525),
.A2(n_457),
.B(n_456),
.Y(n_2759)
);

OAI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2533),
.A2(n_459),
.B(n_458),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2582),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2485),
.B(n_459),
.Y(n_2762)
);

OAI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2718),
.A2(n_462),
.B(n_461),
.Y(n_2763)
);

AOI21x1_ASAP7_75t_L g2764 ( 
.A1(n_2505),
.A2(n_464),
.B(n_463),
.Y(n_2764)
);

BUFx3_ASAP7_75t_L g2765 ( 
.A(n_2517),
.Y(n_2765)
);

OAI21x1_ASAP7_75t_L g2766 ( 
.A1(n_2509),
.A2(n_466),
.B(n_465),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2492),
.B(n_2495),
.Y(n_2767)
);

AO31x2_ASAP7_75t_L g2768 ( 
.A1(n_2704),
.A2(n_467),
.A3(n_468),
.B(n_466),
.Y(n_2768)
);

INVx2_ASAP7_75t_SL g2769 ( 
.A(n_2649),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_L g2770 ( 
.A1(n_2508),
.A2(n_468),
.B(n_467),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2552),
.B(n_467),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2496),
.Y(n_2772)
);

AOI31xp67_ASAP7_75t_L g2773 ( 
.A1(n_2719),
.A2(n_470),
.A3(n_471),
.B(n_469),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_2500),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2548),
.Y(n_2775)
);

INVx5_ASAP7_75t_L g2776 ( 
.A(n_2567),
.Y(n_2776)
);

AOI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2682),
.A2(n_472),
.B(n_471),
.Y(n_2777)
);

OAI21x1_ASAP7_75t_L g2778 ( 
.A1(n_2512),
.A2(n_2521),
.B(n_2513),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2504),
.Y(n_2779)
);

NAND3x1_ASAP7_75t_L g2780 ( 
.A(n_2529),
.B(n_474),
.C(n_473),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2518),
.Y(n_2781)
);

INVx8_ASAP7_75t_L g2782 ( 
.A(n_2522),
.Y(n_2782)
);

OAI21x1_ASAP7_75t_L g2783 ( 
.A1(n_2541),
.A2(n_476),
.B(n_475),
.Y(n_2783)
);

AO31x2_ASAP7_75t_L g2784 ( 
.A1(n_2738),
.A2(n_478),
.A3(n_479),
.B(n_477),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2530),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2561),
.Y(n_2786)
);

OAI21x1_ASAP7_75t_L g2787 ( 
.A1(n_2715),
.A2(n_2532),
.B(n_2549),
.Y(n_2787)
);

INVx3_ASAP7_75t_L g2788 ( 
.A(n_2597),
.Y(n_2788)
);

AO31x2_ASAP7_75t_L g2789 ( 
.A1(n_2720),
.A2(n_481),
.A3(n_482),
.B(n_480),
.Y(n_2789)
);

INVx3_ASAP7_75t_L g2790 ( 
.A(n_2597),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2564),
.Y(n_2791)
);

OAI21x1_ASAP7_75t_L g2792 ( 
.A1(n_2554),
.A2(n_484),
.B(n_483),
.Y(n_2792)
);

OAI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2746),
.A2(n_485),
.B(n_484),
.Y(n_2793)
);

AO31x2_ASAP7_75t_L g2794 ( 
.A1(n_2727),
.A2(n_487),
.A3(n_488),
.B(n_486),
.Y(n_2794)
);

OAI21x1_ASAP7_75t_L g2795 ( 
.A1(n_2563),
.A2(n_487),
.B(n_486),
.Y(n_2795)
);

AO31x2_ASAP7_75t_L g2796 ( 
.A1(n_2745),
.A2(n_489),
.A3(n_490),
.B(n_488),
.Y(n_2796)
);

INVx4_ASAP7_75t_L g2797 ( 
.A(n_2598),
.Y(n_2797)
);

AND2x4_ASAP7_75t_L g2798 ( 
.A(n_2572),
.B(n_490),
.Y(n_2798)
);

OAI21x1_ASAP7_75t_L g2799 ( 
.A1(n_2705),
.A2(n_492),
.B(n_491),
.Y(n_2799)
);

OAI21x1_ASAP7_75t_L g2800 ( 
.A1(n_2566),
.A2(n_493),
.B(n_492),
.Y(n_2800)
);

INVx5_ASAP7_75t_L g2801 ( 
.A(n_2511),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2511),
.B(n_493),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2560),
.B(n_494),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2743),
.A2(n_496),
.B(n_495),
.Y(n_2804)
);

NOR2x1_ASAP7_75t_SL g2805 ( 
.A(n_2489),
.B(n_496),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2569),
.B(n_497),
.Y(n_2806)
);

AO31x2_ASAP7_75t_L g2807 ( 
.A1(n_2709),
.A2(n_498),
.A3(n_499),
.B(n_497),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2716),
.A2(n_502),
.B(n_501),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2577),
.B(n_501),
.Y(n_2809)
);

AOI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2707),
.A2(n_504),
.B(n_503),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2576),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2580),
.Y(n_2812)
);

AOI21xp5_ASAP7_75t_L g2813 ( 
.A1(n_2706),
.A2(n_505),
.B(n_504),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_SL g2814 ( 
.A(n_2552),
.B(n_505),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2528),
.A2(n_507),
.B(n_506),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2741),
.A2(n_509),
.B(n_508),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2550),
.B(n_508),
.Y(n_2817)
);

BUFx6f_ASAP7_75t_L g2818 ( 
.A(n_2579),
.Y(n_2818)
);

OAI21x1_ASAP7_75t_L g2819 ( 
.A1(n_2589),
.A2(n_511),
.B(n_510),
.Y(n_2819)
);

OAI21x1_ASAP7_75t_L g2820 ( 
.A1(n_2573),
.A2(n_511),
.B(n_510),
.Y(n_2820)
);

AOI221x1_ASAP7_75t_L g2821 ( 
.A1(n_2693),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.C(n_512),
.Y(n_2821)
);

AO31x2_ASAP7_75t_L g2822 ( 
.A1(n_2694),
.A2(n_515),
.A3(n_516),
.B(n_514),
.Y(n_2822)
);

OAI21x1_ASAP7_75t_L g2823 ( 
.A1(n_2562),
.A2(n_516),
.B(n_515),
.Y(n_2823)
);

INVx4_ASAP7_75t_L g2824 ( 
.A(n_2586),
.Y(n_2824)
);

OAI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2689),
.A2(n_517),
.B1(n_518),
.B2(n_516),
.Y(n_2825)
);

INVxp67_ASAP7_75t_L g2826 ( 
.A(n_2498),
.Y(n_2826)
);

OAI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2679),
.A2(n_518),
.B1(n_519),
.B2(n_517),
.Y(n_2827)
);

AOI21x1_ASAP7_75t_L g2828 ( 
.A1(n_2684),
.A2(n_518),
.B(n_517),
.Y(n_2828)
);

BUFx5_ASAP7_75t_L g2829 ( 
.A(n_2634),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2590),
.Y(n_2830)
);

OA21x2_ASAP7_75t_L g2831 ( 
.A1(n_2671),
.A2(n_522),
.B(n_521),
.Y(n_2831)
);

OAI21x1_ASAP7_75t_L g2832 ( 
.A1(n_2547),
.A2(n_524),
.B(n_523),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2593),
.Y(n_2833)
);

AOI211x1_ASAP7_75t_L g2834 ( 
.A1(n_2534),
.A2(n_527),
.B(n_528),
.C(n_526),
.Y(n_2834)
);

OAI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2733),
.A2(n_530),
.B(n_529),
.Y(n_2835)
);

BUFx4f_ASAP7_75t_SL g2836 ( 
.A(n_2602),
.Y(n_2836)
);

AO31x2_ASAP7_75t_L g2837 ( 
.A1(n_2659),
.A2(n_531),
.A3(n_532),
.B(n_530),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2594),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2506),
.Y(n_2839)
);

AO31x2_ASAP7_75t_L g2840 ( 
.A1(n_2666),
.A2(n_534),
.A3(n_535),
.B(n_533),
.Y(n_2840)
);

AO31x2_ASAP7_75t_L g2841 ( 
.A1(n_2575),
.A2(n_537),
.A3(n_538),
.B(n_536),
.Y(n_2841)
);

NOR2xp67_ASAP7_75t_L g2842 ( 
.A(n_2546),
.B(n_542),
.Y(n_2842)
);

NAND2x1p5_ASAP7_75t_L g2843 ( 
.A(n_2581),
.B(n_2624),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2677),
.A2(n_904),
.B1(n_538),
.B2(n_539),
.Y(n_2844)
);

OAI21x1_ASAP7_75t_L g2845 ( 
.A1(n_2639),
.A2(n_540),
.B(n_539),
.Y(n_2845)
);

OAI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2680),
.A2(n_541),
.B1(n_542),
.B2(n_540),
.Y(n_2846)
);

BUFx3_ASAP7_75t_L g2847 ( 
.A(n_2538),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2739),
.A2(n_544),
.B(n_543),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2656),
.A2(n_2653),
.B(n_2712),
.Y(n_2849)
);

OA21x2_ASAP7_75t_L g2850 ( 
.A1(n_2606),
.A2(n_547),
.B(n_546),
.Y(n_2850)
);

INVxp67_ASAP7_75t_L g2851 ( 
.A(n_2523),
.Y(n_2851)
);

OAI21x1_ASAP7_75t_L g2852 ( 
.A1(n_2698),
.A2(n_548),
.B(n_547),
.Y(n_2852)
);

OAI21x1_ASAP7_75t_L g2853 ( 
.A1(n_2735),
.A2(n_550),
.B(n_549),
.Y(n_2853)
);

AO31x2_ASAP7_75t_L g2854 ( 
.A1(n_2633),
.A2(n_552),
.A3(n_553),
.B(n_551),
.Y(n_2854)
);

OR2x2_ASAP7_75t_L g2855 ( 
.A(n_2565),
.B(n_552),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2490),
.B(n_2514),
.Y(n_2856)
);

OAI21x1_ASAP7_75t_L g2857 ( 
.A1(n_2585),
.A2(n_553),
.B(n_552),
.Y(n_2857)
);

BUFx2_ASAP7_75t_L g2858 ( 
.A(n_2526),
.Y(n_2858)
);

OAI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2703),
.A2(n_556),
.B(n_555),
.Y(n_2859)
);

BUFx12f_ASAP7_75t_L g2860 ( 
.A(n_2535),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2601),
.Y(n_2861)
);

BUFx2_ASAP7_75t_L g2862 ( 
.A(n_2603),
.Y(n_2862)
);

INVxp67_ASAP7_75t_SL g2863 ( 
.A(n_2629),
.Y(n_2863)
);

AND4x1_ASAP7_75t_L g2864 ( 
.A(n_2555),
.B(n_32),
.C(n_30),
.D(n_31),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2607),
.A2(n_559),
.B(n_558),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2608),
.A2(n_562),
.B(n_560),
.Y(n_2866)
);

BUFx12f_ASAP7_75t_L g2867 ( 
.A(n_2574),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2658),
.A2(n_564),
.B(n_563),
.Y(n_2868)
);

AOI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2699),
.A2(n_565),
.B(n_564),
.Y(n_2869)
);

OAI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2660),
.A2(n_566),
.B(n_565),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2619),
.Y(n_2871)
);

CKINVDCx20_ASAP7_75t_R g2872 ( 
.A(n_2571),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2484),
.B(n_567),
.Y(n_2873)
);

BUFx12f_ASAP7_75t_L g2874 ( 
.A(n_2657),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2497),
.B(n_569),
.Y(n_2875)
);

INVxp67_ASAP7_75t_SL g2876 ( 
.A(n_2591),
.Y(n_2876)
);

BUFx3_ASAP7_75t_L g2877 ( 
.A(n_2623),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2493),
.B(n_570),
.Y(n_2878)
);

OAI21x1_ASAP7_75t_L g2879 ( 
.A1(n_2632),
.A2(n_572),
.B(n_571),
.Y(n_2879)
);

OAI21x1_ASAP7_75t_L g2880 ( 
.A1(n_2642),
.A2(n_573),
.B(n_571),
.Y(n_2880)
);

OA21x2_ASAP7_75t_L g2881 ( 
.A1(n_2620),
.A2(n_2622),
.B(n_2568),
.Y(n_2881)
);

AO31x2_ASAP7_75t_L g2882 ( 
.A1(n_2637),
.A2(n_574),
.A3(n_576),
.B(n_573),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2645),
.Y(n_2883)
);

OAI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2537),
.A2(n_574),
.B(n_573),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2662),
.A2(n_576),
.B1(n_577),
.B2(n_574),
.Y(n_2885)
);

OA21x2_ASAP7_75t_L g2886 ( 
.A1(n_2685),
.A2(n_579),
.B(n_578),
.Y(n_2886)
);

OAI21x1_ASAP7_75t_L g2887 ( 
.A1(n_2701),
.A2(n_580),
.B(n_579),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2681),
.B(n_581),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2636),
.B(n_582),
.Y(n_2889)
);

OA21x2_ASAP7_75t_L g2890 ( 
.A1(n_2688),
.A2(n_584),
.B(n_583),
.Y(n_2890)
);

HB1xp67_ASAP7_75t_L g2891 ( 
.A(n_2627),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_2491),
.Y(n_2892)
);

AOI21xp5_ASAP7_75t_L g2893 ( 
.A1(n_2708),
.A2(n_586),
.B(n_585),
.Y(n_2893)
);

CKINVDCx8_ASAP7_75t_R g2894 ( 
.A(n_2650),
.Y(n_2894)
);

OAI21x1_ASAP7_75t_L g2895 ( 
.A1(n_2697),
.A2(n_589),
.B(n_588),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2588),
.B(n_588),
.Y(n_2896)
);

OAI21x1_ASAP7_75t_L g2897 ( 
.A1(n_2621),
.A2(n_589),
.B(n_588),
.Y(n_2897)
);

AND2x6_ASAP7_75t_L g2898 ( 
.A(n_2617),
.B(n_590),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2519),
.B(n_2674),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_SL g2900 ( 
.A1(n_2668),
.A2(n_591),
.B(n_590),
.Y(n_2900)
);

OAI21x1_ASAP7_75t_SL g2901 ( 
.A1(n_2604),
.A2(n_592),
.B(n_591),
.Y(n_2901)
);

AO31x2_ASAP7_75t_L g2902 ( 
.A1(n_2647),
.A2(n_595),
.A3(n_596),
.B(n_594),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2722),
.A2(n_595),
.B(n_594),
.Y(n_2903)
);

OAI21x1_ASAP7_75t_L g2904 ( 
.A1(n_2643),
.A2(n_596),
.B(n_594),
.Y(n_2904)
);

OAI21x1_ASAP7_75t_L g2905 ( 
.A1(n_2665),
.A2(n_598),
.B(n_597),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2558),
.B(n_598),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2516),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2644),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2531),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2600),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2690),
.B(n_599),
.Y(n_2911)
);

OAI21x1_ASAP7_75t_L g2912 ( 
.A1(n_2710),
.A2(n_602),
.B(n_601),
.Y(n_2912)
);

INVxp67_ASAP7_75t_L g2913 ( 
.A(n_2507),
.Y(n_2913)
);

NAND3xp33_ASAP7_75t_L g2914 ( 
.A(n_2675),
.B(n_604),
.C(n_603),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2678),
.B(n_604),
.Y(n_2915)
);

INVx5_ASAP7_75t_L g2916 ( 
.A(n_2600),
.Y(n_2916)
);

OAI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2652),
.A2(n_606),
.B(n_605),
.Y(n_2917)
);

NOR2x1_ASAP7_75t_SL g2918 ( 
.A(n_2683),
.B(n_607),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2583),
.B(n_2676),
.Y(n_2919)
);

AOI221x1_ASAP7_75t_L g2920 ( 
.A1(n_2540),
.A2(n_610),
.B1(n_611),
.B2(n_609),
.C(n_608),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2609),
.A2(n_613),
.B(n_612),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2609),
.A2(n_613),
.B(n_612),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2654),
.B(n_614),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2545),
.B(n_614),
.Y(n_2924)
);

OAI21x1_ASAP7_75t_L g2925 ( 
.A1(n_2536),
.A2(n_616),
.B(n_615),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2551),
.B(n_615),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2543),
.B(n_617),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2631),
.A2(n_618),
.B1(n_619),
.B2(n_617),
.Y(n_2928)
);

AO31x2_ASAP7_75t_L g2929 ( 
.A1(n_2737),
.A2(n_619),
.A3(n_620),
.B(n_618),
.Y(n_2929)
);

BUFx6f_ASAP7_75t_L g2930 ( 
.A(n_2487),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2599),
.B(n_620),
.Y(n_2931)
);

BUFx2_ASAP7_75t_L g2932 ( 
.A(n_2487),
.Y(n_2932)
);

OAI21x1_ASAP7_75t_L g2933 ( 
.A1(n_2646),
.A2(n_622),
.B(n_621),
.Y(n_2933)
);

OAI21x1_ASAP7_75t_L g2934 ( 
.A1(n_2713),
.A2(n_623),
.B(n_622),
.Y(n_2934)
);

OAI21x1_ASAP7_75t_L g2935 ( 
.A1(n_2714),
.A2(n_623),
.B(n_622),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2544),
.B(n_624),
.Y(n_2936)
);

BUFx3_ASAP7_75t_L g2937 ( 
.A(n_2487),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2611),
.B(n_625),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2494),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2539),
.B(n_626),
.Y(n_2940)
);

AOI22xp33_ASAP7_75t_L g2941 ( 
.A1(n_2612),
.A2(n_629),
.B1(n_630),
.B2(n_628),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2542),
.B(n_629),
.Y(n_2942)
);

AOI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2616),
.A2(n_631),
.B(n_629),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2605),
.B(n_631),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2527),
.B(n_631),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2494),
.B(n_632),
.Y(n_2946)
);

OAI21x1_ASAP7_75t_L g2947 ( 
.A1(n_2702),
.A2(n_634),
.B(n_632),
.Y(n_2947)
);

AO31x2_ASAP7_75t_L g2948 ( 
.A1(n_2648),
.A2(n_2651),
.A3(n_2711),
.B(n_2721),
.Y(n_2948)
);

OR2x6_ASAP7_75t_L g2949 ( 
.A(n_2691),
.B(n_637),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2584),
.B(n_638),
.Y(n_2950)
);

AO32x2_ASAP7_75t_L g2951 ( 
.A1(n_2655),
.A2(n_641),
.A3(n_642),
.B1(n_640),
.B2(n_639),
.Y(n_2951)
);

NAND2xp33_ASAP7_75t_R g2952 ( 
.A(n_2499),
.B(n_639),
.Y(n_2952)
);

OAI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2670),
.A2(n_644),
.B1(n_645),
.B2(n_643),
.Y(n_2953)
);

OAI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2724),
.A2(n_644),
.B(n_643),
.Y(n_2954)
);

AO32x2_ASAP7_75t_L g2955 ( 
.A1(n_2661),
.A2(n_648),
.A3(n_650),
.B1(n_647),
.B2(n_646),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2625),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2557),
.B(n_647),
.Y(n_2957)
);

OAI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2726),
.A2(n_2592),
.B(n_2626),
.Y(n_2958)
);

INVx5_ASAP7_75t_L g2959 ( 
.A(n_2628),
.Y(n_2959)
);

OAI21x1_ASAP7_75t_L g2960 ( 
.A1(n_2578),
.A2(n_652),
.B(n_651),
.Y(n_2960)
);

OAI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2732),
.A2(n_652),
.B(n_651),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2687),
.B(n_653),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2628),
.Y(n_2963)
);

CKINVDCx16_ASAP7_75t_R g2964 ( 
.A(n_2663),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2729),
.A2(n_655),
.B1(n_656),
.B2(n_653),
.Y(n_2965)
);

AOI221x1_ASAP7_75t_L g2966 ( 
.A1(n_2570),
.A2(n_659),
.B1(n_660),
.B2(n_658),
.C(n_657),
.Y(n_2966)
);

BUFx6f_ASAP7_75t_L g2967 ( 
.A(n_2515),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2641),
.Y(n_2968)
);

BUFx6f_ASAP7_75t_L g2969 ( 
.A(n_2524),
.Y(n_2969)
);

OAI21x1_ASAP7_75t_L g2970 ( 
.A1(n_2630),
.A2(n_660),
.B(n_659),
.Y(n_2970)
);

HB1xp67_ASAP7_75t_L g2971 ( 
.A(n_2761),
.Y(n_2971)
);

OAI21x1_ASAP7_75t_SL g2972 ( 
.A1(n_2918),
.A2(n_2596),
.B(n_2595),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2772),
.Y(n_2973)
);

HB1xp67_ASAP7_75t_L g2974 ( 
.A(n_2858),
.Y(n_2974)
);

INVxp67_ASAP7_75t_SL g2975 ( 
.A(n_2774),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2779),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2847),
.B(n_2524),
.Y(n_2977)
);

NAND2x1p5_ASAP7_75t_L g2978 ( 
.A(n_2797),
.B(n_2524),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_L g2979 ( 
.A1(n_2949),
.A2(n_2729),
.B1(n_2728),
.B2(n_2740),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2781),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2785),
.Y(n_2981)
);

INVx6_ASAP7_75t_L g2982 ( 
.A(n_2782),
.Y(n_2982)
);

OAI21x1_ASAP7_75t_L g2983 ( 
.A1(n_2787),
.A2(n_2618),
.B(n_2614),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2856),
.B(n_2909),
.Y(n_2984)
);

OAI21x1_ASAP7_75t_L g2985 ( 
.A1(n_2752),
.A2(n_2723),
.B(n_2717),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_L g2986 ( 
.A1(n_2778),
.A2(n_2734),
.B(n_2736),
.Y(n_2986)
);

INVx3_ASAP7_75t_L g2987 ( 
.A(n_2765),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2908),
.B(n_2692),
.Y(n_2988)
);

OAI22xp33_ASAP7_75t_L g2989 ( 
.A1(n_2894),
.A2(n_2686),
.B1(n_2728),
.B2(n_2556),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2907),
.B(n_2695),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2782),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2812),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2889),
.B(n_2695),
.Y(n_2993)
);

OR2x6_ASAP7_75t_L g2994 ( 
.A(n_2874),
.B(n_2725),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2751),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2830),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2833),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2775),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2838),
.Y(n_2999)
);

BUFx2_ASAP7_75t_L g3000 ( 
.A(n_2862),
.Y(n_3000)
);

AO21x2_ASAP7_75t_L g3001 ( 
.A1(n_2849),
.A2(n_2587),
.B(n_2610),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2786),
.Y(n_3002)
);

AOI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2919),
.A2(n_2672),
.B(n_2615),
.Y(n_3003)
);

OA21x2_ASAP7_75t_L g3004 ( 
.A1(n_2760),
.A2(n_2730),
.B(n_2696),
.Y(n_3004)
);

OAI21x1_ASAP7_75t_L g3005 ( 
.A1(n_2763),
.A2(n_2613),
.B(n_2501),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2767),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2791),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2898),
.A2(n_2731),
.B1(n_2640),
.B2(n_2744),
.Y(n_3008)
);

OAI21x1_ASAP7_75t_L g3009 ( 
.A1(n_2755),
.A2(n_2667),
.B(n_2635),
.Y(n_3009)
);

BUFx8_ASAP7_75t_L g3010 ( 
.A(n_2860),
.Y(n_3010)
);

NAND2x1p5_ASAP7_75t_L g3011 ( 
.A(n_2749),
.B(n_2669),
.Y(n_3011)
);

AOI22xp33_ASAP7_75t_L g3012 ( 
.A1(n_2898),
.A2(n_2740),
.B1(n_2742),
.B2(n_2510),
.Y(n_3012)
);

OAI21x1_ASAP7_75t_L g3013 ( 
.A1(n_2799),
.A2(n_662),
.B(n_661),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2871),
.Y(n_3014)
);

CKINVDCx20_ASAP7_75t_R g3015 ( 
.A(n_2872),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2883),
.Y(n_3016)
);

AO31x2_ASAP7_75t_L g3017 ( 
.A1(n_2920),
.A2(n_901),
.A3(n_665),
.B(n_666),
.Y(n_3017)
);

HB1xp67_ASAP7_75t_L g3018 ( 
.A(n_2891),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2766),
.A2(n_666),
.B(n_663),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2964),
.B(n_31),
.Y(n_3020)
);

INVx8_ASAP7_75t_L g3021 ( 
.A(n_2867),
.Y(n_3021)
);

O2A1O1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2825),
.A2(n_668),
.B(n_669),
.C(n_667),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2898),
.A2(n_669),
.B1(n_670),
.B2(n_668),
.Y(n_3023)
);

AO31x2_ASAP7_75t_L g3024 ( 
.A1(n_2805),
.A2(n_900),
.A3(n_670),
.B(n_671),
.Y(n_3024)
);

OAI21x1_ASAP7_75t_L g3025 ( 
.A1(n_2759),
.A2(n_672),
.B(n_671),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2876),
.Y(n_3026)
);

AND2x4_ASAP7_75t_L g3027 ( 
.A(n_2801),
.B(n_673),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_2758),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2863),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2899),
.Y(n_3030)
);

OA21x2_ASAP7_75t_L g3031 ( 
.A1(n_2958),
.A2(n_676),
.B(n_674),
.Y(n_3031)
);

OAI21x1_ASAP7_75t_L g3032 ( 
.A1(n_2804),
.A2(n_678),
.B(n_677),
.Y(n_3032)
);

AO31x2_ASAP7_75t_L g3033 ( 
.A1(n_2932),
.A2(n_680),
.A3(n_681),
.B(n_679),
.Y(n_3033)
);

OAI21x1_ASAP7_75t_L g3034 ( 
.A1(n_2808),
.A2(n_2832),
.B(n_2925),
.Y(n_3034)
);

OAI21x1_ASAP7_75t_L g3035 ( 
.A1(n_2843),
.A2(n_681),
.B(n_680),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2851),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2910),
.Y(n_3037)
);

CKINVDCx5p33_ASAP7_75t_R g3038 ( 
.A(n_2839),
.Y(n_3038)
);

CKINVDCx6p67_ASAP7_75t_R g3039 ( 
.A(n_2776),
.Y(n_3039)
);

BUFx12f_ASAP7_75t_L g3040 ( 
.A(n_2824),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2877),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2757),
.Y(n_3042)
);

OAI21x1_ASAP7_75t_L g3043 ( 
.A1(n_2764),
.A2(n_683),
.B(n_682),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2754),
.B(n_2861),
.Y(n_3044)
);

OAI21x1_ASAP7_75t_L g3045 ( 
.A1(n_2853),
.A2(n_685),
.B(n_684),
.Y(n_3045)
);

OAI21x1_ASAP7_75t_SL g3046 ( 
.A1(n_2835),
.A2(n_2901),
.B(n_2885),
.Y(n_3046)
);

CKINVDCx11_ASAP7_75t_R g3047 ( 
.A(n_2802),
.Y(n_3047)
);

BUFx2_ASAP7_75t_L g3048 ( 
.A(n_2788),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2896),
.B(n_686),
.Y(n_3049)
);

BUFx2_ASAP7_75t_L g3050 ( 
.A(n_2790),
.Y(n_3050)
);

BUFx2_ASAP7_75t_SL g3051 ( 
.A(n_2769),
.Y(n_3051)
);

OAI21x1_ASAP7_75t_L g3052 ( 
.A1(n_2819),
.A2(n_688),
.B(n_687),
.Y(n_3052)
);

AO31x2_ASAP7_75t_L g3053 ( 
.A1(n_2939),
.A2(n_899),
.A3(n_688),
.B(n_689),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2826),
.B(n_2913),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2965),
.A2(n_688),
.B1(n_689),
.B2(n_687),
.Y(n_3055)
);

OA21x2_ASAP7_75t_L g3056 ( 
.A1(n_2821),
.A2(n_690),
.B(n_689),
.Y(n_3056)
);

OAI21x1_ASAP7_75t_L g3057 ( 
.A1(n_2956),
.A2(n_691),
.B(n_690),
.Y(n_3057)
);

OA21x2_ASAP7_75t_L g3058 ( 
.A1(n_2813),
.A2(n_691),
.B(n_690),
.Y(n_3058)
);

INVx5_ASAP7_75t_L g3059 ( 
.A(n_2818),
.Y(n_3059)
);

OR2x6_ASAP7_75t_L g3060 ( 
.A(n_2900),
.B(n_692),
.Y(n_3060)
);

OAI21x1_ASAP7_75t_L g3061 ( 
.A1(n_2963),
.A2(n_694),
.B(n_693),
.Y(n_3061)
);

NOR2x1_ASAP7_75t_R g3062 ( 
.A(n_2892),
.B(n_693),
.Y(n_3062)
);

OAI21x1_ASAP7_75t_L g3063 ( 
.A1(n_2968),
.A2(n_695),
.B(n_694),
.Y(n_3063)
);

BUFx2_ASAP7_75t_SL g3064 ( 
.A(n_2811),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2855),
.B(n_694),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2803),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2806),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2809),
.Y(n_3068)
);

INVx3_ASAP7_75t_L g3069 ( 
.A(n_2836),
.Y(n_3069)
);

OA21x2_ASAP7_75t_L g3070 ( 
.A1(n_2777),
.A2(n_700),
.B(n_699),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2937),
.Y(n_3071)
);

OAI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2914),
.A2(n_701),
.B(n_699),
.Y(n_3072)
);

OAI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2884),
.A2(n_703),
.B(n_702),
.Y(n_3073)
);

OAI21x1_ASAP7_75t_L g3074 ( 
.A1(n_2857),
.A2(n_703),
.B(n_702),
.Y(n_3074)
);

OAI21x1_ASAP7_75t_L g3075 ( 
.A1(n_2879),
.A2(n_2880),
.B(n_2820),
.Y(n_3075)
);

OA21x2_ASAP7_75t_L g3076 ( 
.A1(n_2793),
.A2(n_705),
.B(n_704),
.Y(n_3076)
);

BUFx2_ASAP7_75t_L g3077 ( 
.A(n_2930),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2807),
.Y(n_3078)
);

INVx5_ASAP7_75t_L g3079 ( 
.A(n_2916),
.Y(n_3079)
);

OAI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2842),
.A2(n_708),
.B1(n_709),
.B2(n_707),
.Y(n_3080)
);

AOI21x1_ASAP7_75t_L g3081 ( 
.A1(n_2869),
.A2(n_710),
.B(n_709),
.Y(n_3081)
);

INVx6_ASAP7_75t_L g3082 ( 
.A(n_2916),
.Y(n_3082)
);

CKINVDCx6p67_ASAP7_75t_R g3083 ( 
.A(n_2798),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2888),
.Y(n_3084)
);

OAI221xp5_ASAP7_75t_L g3085 ( 
.A1(n_2864),
.A2(n_714),
.B1(n_715),
.B2(n_713),
.C(n_712),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2967),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2906),
.B(n_716),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2931),
.B(n_893),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2969),
.Y(n_3089)
);

AOI221xp5_ASAP7_75t_L g3090 ( 
.A1(n_2827),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2768),
.Y(n_3091)
);

OA21x2_ASAP7_75t_L g3092 ( 
.A1(n_2893),
.A2(n_719),
.B(n_717),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2789),
.Y(n_3093)
);

INVxp67_ASAP7_75t_L g3094 ( 
.A(n_2915),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2789),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2923),
.B(n_892),
.Y(n_3096)
);

OAI21x1_ASAP7_75t_L g3097 ( 
.A1(n_2792),
.A2(n_721),
.B(n_720),
.Y(n_3097)
);

INVx6_ASAP7_75t_L g3098 ( 
.A(n_2916),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2794),
.Y(n_3099)
);

OAI21x1_ASAP7_75t_L g3100 ( 
.A1(n_2795),
.A2(n_2828),
.B(n_2800),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2796),
.Y(n_3101)
);

OAI21x1_ASAP7_75t_L g3102 ( 
.A1(n_2770),
.A2(n_725),
.B(n_723),
.Y(n_3102)
);

BUFx2_ASAP7_75t_L g3103 ( 
.A(n_2829),
.Y(n_3103)
);

INVx6_ASAP7_75t_L g3104 ( 
.A(n_2959),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_2783),
.A2(n_730),
.B(n_729),
.Y(n_3105)
);

OAI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_2834),
.A2(n_731),
.B1(n_732),
.B2(n_730),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2784),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2784),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2837),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2837),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2829),
.Y(n_3111)
);

OA21x2_ASAP7_75t_L g3112 ( 
.A1(n_2903),
.A2(n_734),
.B(n_733),
.Y(n_3112)
);

OAI21x1_ASAP7_75t_L g3113 ( 
.A1(n_2933),
.A2(n_737),
.B(n_736),
.Y(n_3113)
);

INVx3_ASAP7_75t_L g3114 ( 
.A(n_2982),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2973),
.Y(n_3115)
);

AND2x4_ASAP7_75t_L g3116 ( 
.A(n_3000),
.B(n_2959),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_3091),
.A2(n_2852),
.B(n_2845),
.Y(n_3117)
);

AO31x2_ASAP7_75t_L g3118 ( 
.A1(n_3109),
.A2(n_2966),
.A3(n_2846),
.B(n_2928),
.Y(n_3118)
);

AO21x2_ASAP7_75t_L g3119 ( 
.A1(n_3110),
.A2(n_2911),
.B(n_2938),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2976),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_3041),
.B(n_2959),
.Y(n_3121)
);

OA21x2_ASAP7_75t_L g3122 ( 
.A1(n_3107),
.A2(n_3108),
.B(n_3078),
.Y(n_3122)
);

AOI21xp33_ASAP7_75t_L g3123 ( 
.A1(n_3001),
.A2(n_2952),
.B(n_2878),
.Y(n_3123)
);

BUFx3_ASAP7_75t_L g3124 ( 
.A(n_3021),
.Y(n_3124)
);

AOI21x1_ASAP7_75t_L g3125 ( 
.A1(n_3003),
.A2(n_2814),
.B(n_2771),
.Y(n_3125)
);

OR2x2_ASAP7_75t_L g3126 ( 
.A(n_2971),
.B(n_2822),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2980),
.Y(n_3127)
);

AOI21x1_ASAP7_75t_L g3128 ( 
.A1(n_3081),
.A2(n_2946),
.B(n_2850),
.Y(n_3128)
);

OAI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2979),
.A2(n_2780),
.B1(n_2844),
.B2(n_2941),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_3026),
.Y(n_3130)
);

AND3x1_ASAP7_75t_L g3131 ( 
.A(n_3069),
.B(n_3020),
.C(n_2987),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2981),
.Y(n_3132)
);

BUFx8_ASAP7_75t_L g3133 ( 
.A(n_3040),
.Y(n_3133)
);

INVx4_ASAP7_75t_L g3134 ( 
.A(n_3021),
.Y(n_3134)
);

BUFx10_ASAP7_75t_L g3135 ( 
.A(n_2991),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3006),
.B(n_2817),
.Y(n_3136)
);

AO31x2_ASAP7_75t_L g3137 ( 
.A1(n_3103),
.A2(n_2953),
.A3(n_2957),
.B(n_2945),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_2989),
.A2(n_2859),
.B1(n_2870),
.B2(n_2868),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2992),
.Y(n_3139)
);

AOI21x1_ASAP7_75t_L g3140 ( 
.A1(n_3031),
.A2(n_2831),
.B(n_2816),
.Y(n_3140)
);

INVxp67_ASAP7_75t_L g3141 ( 
.A(n_3064),
.Y(n_3141)
);

OA21x2_ASAP7_75t_L g3142 ( 
.A1(n_3093),
.A2(n_2935),
.B(n_2934),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2995),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_2975),
.B(n_2822),
.Y(n_3144)
);

OR2x6_ASAP7_75t_L g3145 ( 
.A(n_2994),
.B(n_2887),
.Y(n_3145)
);

OAI21x1_ASAP7_75t_L g3146 ( 
.A1(n_2986),
.A2(n_3034),
.B(n_3100),
.Y(n_3146)
);

AO21x2_ASAP7_75t_L g3147 ( 
.A1(n_3095),
.A2(n_2873),
.B(n_2875),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2998),
.Y(n_3148)
);

NAND2x1p5_ASAP7_75t_L g3149 ( 
.A(n_3079),
.B(n_2848),
.Y(n_3149)
);

OAI21x1_ASAP7_75t_L g3150 ( 
.A1(n_3075),
.A2(n_2823),
.B(n_2947),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2996),
.Y(n_3151)
);

AO21x2_ASAP7_75t_L g3152 ( 
.A1(n_3099),
.A2(n_2748),
.B(n_2750),
.Y(n_3152)
);

AO21x2_ASAP7_75t_L g3153 ( 
.A1(n_3101),
.A2(n_2926),
.B(n_2924),
.Y(n_3153)
);

HB1xp67_ASAP7_75t_L g3154 ( 
.A(n_3018),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2997),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2999),
.Y(n_3156)
);

OAI21x1_ASAP7_75t_L g3157 ( 
.A1(n_3005),
.A2(n_2904),
.B(n_2897),
.Y(n_3157)
);

AO31x2_ASAP7_75t_L g3158 ( 
.A1(n_3048),
.A2(n_2762),
.A3(n_2936),
.B(n_2927),
.Y(n_3158)
);

OAI21x1_ASAP7_75t_L g3159 ( 
.A1(n_2983),
.A2(n_2905),
.B(n_2960),
.Y(n_3159)
);

BUFx2_ASAP7_75t_L g3160 ( 
.A(n_2977),
.Y(n_3160)
);

AO31x2_ASAP7_75t_L g3161 ( 
.A1(n_3050),
.A2(n_2942),
.A3(n_2940),
.B(n_2950),
.Y(n_3161)
);

AOI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_3046),
.A2(n_2961),
.B1(n_2954),
.B2(n_2917),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_3029),
.B(n_2840),
.Y(n_3163)
);

AO31x2_ASAP7_75t_L g3164 ( 
.A1(n_3077),
.A2(n_2810),
.A3(n_2815),
.B(n_2962),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2984),
.B(n_2829),
.Y(n_3165)
);

NOR2x1_ASAP7_75t_SL g3166 ( 
.A(n_3079),
.B(n_2944),
.Y(n_3166)
);

CKINVDCx20_ASAP7_75t_R g3167 ( 
.A(n_3015),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2974),
.B(n_2747),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3014),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_3002),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3016),
.Y(n_3171)
);

NAND2x1p5_ASAP7_75t_L g3172 ( 
.A(n_3059),
.B(n_2970),
.Y(n_3172)
);

AO21x2_ASAP7_75t_L g3173 ( 
.A1(n_3072),
.A2(n_2922),
.B(n_2921),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_3036),
.Y(n_3174)
);

BUFx12f_ASAP7_75t_L g3175 ( 
.A(n_3010),
.Y(n_3175)
);

OR2x6_ASAP7_75t_L g3176 ( 
.A(n_3051),
.B(n_2943),
.Y(n_3176)
);

OAI21x1_ASAP7_75t_L g3177 ( 
.A1(n_3111),
.A2(n_2895),
.B(n_2912),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_3030),
.B(n_2993),
.Y(n_3178)
);

BUFx12f_ASAP7_75t_L g3179 ( 
.A(n_3028),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2972),
.A2(n_2881),
.B(n_2886),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_3012),
.A2(n_2881),
.B(n_2890),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3007),
.Y(n_3182)
);

AOI21x1_ASAP7_75t_L g3183 ( 
.A1(n_3060),
.A2(n_2866),
.B(n_2865),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2990),
.Y(n_3184)
);

INVxp33_ASAP7_75t_L g3185 ( 
.A(n_3047),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3042),
.Y(n_3186)
);

OA21x2_ASAP7_75t_L g3187 ( 
.A1(n_2988),
.A2(n_2773),
.B(n_2841),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_3066),
.B(n_2929),
.Y(n_3188)
);

AO21x1_ASAP7_75t_L g3189 ( 
.A1(n_3027),
.A2(n_2753),
.B(n_2756),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_3044),
.B(n_2841),
.Y(n_3190)
);

OR2x2_ASAP7_75t_L g3191 ( 
.A(n_3178),
.B(n_3184),
.Y(n_3191)
);

CKINVDCx6p67_ASAP7_75t_R g3192 ( 
.A(n_3124),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3115),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3122),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3120),
.Y(n_3195)
);

CKINVDCx5p33_ASAP7_75t_R g3196 ( 
.A(n_3175),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_3154),
.B(n_3054),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3127),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_3130),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3132),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_L g3201 ( 
.A1(n_3146),
.A2(n_2978),
.B(n_3011),
.Y(n_3201)
);

CKINVDCx6p67_ASAP7_75t_R g3202 ( 
.A(n_3134),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_3143),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_3148),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3139),
.Y(n_3205)
);

AND2x4_ASAP7_75t_L g3206 ( 
.A(n_3160),
.B(n_3071),
.Y(n_3206)
);

BUFx3_ASAP7_75t_L g3207 ( 
.A(n_3133),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_3170),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3165),
.B(n_3094),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3151),
.Y(n_3210)
);

OA21x2_ASAP7_75t_L g3211 ( 
.A1(n_3180),
.A2(n_3068),
.B(n_3067),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3182),
.Y(n_3212)
);

BUFx2_ASAP7_75t_L g3213 ( 
.A(n_3116),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3155),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_3121),
.Y(n_3215)
);

AO21x2_ASAP7_75t_L g3216 ( 
.A1(n_3123),
.A2(n_3181),
.B(n_3188),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_3156),
.Y(n_3217)
);

AND2x4_ASAP7_75t_L g3218 ( 
.A(n_3174),
.B(n_3077),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3186),
.B(n_3083),
.Y(n_3219)
);

AND2x4_ASAP7_75t_SL g3220 ( 
.A(n_3135),
.B(n_3039),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3169),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3171),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_3141),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3163),
.Y(n_3224)
);

OAI22xp5_ASAP7_75t_L g3225 ( 
.A1(n_3145),
.A2(n_3131),
.B1(n_3162),
.B2(n_3138),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3168),
.B(n_3084),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3163),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3126),
.Y(n_3228)
);

OR2x2_ASAP7_75t_L g3229 ( 
.A(n_3190),
.B(n_3037),
.Y(n_3229)
);

BUFx4f_ASAP7_75t_L g3230 ( 
.A(n_3114),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3144),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3153),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3152),
.Y(n_3233)
);

CKINVDCx6p67_ASAP7_75t_R g3234 ( 
.A(n_3179),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_SL g3235 ( 
.A(n_3185),
.B(n_3062),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3119),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3147),
.Y(n_3237)
);

HB1xp67_ASAP7_75t_L g3238 ( 
.A(n_3161),
.Y(n_3238)
);

INVx3_ASAP7_75t_L g3239 ( 
.A(n_3145),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3187),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3142),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3136),
.Y(n_3242)
);

AND2x4_ASAP7_75t_L g3243 ( 
.A(n_3166),
.B(n_3086),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3158),
.B(n_3089),
.Y(n_3244)
);

BUFx6f_ASAP7_75t_L g3245 ( 
.A(n_3149),
.Y(n_3245)
);

OR2x6_ASAP7_75t_L g3246 ( 
.A(n_3176),
.B(n_3082),
.Y(n_3246)
);

INVx2_ASAP7_75t_SL g3247 ( 
.A(n_3167),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3117),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_3202),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_L g3250 ( 
.A1(n_3225),
.A2(n_3129),
.B1(n_3189),
.B2(n_3173),
.Y(n_3250)
);

AND2x4_ASAP7_75t_L g3251 ( 
.A(n_3239),
.B(n_3150),
.Y(n_3251)
);

OAI22xp33_ASAP7_75t_L g3252 ( 
.A1(n_3246),
.A2(n_3172),
.B1(n_3008),
.B2(n_3085),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3231),
.B(n_3137),
.Y(n_3253)
);

OAI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3235),
.A2(n_3125),
.B(n_3183),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_3192),
.B(n_3038),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_3223),
.A2(n_3058),
.B1(n_3112),
.B2(n_3092),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3242),
.A2(n_3092),
.B1(n_3112),
.B2(n_3070),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3213),
.B(n_3215),
.Y(n_3258)
);

O2A1O1Ixp5_ASAP7_75t_SL g3259 ( 
.A1(n_3238),
.A2(n_3080),
.B(n_3106),
.C(n_3049),
.Y(n_3259)
);

AO21x2_ASAP7_75t_L g3260 ( 
.A1(n_3194),
.A2(n_3128),
.B(n_3140),
.Y(n_3260)
);

AOI22xp33_ASAP7_75t_L g3261 ( 
.A1(n_3244),
.A2(n_3056),
.B1(n_3004),
.B2(n_3023),
.Y(n_3261)
);

OAI22xp33_ASAP7_75t_L g3262 ( 
.A1(n_3215),
.A2(n_3098),
.B1(n_3104),
.B2(n_3082),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3209),
.B(n_3137),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3228),
.B(n_3118),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3240),
.Y(n_3265)
);

AOI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_3197),
.A2(n_3056),
.B1(n_3004),
.B2(n_3076),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3195),
.Y(n_3267)
);

OR2x6_ASAP7_75t_L g3268 ( 
.A(n_3207),
.B(n_3098),
.Y(n_3268)
);

CKINVDCx20_ASAP7_75t_R g3269 ( 
.A(n_3196),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3195),
.Y(n_3270)
);

AO21x2_ASAP7_75t_L g3271 ( 
.A1(n_3236),
.A2(n_3159),
.B(n_3157),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3217),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3226),
.A2(n_3065),
.B1(n_3087),
.B2(n_3088),
.Y(n_3273)
);

CKINVDCx6p67_ASAP7_75t_R g3274 ( 
.A(n_3234),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_3220),
.Y(n_3275)
);

INVx2_ASAP7_75t_L g3276 ( 
.A(n_3203),
.Y(n_3276)
);

AOI221xp5_ASAP7_75t_L g3277 ( 
.A1(n_3237),
.A2(n_3090),
.B1(n_3022),
.B2(n_3096),
.C(n_3055),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3204),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3212),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_3206),
.B(n_3164),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3193),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3224),
.Y(n_3282)
);

OAI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_3230),
.A2(n_3164),
.B1(n_3118),
.B2(n_3024),
.Y(n_3283)
);

INVx3_ASAP7_75t_L g3284 ( 
.A(n_3245),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_SL g3285 ( 
.A1(n_3211),
.A2(n_3177),
.B1(n_3035),
.B2(n_3009),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3219),
.A2(n_2985),
.B1(n_3043),
.B2(n_3073),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3218),
.A2(n_3052),
.B1(n_3025),
.B2(n_3019),
.Y(n_3287)
);

AOI221xp5_ASAP7_75t_L g3288 ( 
.A1(n_3232),
.A2(n_2955),
.B1(n_2951),
.B2(n_3053),
.C(n_3033),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_3218),
.A2(n_3113),
.B1(n_3013),
.B2(n_3032),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3227),
.B(n_3053),
.Y(n_3290)
);

OAI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3245),
.A2(n_2955),
.B1(n_3024),
.B2(n_3017),
.Y(n_3291)
);

AOI21xp33_ASAP7_75t_L g3292 ( 
.A1(n_3216),
.A2(n_3102),
.B(n_3097),
.Y(n_3292)
);

INVxp67_ASAP7_75t_L g3293 ( 
.A(n_3247),
.Y(n_3293)
);

OAI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_3243),
.A2(n_3017),
.B1(n_2929),
.B2(n_2882),
.Y(n_3294)
);

AOI221xp5_ASAP7_75t_L g3295 ( 
.A1(n_3232),
.A2(n_742),
.B1(n_743),
.B2(n_741),
.C(n_739),
.Y(n_3295)
);

OAI221xp5_ASAP7_75t_L g3296 ( 
.A1(n_3233),
.A2(n_2948),
.B1(n_2854),
.B2(n_2902),
.C(n_2882),
.Y(n_3296)
);

AOI222xp33_ASAP7_75t_L g3297 ( 
.A1(n_3233),
.A2(n_3105),
.B1(n_3045),
.B2(n_3057),
.C1(n_3063),
.C2(n_3061),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3198),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3200),
.Y(n_3299)
);

HB1xp67_ASAP7_75t_L g3300 ( 
.A(n_3258),
.Y(n_3300)
);

AND2x4_ASAP7_75t_L g3301 ( 
.A(n_3280),
.B(n_3241),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3250),
.A2(n_3191),
.B1(n_3243),
.B2(n_3229),
.Y(n_3302)
);

AND2x4_ASAP7_75t_L g3303 ( 
.A(n_3251),
.B(n_3201),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3282),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3267),
.Y(n_3305)
);

INVxp67_ASAP7_75t_L g3306 ( 
.A(n_3268),
.Y(n_3306)
);

OR2x2_ASAP7_75t_L g3307 ( 
.A(n_3264),
.B(n_3253),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3263),
.B(n_3199),
.Y(n_3308)
);

NOR2x1_ASAP7_75t_L g3309 ( 
.A(n_3268),
.B(n_3205),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_3265),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3270),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3251),
.B(n_3210),
.Y(n_3312)
);

AND2x2_ASAP7_75t_L g3313 ( 
.A(n_3284),
.B(n_3214),
.Y(n_3313)
);

BUFx6f_ASAP7_75t_SL g3314 ( 
.A(n_3274),
.Y(n_3314)
);

OR2x2_ASAP7_75t_L g3315 ( 
.A(n_3290),
.B(n_3208),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3272),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3279),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3281),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3276),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3298),
.Y(n_3320)
);

NOR2xp67_ASAP7_75t_L g3321 ( 
.A(n_3249),
.B(n_3248),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3299),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3278),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_L g3324 ( 
.A(n_3275),
.B(n_3221),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_3260),
.B(n_3222),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3293),
.B(n_3248),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3271),
.Y(n_3327)
);

AND2x4_ASAP7_75t_L g3328 ( 
.A(n_3254),
.B(n_3074),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3283),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3273),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3294),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3296),
.Y(n_3332)
);

INVx2_ASAP7_75t_SL g3333 ( 
.A(n_3255),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3285),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_3314),
.B(n_3269),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3306),
.B(n_3261),
.Y(n_3336)
);

OR2x2_ASAP7_75t_L g3337 ( 
.A(n_3331),
.B(n_3257),
.Y(n_3337)
);

NAND2x1p5_ASAP7_75t_L g3338 ( 
.A(n_3309),
.B(n_3262),
.Y(n_3338)
);

AND2x4_ASAP7_75t_L g3339 ( 
.A(n_3333),
.B(n_3286),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3300),
.B(n_3292),
.Y(n_3340)
);

OR2x2_ASAP7_75t_L g3341 ( 
.A(n_3331),
.B(n_3256),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_3312),
.B(n_3266),
.Y(n_3342)
);

AND2x4_ASAP7_75t_L g3343 ( 
.A(n_3329),
.B(n_3289),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3314),
.B(n_3252),
.Y(n_3344)
);

HB1xp67_ASAP7_75t_L g3345 ( 
.A(n_3304),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3330),
.B(n_3288),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3332),
.B(n_3291),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3326),
.B(n_3287),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3308),
.B(n_3297),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3301),
.B(n_3277),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3316),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3310),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3301),
.B(n_3259),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3313),
.B(n_3295),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_3317),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3305),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3311),
.Y(n_3357)
);

HB1xp67_ASAP7_75t_L g3358 ( 
.A(n_3325),
.Y(n_3358)
);

AND2x4_ASAP7_75t_SL g3359 ( 
.A(n_3324),
.B(n_742),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3319),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3318),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3318),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3303),
.B(n_37),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3334),
.B(n_37),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3320),
.Y(n_3365)
);

NOR2x1p5_ASAP7_75t_L g3366 ( 
.A(n_3328),
.B(n_744),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_3328),
.B(n_744),
.Y(n_3367)
);

NAND2x1p5_ASAP7_75t_L g3368 ( 
.A(n_3321),
.B(n_744),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3344),
.B(n_3302),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3338),
.B(n_3307),
.Y(n_3370)
);

AOI221xp5_ASAP7_75t_L g3371 ( 
.A1(n_3346),
.A2(n_3327),
.B1(n_3322),
.B2(n_3323),
.C(n_3315),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3345),
.Y(n_3372)
);

OAI21xp33_ASAP7_75t_L g3373 ( 
.A1(n_3347),
.A2(n_38),
.B(n_39),
.Y(n_3373)
);

OR2x2_ASAP7_75t_L g3374 ( 
.A(n_3337),
.B(n_3341),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3350),
.B(n_3336),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3366),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3363),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3339),
.B(n_40),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3355),
.Y(n_3379)
);

OR2x2_ASAP7_75t_L g3380 ( 
.A(n_3364),
.B(n_41),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3365),
.Y(n_3381)
);

OAI31xp33_ASAP7_75t_SL g3382 ( 
.A1(n_3367),
.A2(n_43),
.A3(n_41),
.B(n_42),
.Y(n_3382)
);

AND2x4_ASAP7_75t_SL g3383 ( 
.A(n_3335),
.B(n_42),
.Y(n_3383)
);

INVx3_ASAP7_75t_L g3384 ( 
.A(n_3368),
.Y(n_3384)
);

BUFx3_ASAP7_75t_L g3385 ( 
.A(n_3359),
.Y(n_3385)
);

INVx2_ASAP7_75t_SL g3386 ( 
.A(n_3366),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3354),
.B(n_43),
.Y(n_3387)
);

OAI31xp33_ASAP7_75t_L g3388 ( 
.A1(n_3343),
.A2(n_46),
.A3(n_44),
.B(n_45),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_SL g3389 ( 
.A(n_3353),
.B(n_46),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3375),
.B(n_3348),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3378),
.Y(n_3391)
);

AND2x2_ASAP7_75t_L g3392 ( 
.A(n_3370),
.B(n_3342),
.Y(n_3392)
);

INVx1_ASAP7_75t_SL g3393 ( 
.A(n_3383),
.Y(n_3393)
);

NAND3xp33_ASAP7_75t_L g3394 ( 
.A(n_3389),
.B(n_3358),
.C(n_3340),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_3384),
.B(n_3349),
.Y(n_3395)
);

INVx1_ASAP7_75t_SL g3396 ( 
.A(n_3385),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3374),
.B(n_3361),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3388),
.B(n_3362),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3372),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3379),
.B(n_3362),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3379),
.Y(n_3401)
);

OR2x2_ASAP7_75t_L g3402 ( 
.A(n_3387),
.B(n_3351),
.Y(n_3402)
);

AND2x4_ASAP7_75t_L g3403 ( 
.A(n_3386),
.B(n_3352),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3377),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3369),
.B(n_3360),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3381),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3380),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3396),
.B(n_3373),
.Y(n_3408)
);

NAND4xp25_ASAP7_75t_L g3409 ( 
.A(n_3394),
.B(n_3382),
.C(n_3376),
.D(n_3371),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3393),
.B(n_3395),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3403),
.Y(n_3411)
);

OR2x6_ASAP7_75t_L g3412 ( 
.A(n_3407),
.B(n_3356),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3391),
.Y(n_3413)
);

OR2x2_ASAP7_75t_L g3414 ( 
.A(n_3398),
.B(n_3357),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3405),
.B(n_46),
.Y(n_3415)
);

OR2x2_ASAP7_75t_L g3416 ( 
.A(n_3397),
.B(n_47),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_L g3417 ( 
.A(n_3392),
.B(n_48),
.Y(n_3417)
);

OAI322xp33_ASAP7_75t_L g3418 ( 
.A1(n_3399),
.A2(n_3397),
.A3(n_3390),
.B1(n_3404),
.B2(n_3394),
.C1(n_3401),
.C2(n_3402),
.Y(n_3418)
);

AND2x4_ASAP7_75t_L g3419 ( 
.A(n_3406),
.B(n_50),
.Y(n_3419)
);

INVxp67_ASAP7_75t_L g3420 ( 
.A(n_3400),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3400),
.Y(n_3421)
);

NOR2xp33_ASAP7_75t_L g3422 ( 
.A(n_3396),
.B(n_50),
.Y(n_3422)
);

OR2x2_ASAP7_75t_L g3423 ( 
.A(n_3416),
.B(n_51),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3410),
.B(n_51),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3422),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3411),
.Y(n_3426)
);

INVx1_ASAP7_75t_SL g3427 ( 
.A(n_3408),
.Y(n_3427)
);

AND2x4_ASAP7_75t_L g3428 ( 
.A(n_3419),
.B(n_55),
.Y(n_3428)
);

OAI21xp33_ASAP7_75t_L g3429 ( 
.A1(n_3409),
.A2(n_55),
.B(n_56),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3415),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3412),
.Y(n_3431)
);

INVxp67_ASAP7_75t_L g3432 ( 
.A(n_3417),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3413),
.B(n_57),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3414),
.Y(n_3434)
);

OAI31xp33_ASAP7_75t_L g3435 ( 
.A1(n_3429),
.A2(n_3421),
.A3(n_3420),
.B(n_3418),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3426),
.Y(n_3436)
);

AOI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3427),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3431),
.Y(n_3438)
);

OAI22xp33_ASAP7_75t_SL g3439 ( 
.A1(n_3430),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_3439)
);

NOR2x1_ASAP7_75t_L g3440 ( 
.A(n_3423),
.B(n_63),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3428),
.B(n_64),
.Y(n_3441)
);

AOI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3425),
.A2(n_3433),
.B1(n_3432),
.B2(n_3434),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3428),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3424),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3424),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3424),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3424),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3436),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3441),
.Y(n_3449)
);

AOI21xp33_ASAP7_75t_SL g3450 ( 
.A1(n_3435),
.A2(n_69),
.B(n_70),
.Y(n_3450)
);

AOI22xp33_ASAP7_75t_SL g3451 ( 
.A1(n_3438),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3443),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3437),
.Y(n_3453)
);

NAND2x1p5_ASAP7_75t_L g3454 ( 
.A(n_3440),
.B(n_746),
.Y(n_3454)
);

AO32x1_ASAP7_75t_L g3455 ( 
.A1(n_3444),
.A2(n_73),
.A3(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_3455)
);

OAI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3435),
.A2(n_71),
.B(n_72),
.Y(n_3456)
);

OAI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3442),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3439),
.Y(n_3458)
);

AOI211x1_ASAP7_75t_L g3459 ( 
.A1(n_3456),
.A2(n_3445),
.B(n_3447),
.C(n_3446),
.Y(n_3459)
);

AOI21xp33_ASAP7_75t_L g3460 ( 
.A1(n_3458),
.A2(n_80),
.B(n_81),
.Y(n_3460)
);

OA21x2_ASAP7_75t_L g3461 ( 
.A1(n_3448),
.A2(n_82),
.B(n_83),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3451),
.B(n_82),
.Y(n_3462)
);

AOI22xp5_ASAP7_75t_L g3463 ( 
.A1(n_3453),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3455),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3457),
.B(n_87),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_3455),
.A2(n_88),
.B(n_89),
.Y(n_3466)
);

NOR2xp67_ASAP7_75t_L g3467 ( 
.A(n_3452),
.B(n_89),
.Y(n_3467)
);

OAI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3454),
.A2(n_750),
.B1(n_748),
.B2(n_749),
.C(n_751),
.Y(n_3468)
);

AOI21xp33_ASAP7_75t_L g3469 ( 
.A1(n_3449),
.A2(n_752),
.B(n_753),
.Y(n_3469)
);

AOI211xp5_ASAP7_75t_L g3470 ( 
.A1(n_3450),
.A2(n_757),
.B(n_755),
.C(n_756),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3450),
.B(n_755),
.Y(n_3471)
);

NAND3xp33_ASAP7_75t_SL g3472 ( 
.A(n_3456),
.B(n_892),
.C(n_760),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3461),
.Y(n_3473)
);

NAND3xp33_ASAP7_75t_L g3474 ( 
.A(n_3470),
.B(n_763),
.C(n_764),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3472),
.A2(n_767),
.B1(n_765),
.B2(n_766),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3461),
.Y(n_3476)
);

AOI311xp33_ASAP7_75t_L g3477 ( 
.A1(n_3464),
.A2(n_891),
.A3(n_768),
.B(n_766),
.C(n_767),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_3471),
.B(n_769),
.Y(n_3478)
);

NAND4xp75_ASAP7_75t_L g3479 ( 
.A(n_3459),
.B(n_772),
.C(n_770),
.D(n_771),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3465),
.Y(n_3480)
);

OAI21xp33_ASAP7_75t_SL g3481 ( 
.A1(n_3467),
.A2(n_774),
.B(n_775),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3462),
.Y(n_3482)
);

AOI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3468),
.A2(n_779),
.B1(n_777),
.B2(n_778),
.Y(n_3483)
);

AOI31xp33_ASAP7_75t_L g3484 ( 
.A1(n_3469),
.A2(n_781),
.A3(n_779),
.B(n_780),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3463),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3466),
.B(n_782),
.Y(n_3486)
);

AOI21xp33_ASAP7_75t_SL g3487 ( 
.A1(n_3460),
.A2(n_783),
.B(n_784),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3473),
.B(n_784),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_R g3489 ( 
.A(n_3480),
.B(n_786),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3476),
.Y(n_3490)
);

O2A1O1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3486),
.A2(n_790),
.B(n_788),
.C(n_789),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_3477),
.B(n_791),
.Y(n_3492)
);

CKINVDCx6p67_ASAP7_75t_R g3493 ( 
.A(n_3482),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3479),
.Y(n_3494)
);

OAI32xp33_ASAP7_75t_L g3495 ( 
.A1(n_3481),
.A2(n_791),
.A3(n_792),
.B1(n_793),
.B2(n_794),
.Y(n_3495)
);

AOI211x1_ASAP7_75t_L g3496 ( 
.A1(n_3474),
.A2(n_795),
.B(n_793),
.C(n_794),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_L g3497 ( 
.A(n_3484),
.B(n_795),
.Y(n_3497)
);

AOI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_3478),
.A2(n_798),
.B1(n_796),
.B2(n_797),
.Y(n_3498)
);

OAI221xp5_ASAP7_75t_L g3499 ( 
.A1(n_3475),
.A2(n_796),
.B1(n_797),
.B2(n_798),
.C(n_799),
.Y(n_3499)
);

OAI21xp5_ASAP7_75t_SL g3500 ( 
.A1(n_3483),
.A2(n_797),
.B(n_799),
.Y(n_3500)
);

AOI21xp33_ASAP7_75t_SL g3501 ( 
.A1(n_3485),
.A2(n_800),
.B(n_801),
.Y(n_3501)
);

A2O1A1Ixp33_ASAP7_75t_L g3502 ( 
.A1(n_3487),
.A2(n_803),
.B(n_801),
.C(n_802),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3490),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_R g3504 ( 
.A(n_3494),
.B(n_890),
.Y(n_3504)
);

O2A1O1Ixp33_ASAP7_75t_L g3505 ( 
.A1(n_3492),
.A2(n_3502),
.B(n_3495),
.C(n_3488),
.Y(n_3505)
);

NOR4xp75_ASAP7_75t_L g3506 ( 
.A(n_3499),
.B(n_887),
.C(n_806),
.D(n_804),
.Y(n_3506)
);

NOR3xp33_ASAP7_75t_L g3507 ( 
.A(n_3491),
.B(n_805),
.C(n_806),
.Y(n_3507)
);

AOI221xp5_ASAP7_75t_L g3508 ( 
.A1(n_3501),
.A2(n_807),
.B1(n_808),
.B2(n_809),
.C(n_810),
.Y(n_3508)
);

NOR2xp33_ASAP7_75t_L g3509 ( 
.A(n_3497),
.B(n_809),
.Y(n_3509)
);

OR2x2_ASAP7_75t_L g3510 ( 
.A(n_3493),
.B(n_885),
.Y(n_3510)
);

A2O1A1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_3500),
.A2(n_814),
.B(n_812),
.C(n_813),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3503),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3510),
.Y(n_3513)
);

AOI22xp5_ASAP7_75t_L g3514 ( 
.A1(n_3509),
.A2(n_3498),
.B1(n_3496),
.B2(n_3489),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3511),
.B(n_815),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3506),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3505),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3504),
.Y(n_3518)
);

NOR2x1_ASAP7_75t_L g3519 ( 
.A(n_3507),
.B(n_817),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3508),
.B(n_819),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3512),
.Y(n_3521)
);

XNOR2x1_ASAP7_75t_L g3522 ( 
.A(n_3519),
.B(n_820),
.Y(n_3522)
);

AO22x1_ASAP7_75t_L g3523 ( 
.A1(n_3516),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.Y(n_3523)
);

OAI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_3517),
.A2(n_823),
.B(n_824),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3520),
.Y(n_3525)
);

INVxp67_ASAP7_75t_SL g3526 ( 
.A(n_3515),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3513),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3518),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3514),
.Y(n_3529)
);

AOI221x1_ASAP7_75t_L g3530 ( 
.A1(n_3529),
.A2(n_825),
.B1(n_826),
.B2(n_827),
.C(n_828),
.Y(n_3530)
);

AOI222xp33_ASAP7_75t_L g3531 ( 
.A1(n_3523),
.A2(n_827),
.B1(n_829),
.B2(n_830),
.C1(n_831),
.C2(n_832),
.Y(n_3531)
);

AOI22xp5_ASAP7_75t_L g3532 ( 
.A1(n_3527),
.A2(n_832),
.B1(n_829),
.B2(n_831),
.Y(n_3532)
);

AOI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3521),
.A2(n_832),
.B1(n_829),
.B2(n_831),
.Y(n_3533)
);

NAND4xp25_ASAP7_75t_L g3534 ( 
.A(n_3525),
.B(n_835),
.C(n_833),
.D(n_834),
.Y(n_3534)
);

NOR3x1_ASAP7_75t_L g3535 ( 
.A(n_3526),
.B(n_833),
.C(n_834),
.Y(n_3535)
);

NOR3xp33_ASAP7_75t_L g3536 ( 
.A(n_3534),
.B(n_3528),
.C(n_3524),
.Y(n_3536)
);

NOR2x1p5_ASAP7_75t_L g3537 ( 
.A(n_3535),
.B(n_3522),
.Y(n_3537)
);

OA22x2_ASAP7_75t_L g3538 ( 
.A1(n_3533),
.A2(n_836),
.B1(n_833),
.B2(n_835),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3531),
.B(n_835),
.Y(n_3539)
);

INVx3_ASAP7_75t_L g3540 ( 
.A(n_3538),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_3536),
.A2(n_3532),
.B1(n_3530),
.B2(n_838),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3539),
.Y(n_3542)
);

XNOR2x1_ASAP7_75t_L g3543 ( 
.A(n_3537),
.B(n_837),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3543),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3544),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_SL g3546 ( 
.A1(n_3545),
.A2(n_3542),
.B1(n_3540),
.B2(n_3541),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3545),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3546),
.Y(n_3548)
);

NAND2x1p5_ASAP7_75t_L g3549 ( 
.A(n_3548),
.B(n_3547),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3549),
.Y(n_3550)
);

AOI22xp33_ASAP7_75t_L g3551 ( 
.A1(n_3550),
.A2(n_839),
.B1(n_840),
.B2(n_841),
.Y(n_3551)
);

NOR2xp67_ASAP7_75t_L g3552 ( 
.A(n_3551),
.B(n_840),
.Y(n_3552)
);

NOR4xp25_ASAP7_75t_L g3553 ( 
.A(n_3552),
.B(n_842),
.C(n_843),
.D(n_844),
.Y(n_3553)
);

AOI211xp5_ASAP7_75t_L g3554 ( 
.A1(n_3553),
.A2(n_842),
.B(n_843),
.C(n_844),
.Y(n_3554)
);


endmodule