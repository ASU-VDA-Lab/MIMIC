module fake_jpeg_23268_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_102;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_4),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_32),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_50),
.B1(n_37),
.B2(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_22),
.B1(n_30),
.B2(n_23),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_25),
.B1(n_20),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_81),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_23),
.B1(n_62),
.B2(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_91),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_23),
.B1(n_29),
.B2(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_96),
.B1(n_41),
.B2(n_45),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_37),
.B1(n_41),
.B2(n_39),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_100),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_64),
.C(n_59),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_0),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_42),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_61),
.Y(n_130)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_45),
.A2(n_41),
.B1(n_24),
.B2(n_19),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_83),
.Y(n_138)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_94),
.B1(n_92),
.B2(n_95),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_45),
.B1(n_24),
.B2(n_18),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_123),
.B1(n_127),
.B2(n_105),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_43),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_89),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_9),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_81),
.B1(n_78),
.B2(n_75),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_32),
.B(n_35),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_33),
.B(n_32),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_56),
.B1(n_65),
.B2(n_18),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_74),
.B1(n_27),
.B2(n_34),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_96),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_86),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_136),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_135),
.A2(n_150),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_141),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_139),
.B(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_144),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_159),
.B(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_72),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_113),
.B(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_99),
.B1(n_79),
.B2(n_104),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_155),
.B1(n_162),
.B2(n_118),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_109),
.A2(n_79),
.B1(n_88),
.B2(n_99),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_71),
.B(n_36),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_36),
.C(n_103),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_27),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_8),
.B(n_14),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_125),
.B1(n_111),
.B2(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_36),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_165),
.B(n_174),
.Y(n_217)
);

OAI322xp33_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_114),
.A3(n_115),
.B1(n_126),
.B2(n_121),
.C1(n_130),
.C2(n_111),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_176),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_164),
.B1(n_160),
.B2(n_145),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_169),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_129),
.B(n_115),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_189),
.B(n_190),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_119),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_32),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_6),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_184),
.B1(n_155),
.B2(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_118),
.B1(n_116),
.B2(n_120),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_140),
.A2(n_116),
.B(n_120),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_142),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_8),
.B(n_14),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_190),
.B(n_166),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_162),
.A3(n_135),
.B1(n_157),
.B2(n_149),
.C1(n_163),
.C2(n_141),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_182),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_202),
.B(n_189),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_205),
.B(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_209),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_154),
.C(n_146),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_216),
.C(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_168),
.A2(n_138),
.B1(n_161),
.B2(n_139),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_213),
.B1(n_219),
.B2(n_195),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_139),
.B1(n_120),
.B2(n_102),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_102),
.C(n_1),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_166),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_170),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_229),
.B(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_227),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_232),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_170),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_238),
.C(n_239),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

NAND2x1_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_173),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_240),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_196),
.B1(n_201),
.B2(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_180),
.B1(n_183),
.B2(n_185),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_179),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_208),
.C(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_248),
.C(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_199),
.C(n_218),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_209),
.C(n_169),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_212),
.C(n_211),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_212),
.C(n_203),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_220),
.C(n_197),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_227),
.B1(n_241),
.B2(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_237),
.C(n_224),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_262),
.C(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_243),
.B(n_205),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_197),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_270),
.B(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_266),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_228),
.B1(n_231),
.B2(n_223),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_174),
.B1(n_187),
.B2(n_171),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_251),
.C(n_256),
.Y(n_279)
);

FAx1_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_230),
.CI(n_191),
.CON(n_270),
.SN(n_270)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_242),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_246),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_270),
.B1(n_9),
.B2(n_11),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_244),
.C(n_248),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_187),
.C(n_165),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_191),
.C(n_8),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_270),
.B(n_261),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_5),
.B(n_12),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_290),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_7),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_273),
.B1(n_278),
.B2(n_275),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_296),
.B(n_288),
.C(n_13),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_7),
.B(n_12),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_5),
.B(n_11),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_2),
.B(n_3),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_5),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_288),
.B(n_12),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_300),
.Y(n_302)
);

OAI321xp33_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_174),
.C(n_170),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_298),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_302),
.Y(n_304)
);


endmodule