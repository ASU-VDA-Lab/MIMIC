module fake_jpeg_18488_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_45),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_23),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_50),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_23),
.B(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_20),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_80),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_16),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_79),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx2_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_90),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_82),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_86),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_101),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_83),
.B1(n_66),
.B2(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_96),
.A2(n_104),
.B1(n_107),
.B2(n_115),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_61),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_44),
.B1(n_37),
.B2(n_42),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_44),
.B(n_37),
.C(n_42),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_87),
.B1(n_72),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_109),
.A2(n_110),
.B1(n_140),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_36),
.B1(n_39),
.B2(n_15),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_31),
.B1(n_39),
.B2(n_15),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_39),
.B1(n_43),
.B2(n_18),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_130),
.B1(n_138),
.B2(n_9),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_118),
.B(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_55),
.A2(n_39),
.B1(n_43),
.B2(n_4),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_46),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_47),
.B(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_8),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_54),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_57),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_62),
.B(n_6),
.C(n_7),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_48),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_147),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_69),
.B1(n_86),
.B2(n_80),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_148),
.B1(n_158),
.B2(n_159),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_100),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_91),
.B1(n_78),
.B2(n_77),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_56),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_157),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_92),
.A2(n_73),
.B1(n_67),
.B2(n_75),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_139),
.B1(n_111),
.B2(n_93),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_168),
.Y(n_199)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_65),
.B1(n_82),
.B2(n_9),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_113),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_165),
.B(n_167),
.Y(n_222)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_99),
.B(n_7),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_177),
.Y(n_194)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_187),
.B1(n_114),
.B2(n_122),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_7),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_130),
.B(n_121),
.Y(n_200)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_181),
.Y(n_206)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_10),
.B1(n_13),
.B2(n_97),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_134),
.B1(n_144),
.B2(n_98),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_13),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_191),
.Y(n_220)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_13),
.B(n_107),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_186),
.B1(n_180),
.B2(n_163),
.Y(n_227)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_135),
.B(n_105),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_103),
.B(n_139),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_134),
.B1(n_119),
.B2(n_103),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_193),
.A2(n_200),
.B1(n_210),
.B2(n_212),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_203),
.B(n_191),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_150),
.B1(n_178),
.B2(n_156),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_156),
.A2(n_114),
.B1(n_106),
.B2(n_137),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_153),
.A2(n_106),
.B1(n_114),
.B2(n_137),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_219),
.B1(n_224),
.B2(n_225),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_171),
.A2(n_98),
.B1(n_120),
.B2(n_95),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_153),
.A2(n_95),
.B1(n_121),
.B2(n_122),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_159),
.A2(n_102),
.B1(n_158),
.B2(n_161),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_227),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_233),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_160),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_154),
.B(n_184),
.C(n_160),
.D(n_185),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_246),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_239),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g237 ( 
.A(n_222),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_154),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_189),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_243),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_155),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_169),
.C(n_185),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_199),
.B1(n_224),
.B2(n_223),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_166),
.Y(n_248)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

AO22x1_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_191),
.B1(n_183),
.B2(n_182),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_170),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_251),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_162),
.C(n_179),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_254),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_176),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_181),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_188),
.C(n_152),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_188),
.B(n_192),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_223),
.B(n_206),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_196),
.B1(n_203),
.B2(n_192),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_232),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_196),
.B1(n_208),
.B2(n_219),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_277),
.B(n_278),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_202),
.B(n_201),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_236),
.A2(n_206),
.B1(n_201),
.B2(n_212),
.Y(n_278)
);

AO22x1_ASAP7_75t_SL g279 ( 
.A1(n_250),
.A2(n_217),
.B1(n_228),
.B2(n_198),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_284),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_259),
.B1(n_250),
.B2(n_234),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_258),
.B1(n_238),
.B2(n_249),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_288),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_292),
.B(n_300),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_301),
.B1(n_281),
.B2(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_239),
.B(n_235),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_303),
.B(n_304),
.Y(n_320)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_299),
.Y(n_322)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_252),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_253),
.B1(n_243),
.B2(n_257),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_306),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_233),
.B(n_244),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_207),
.B(n_254),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_246),
.C(n_231),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_308),
.C(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_255),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_307),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_197),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_217),
.C(n_230),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_311),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_221),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_276),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_230),
.C(n_188),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_292),
.C(n_309),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_221),
.B(n_232),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_265),
.B1(n_282),
.B2(n_285),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_316),
.A2(n_326),
.B1(n_335),
.B2(n_298),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_323),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_311),
.B1(n_295),
.B2(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_321),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_295),
.A2(n_283),
.B1(n_286),
.B2(n_281),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_262),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_329),
.C(n_314),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_286),
.B1(n_276),
.B2(n_289),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_294),
.B(n_297),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_275),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_334),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_230),
.C(n_271),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_310),
.A2(n_275),
.B1(n_287),
.B2(n_271),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_302),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_282),
.B1(n_205),
.B2(n_245),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_307),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_337),
.Y(n_345)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_354),
.C(n_355),
.Y(n_360)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_298),
.B(n_315),
.C(n_303),
.D(n_296),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_342),
.B(n_329),
.Y(n_361)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_346),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_308),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_353),
.B1(n_320),
.B2(n_330),
.Y(n_358)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_351),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_312),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_327),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_299),
.C(n_291),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_291),
.C(n_204),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_346),
.A2(n_316),
.B1(n_326),
.B2(n_332),
.Y(n_356)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_366),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_324),
.C(n_328),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_368),
.C(n_360),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_323),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_367),
.B(n_352),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_317),
.C(n_321),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_357),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_372),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_362),
.A2(n_347),
.B(n_343),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_330),
.B(n_369),
.Y(n_387)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_369),
.Y(n_376)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_365),
.C(n_340),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_360),
.B(n_345),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_366),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_339),
.B(n_349),
.Y(n_379)
);

AOI21x1_ASAP7_75t_SL g388 ( 
.A1(n_379),
.A2(n_380),
.B(n_350),
.Y(n_388)
);

NAND4xp25_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_342),
.C(n_338),
.D(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_381),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_348),
.B1(n_339),
.B2(n_363),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_382),
.B(n_383),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_368),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_380),
.B1(n_356),
.B2(n_376),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_385),
.C(n_377),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_388),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_392),
.B(n_394),
.Y(n_397)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_370),
.Y(n_393)
);

AOI31xp33_ASAP7_75t_L g399 ( 
.A1(n_393),
.A2(n_379),
.A3(n_387),
.B(n_383),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_367),
.C(n_364),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_389),
.A2(n_373),
.B(n_359),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_396),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_374),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_399),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_390),
.C(n_388),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_401),
.B(n_403),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_390),
.C(n_391),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_391),
.B(n_351),
.Y(n_405)
);

OAI321xp33_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_364),
.A3(n_319),
.B1(n_228),
.B2(n_204),
.C(n_266),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_404),
.B(n_211),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_408),
.A2(n_211),
.B(n_402),
.Y(n_409)
);


endmodule