module fake_jpeg_13266_n_492 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_492);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_492;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_58),
.B(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_61),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_1),
.C(n_2),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_65),
.A2(n_50),
.B(n_45),
.C(n_7),
.Y(n_171)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_49),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_67),
.B(n_108),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g124 ( 
.A(n_74),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_75),
.Y(n_184)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_77),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_2),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_40),
.B(n_3),
.CON(n_90),
.SN(n_90)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_48),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_41),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_97),
.Y(n_187)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g181 ( 
.A(n_99),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_27),
.B(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_113),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_46),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_27),
.B(n_4),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_4),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_117),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_33),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_118),
.B(n_119),
.Y(n_190)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_61),
.B(n_67),
.C(n_105),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_120),
.A2(n_176),
.B(n_118),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_29),
.B1(n_54),
.B2(n_51),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_125),
.A2(n_163),
.B1(n_165),
.B2(n_173),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_83),
.A2(n_29),
.B1(n_31),
.B2(n_81),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_134),
.A2(n_147),
.B(n_171),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_29),
.B1(n_53),
.B2(n_52),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_136),
.A2(n_137),
.B1(n_141),
.B2(n_144),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_75),
.A2(n_55),
.B1(n_53),
.B2(n_52),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_138),
.B(n_169),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_39),
.B1(n_54),
.B2(n_51),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_143),
.B(n_17),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_55),
.B1(n_38),
.B2(n_36),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_23),
.B1(n_45),
.B2(n_41),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_39),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_86),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_56),
.A2(n_21),
.B1(n_45),
.B2(n_50),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_74),
.A2(n_35),
.B(n_28),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_64),
.A2(n_45),
.B1(n_50),
.B2(n_7),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_172),
.A2(n_177),
.B1(n_176),
.B2(n_144),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_57),
.A2(n_45),
.B1(n_5),
.B2(n_7),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_69),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_62),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_108),
.B(n_8),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_73),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_180),
.A2(n_188),
.B1(n_173),
.B2(n_177),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_82),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_68),
.B(n_92),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_191),
.B(n_192),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_68),
.B(n_11),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_85),
.B(n_13),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_194),
.B(n_196),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_85),
.B(n_14),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_92),
.B(n_16),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_197),
.B(n_190),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_215),
.Y(n_270)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_181),
.Y(n_199)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_122),
.B(n_97),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_201),
.B(n_228),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_202),
.B(n_248),
.Y(n_267)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_120),
.A2(n_119),
.B1(n_87),
.B2(n_88),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_205),
.A2(n_213),
.B1(n_227),
.B2(n_234),
.Y(n_298)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_123),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_232),
.Y(n_277)
);

OR2x4_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_71),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_211),
.A2(n_216),
.B(n_225),
.Y(n_289)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_123),
.A2(n_89),
.B1(n_78),
.B2(n_118),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_155),
.A2(n_100),
.B1(n_93),
.B2(n_94),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_214),
.A2(n_235),
.B1(n_167),
.B2(n_158),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_140),
.B(n_97),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_218),
.B(n_261),
.C(n_225),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_133),
.B(n_17),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_222),
.Y(n_265)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx6_ASAP7_75t_SL g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_221),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_135),
.B(n_154),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_239),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_139),
.B(n_109),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_156),
.A2(n_99),
.B1(n_101),
.B2(n_104),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_121),
.B(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_114),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_233),
.Y(n_271)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_143),
.B(n_99),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_165),
.A2(n_160),
.B1(n_131),
.B2(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_142),
.B(n_139),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_244),
.Y(n_286)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_252),
.Y(n_281)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_243),
.A2(n_219),
.B1(n_222),
.B2(n_249),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_170),
.B(n_188),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_137),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_249),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_152),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_250),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_159),
.A2(n_182),
.B1(n_147),
.B2(n_150),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_151),
.B(n_179),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_124),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_124),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_251),
.B(n_254),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_187),
.B(n_153),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_136),
.B(n_129),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_257),
.Y(n_311)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_129),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_255),
.B(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_159),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_259),
.B(n_260),
.Y(n_293)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_153),
.B(n_145),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_146),
.C(n_162),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_134),
.B(n_146),
.C(n_162),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_263),
.A2(n_216),
.B(n_225),
.C(n_236),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_264),
.A2(n_266),
.B1(n_269),
.B2(n_304),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_167),
.B1(n_158),
.B2(n_195),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_208),
.A2(n_195),
.B1(n_184),
.B2(n_157),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_146),
.B(n_162),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_278),
.A2(n_280),
.B(n_303),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_309),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_240),
.A2(n_184),
.B(n_157),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_241),
.A2(n_175),
.B1(n_128),
.B2(n_174),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_285),
.B1(n_296),
.B2(n_307),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_241),
.A2(n_175),
.B1(n_128),
.B2(n_174),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_243),
.A2(n_244),
.B1(n_211),
.B2(n_253),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_218),
.B(n_200),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_310),
.C(n_309),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_233),
.B(n_216),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_214),
.A2(n_202),
.B1(n_231),
.B2(n_224),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_305),
.A2(n_221),
.B(n_199),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_258),
.A2(n_247),
.B1(n_255),
.B2(n_206),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_286),
.B1(n_289),
.B2(n_303),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_252),
.B(n_237),
.C(n_226),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_265),
.B(n_252),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_313),
.B(n_316),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_209),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_314),
.B(n_318),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_277),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_334),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_265),
.B(n_203),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_198),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_339),
.C(n_333),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_210),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_271),
.B(n_232),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_319),
.B(n_320),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_207),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_271),
.B(n_238),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_322),
.B(n_329),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_264),
.A2(n_257),
.B1(n_260),
.B2(n_220),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_325),
.A2(n_328),
.B1(n_332),
.B2(n_345),
.Y(n_376)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_277),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_338),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_304),
.A2(n_254),
.B1(n_217),
.B2(n_204),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_204),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_307),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_333),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_267),
.A2(n_280),
.B1(n_269),
.B2(n_296),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_336),
.A2(n_273),
.B1(n_301),
.B2(n_288),
.Y(n_357)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_281),
.B(n_310),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_286),
.C(n_290),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_287),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_295),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_342),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_268),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_344),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_281),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_267),
.A2(n_266),
.B1(n_298),
.B2(n_285),
.Y(n_345)
);

O2A1O1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_281),
.A2(n_292),
.B(n_305),
.C(n_288),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_347),
.A2(n_350),
.B(n_313),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_284),
.A2(n_312),
.B1(n_306),
.B2(n_282),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_272),
.B1(n_300),
.B2(n_297),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_282),
.B(n_312),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_349),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_306),
.B(n_279),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_330),
.A2(n_294),
.B1(n_273),
.B2(n_301),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_359),
.B1(n_374),
.B2(n_379),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_339),
.A2(n_275),
.B(n_283),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_321),
.B(n_350),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_330),
.A2(n_272),
.B1(n_300),
.B2(n_283),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_371),
.C(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_349),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_370),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_343),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_323),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_320),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_316),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_332),
.A2(n_276),
.B1(n_297),
.B2(n_345),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_378),
.A2(n_348),
.B1(n_315),
.B2(n_319),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_331),
.A2(n_276),
.B1(n_346),
.B2(n_336),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_338),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_383),
.C(n_402),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_338),
.C(n_346),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_384),
.B(n_389),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_356),
.Y(n_412)
);

AO32x1_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_380),
.A3(n_379),
.B1(n_364),
.B2(n_373),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_390),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_378),
.A2(n_318),
.B(n_347),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_368),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_347),
.B(n_344),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_405),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_324),
.B1(n_328),
.B2(n_325),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_376),
.B1(n_351),
.B2(n_352),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_322),
.Y(n_394)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_396),
.A2(n_404),
.B1(n_370),
.B2(n_357),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_351),
.B(n_340),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_398),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_372),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_403),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_367),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_376),
.A2(n_324),
.B1(n_341),
.B2(n_327),
.Y(n_404)
);

OAI32xp33_ASAP7_75t_L g405 ( 
.A1(n_364),
.A2(n_314),
.A3(n_327),
.B1(n_329),
.B2(n_338),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_366),
.C(n_367),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_412),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_410),
.B(n_422),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_371),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_420),
.C(n_401),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_414),
.A2(n_424),
.B1(n_393),
.B2(n_385),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_413),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_419),
.A2(n_425),
.B1(n_426),
.B2(n_396),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_367),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_372),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_404),
.A2(n_354),
.B1(n_369),
.B2(n_374),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_387),
.A2(n_369),
.B1(n_352),
.B2(n_377),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_387),
.A2(n_377),
.B1(n_361),
.B2(n_367),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_417),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_430),
.Y(n_443)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_417),
.Y(n_428)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_428),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_416),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_431),
.A2(n_435),
.B1(n_440),
.B2(n_414),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_407),
.B(n_384),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_432),
.B(n_442),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_385),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_436),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_426),
.A2(n_388),
.B1(n_400),
.B2(n_398),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_386),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_438),
.C(n_441),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_411),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_388),
.B1(n_391),
.B2(n_392),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_394),
.C(n_389),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_424),
.A2(n_381),
.B1(n_403),
.B2(n_399),
.Y(n_442)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_429),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_451),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_416),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_448),
.B(n_453),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g449 ( 
.A1(n_434),
.A2(n_408),
.B(n_409),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_415),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_437),
.B(n_408),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_335),
.Y(n_453)
);

AOI321xp33_ASAP7_75t_L g455 ( 
.A1(n_428),
.A2(n_421),
.A3(n_409),
.B1(n_433),
.B2(n_412),
.C(n_406),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_455),
.A2(n_440),
.B1(n_438),
.B2(n_435),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_460),
.Y(n_467)
);

HAxp5_ASAP7_75t_SL g457 ( 
.A(n_455),
.B(n_433),
.CON(n_457),
.SN(n_457)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_464),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_430),
.B1(n_427),
.B2(n_423),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_459),
.A2(n_446),
.B1(n_449),
.B2(n_443),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_436),
.Y(n_460)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_463),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_420),
.C(n_423),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_468),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_454),
.C(n_452),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_461),
.B(n_450),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_469),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_462),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_462),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_444),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_456),
.C(n_458),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_474),
.B(n_477),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_471),
.A2(n_461),
.B(n_458),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_479),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_463),
.C(n_459),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_483),
.C(n_474),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_469),
.C(n_472),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_484),
.B(n_485),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_465),
.C(n_381),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_465),
.C(n_395),
.Y(n_486)
);

OAI31xp33_ASAP7_75t_SL g488 ( 
.A1(n_486),
.A2(n_481),
.A3(n_405),
.B(n_335),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_355),
.B1(n_335),
.B2(n_353),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_355),
.B(n_487),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_335),
.B(n_353),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_326),
.Y(n_492)
);


endmodule