module fake_jpeg_31595_n_541 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_541);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_10),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_1),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_2),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_35),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_104),
.Y(n_126)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_100),
.Y(n_138)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_2),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_22),
.A2(n_23),
.B(n_49),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_106),
.Y(n_157)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_108),
.Y(n_143)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_110),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_28),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_45),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_35),
.B(n_2),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_34),
.B1(n_50),
.B2(n_49),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_161),
.B1(n_89),
.B2(n_100),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_50),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_82),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_54),
.B1(n_31),
.B2(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_124),
.A2(n_150),
.B1(n_171),
.B2(n_73),
.Y(n_200)
);

HAxp5_ASAP7_75t_SL g136 ( 
.A(n_80),
.B(n_54),
.CON(n_136),
.SN(n_136)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_141),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_31),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_40),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_147),
.B(n_154),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_98),
.A2(n_54),
.B1(n_36),
.B2(n_23),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_36),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_76),
.A2(n_22),
.B1(n_45),
.B2(n_5),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_99),
.B(n_3),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_55),
.C(n_56),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_57),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_169),
.B1(n_79),
.B2(n_96),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_61),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_20),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_8),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_63),
.A2(n_29),
.B1(n_20),
.B2(n_8),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_174),
.Y(n_266)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_181),
.Y(n_253)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_180),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_182),
.B(n_185),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_160),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_183),
.Y(n_274)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_187),
.A2(n_193),
.B1(n_226),
.B2(n_198),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_188),
.B(n_196),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_119),
.B(n_81),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_189),
.B(n_201),
.Y(n_263)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_192),
.Y(n_259)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_127),
.B(n_93),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_200),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_120),
.Y(n_207)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_209),
.B(n_210),
.Y(n_265)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_212),
.B1(n_217),
.B2(n_221),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_136),
.A2(n_104),
.B1(n_72),
.B2(n_67),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_157),
.A2(n_126),
.B(n_130),
.C(n_164),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_230),
.B(n_169),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_228),
.Y(n_238)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_218),
.Y(n_247)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_157),
.A2(n_66),
.B1(n_91),
.B2(n_88),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_117),
.A2(n_88),
.B1(n_29),
.B2(n_20),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_171),
.A2(n_29),
.B1(n_7),
.B2(n_8),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_130),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_152),
.B1(n_111),
.B2(n_112),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_170),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_240),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_117),
.B1(n_121),
.B2(n_112),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_234),
.A2(n_193),
.B1(n_212),
.B2(n_220),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_L g303 ( 
.A(n_239),
.B(n_177),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_114),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_196),
.B(n_135),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_267),
.Y(n_298)
);

AOI32xp33_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_111),
.A3(n_137),
.B1(n_158),
.B2(n_144),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_224),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_135),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_165),
.B1(n_162),
.B2(n_159),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_229),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_277),
.Y(n_323)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_225),
.B1(n_200),
.B2(n_202),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_284),
.B1(n_295),
.B2(n_308),
.Y(n_316)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_202),
.C(n_188),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_241),
.C(n_247),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_283),
.A2(n_301),
.B1(n_237),
.B2(n_242),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_225),
.B1(n_161),
.B2(n_162),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_261),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_289),
.Y(n_342)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_255),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_194),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_238),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g343 ( 
.A1(n_292),
.A2(n_303),
.B(n_191),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_307),
.B1(n_268),
.B2(n_242),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_258),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_296),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_139),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_207),
.B(n_118),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_300),
.A2(n_269),
.B(n_209),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_270),
.A2(n_199),
.B1(n_217),
.B2(n_205),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_302),
.B(n_304),
.Y(n_319)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_231),
.A2(n_178),
.B(n_221),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_241),
.B(n_254),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_175),
.B1(n_184),
.B2(n_139),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_245),
.A2(n_236),
.B1(n_259),
.B2(n_238),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_256),
.B1(n_250),
.B2(n_248),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_253),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_310),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_313),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_254),
.C(n_247),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_320),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_331),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_273),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_235),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_294),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_232),
.B1(n_208),
.B2(n_174),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_326),
.A2(n_336),
.B1(n_288),
.B2(n_289),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_232),
.B1(n_268),
.B2(n_250),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_329),
.B1(n_337),
.B2(n_277),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_280),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_282),
.A2(n_233),
.B1(n_243),
.B2(n_183),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_233),
.B1(n_243),
.B2(n_269),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_301),
.A2(n_211),
.B1(n_266),
.B2(n_237),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_SL g353 ( 
.A(n_339),
.B(n_343),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_300),
.A2(n_256),
.B(n_235),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_341),
.A2(n_306),
.B(n_297),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_314),
.B(n_310),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_344),
.B(n_349),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_345),
.A2(n_346),
.B(n_367),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_298),
.B(n_294),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_314),
.B(n_275),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_323),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_350),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_323),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_351),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_334),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_368),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_356),
.A2(n_361),
.B1(n_331),
.B2(n_340),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_369),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_373),
.B1(n_327),
.B2(n_337),
.Y(n_391)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_362),
.Y(n_403)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_363),
.Y(n_377)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_287),
.B(n_276),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_321),
.B(n_313),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_297),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_304),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_341),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_286),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_372),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_316),
.A2(n_278),
.B1(n_285),
.B2(n_266),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_330),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_330),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_361),
.A2(n_316),
.B1(n_336),
.B2(n_326),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_381),
.A2(n_394),
.B1(n_407),
.B2(n_358),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_312),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_392),
.C(n_393),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_395),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_355),
.A2(n_309),
.B1(n_340),
.B2(n_322),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_384),
.A2(n_352),
.B(n_371),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_401),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_329),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_325),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_338),
.C(n_335),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_338),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_366),
.Y(n_429)
);

XNOR2x2_ASAP7_75t_SL g399 ( 
.A(n_357),
.B(n_273),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_352),
.A2(n_333),
.B(n_322),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_400),
.A2(n_401),
.B(n_404),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_373),
.A2(n_322),
.B1(n_333),
.B2(n_302),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_350),
.B(n_305),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_362),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_346),
.A2(n_299),
.B1(n_246),
.B2(n_216),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_387),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_408),
.Y(n_447)
);

BUFx12_ASAP7_75t_L g410 ( 
.A(n_400),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_365),
.Y(n_414)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_415),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_364),
.Y(n_416)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_388),
.A2(n_355),
.B1(n_353),
.B2(n_367),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_407),
.B1(n_404),
.B2(n_383),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_419),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_396),
.A2(n_353),
.B(n_367),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_377),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_422),
.A2(n_423),
.B1(n_425),
.B2(n_426),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_389),
.Y(n_423)
);

INVx13_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_380),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_345),
.B(n_369),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_427),
.A2(n_430),
.B(n_432),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_431),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_372),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_363),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_377),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_381),
.A2(n_375),
.B1(n_360),
.B2(n_359),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_180),
.B(n_264),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_391),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_395),
.C(n_392),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_448),
.C(n_449),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_451),
.B1(n_452),
.B2(n_459),
.Y(n_478)
);

FAx1_ASAP7_75t_SL g444 ( 
.A(n_416),
.B(n_393),
.CI(n_397),
.CON(n_444),
.SN(n_444)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_456),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_415),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_382),
.C(n_406),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_406),
.C(n_385),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_376),
.C(n_390),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_414),
.C(n_433),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_423),
.A2(n_376),
.B1(n_378),
.B2(n_403),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_417),
.A2(n_408),
.B1(n_411),
.B2(n_428),
.Y(n_452)
);

FAx1_ASAP7_75t_SL g456 ( 
.A(n_412),
.B(n_251),
.CI(n_264),
.CON(n_456),
.SN(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_251),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_443),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_411),
.A2(n_246),
.B1(n_206),
.B2(n_11),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_441),
.A2(n_421),
.B1(n_422),
.B2(n_418),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_460),
.A2(n_440),
.B1(n_458),
.B2(n_419),
.Y(n_482)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_426),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_465),
.Y(n_481)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_464),
.Y(n_487)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_468),
.C(n_472),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_431),
.C(n_427),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_471),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_456),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_476),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_438),
.C(n_443),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_474),
.Y(n_494)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_452),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_475),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_489),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_445),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_488),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_485),
.Y(n_508)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_483),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_457),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_446),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_421),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_453),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_425),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_464),
.A2(n_447),
.B1(n_421),
.B2(n_410),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_493),
.A2(n_419),
.B1(n_409),
.B2(n_435),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_496),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_466),
.C(n_471),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_499),
.C(n_484),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_491),
.A2(n_466),
.B(n_420),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_478),
.C(n_444),
.Y(n_499)
);

FAx1_ASAP7_75t_SL g501 ( 
.A(n_481),
.B(n_430),
.CI(n_436),
.CON(n_501),
.SN(n_501)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_501),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_490),
.A2(n_409),
.B1(n_434),
.B2(n_410),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_506),
.B1(n_492),
.B2(n_487),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_425),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_507),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_480),
.A2(n_410),
.B1(n_444),
.B2(n_432),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_494),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_509),
.A2(n_510),
.B1(n_9),
.B2(n_12),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_493),
.A2(n_244),
.B1(n_10),
.B2(n_11),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_513),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_484),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_515),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_504),
.A2(n_485),
.B1(n_244),
.B2(n_15),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_516),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_506),
.A2(n_244),
.B(n_14),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_518),
.A2(n_499),
.B(n_507),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_13),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_508),
.C(n_500),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_16),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_522),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_525),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_497),
.C(n_15),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_517),
.C(n_527),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_518),
.B(n_521),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_528),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_531),
.B(n_523),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_534),
.B(n_535),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_SL g535 ( 
.A(n_530),
.B(n_520),
.C(n_511),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_536),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_537),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_532),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_SL g540 ( 
.A1(n_539),
.A2(n_514),
.B(n_519),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_16),
.B(n_498),
.Y(n_541)
);


endmodule