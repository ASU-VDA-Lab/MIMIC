module fake_jpeg_6640_n_281 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_38),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_23),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_34),
.Y(n_102)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_62),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_66),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_22),
.B1(n_40),
.B2(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_72),
.A2(n_86),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_22),
.B1(n_33),
.B2(n_39),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_84),
.B1(n_25),
.B2(n_21),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_33),
.C(n_39),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_88),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_83),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_17),
.B(n_3),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_106),
.B(n_17),
.C(n_5),
.Y(n_123)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_18),
.B1(n_36),
.B2(n_35),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_31),
.B1(n_38),
.B2(n_36),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_89),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_44),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_37),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_17),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_53),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_107),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_95),
.B1(n_101),
.B2(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_131),
.B1(n_134),
.B2(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_118),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_117),
.A2(n_142),
.B1(n_116),
.B2(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_126),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_123),
.B1(n_129),
.B2(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_131),
.Y(n_173)
);

OAI22x1_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_127),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_4),
.B(n_6),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_132),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_83),
.B1(n_99),
.B2(n_70),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_82),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_95),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_77),
.B(n_8),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_104),
.B(n_122),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_9),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_117),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_152),
.B1(n_154),
.B2(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_153),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_79),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_141),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_90),
.B1(n_74),
.B2(n_105),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_90),
.B1(n_107),
.B2(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_165),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_71),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_160),
.B(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_103),
.B1(n_94),
.B2(n_76),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_162),
.B1(n_168),
.B2(n_127),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_104),
.B1(n_69),
.B2(n_13),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_69),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_118),
.B(n_137),
.CI(n_108),
.CON(n_165),
.SN(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_137),
.B1(n_123),
.B2(n_136),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_126),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_194),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_119),
.B(n_139),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_195),
.B(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_200),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_133),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_132),
.B1(n_128),
.B2(n_127),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_109),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_144),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_131),
.B1(n_134),
.B2(n_116),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_168),
.C(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_190),
.C(n_199),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_145),
.B1(n_148),
.B2(n_172),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_206),
.B1(n_188),
.B2(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_172),
.B1(n_147),
.B2(n_153),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_181),
.B(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_214),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_157),
.B(n_162),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_219),
.B(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_175),
.A2(n_150),
.B(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_204),
.C(n_218),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_234),
.B(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_197),
.C(n_198),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_230),
.C(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_232),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_193),
.B1(n_200),
.B2(n_178),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_210),
.C(n_216),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_178),
.B1(n_183),
.B2(n_176),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_226),
.B(n_220),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_213),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_189),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_218),
.B(n_221),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_180),
.C(n_219),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_247),
.B(n_203),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_209),
.C(n_207),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_209),
.C(n_207),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_215),
.B(n_238),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_233),
.B(n_220),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_236),
.B(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_243),
.B1(n_229),
.B2(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_237),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_254),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_260),
.B(n_217),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_224),
.Y(n_265)
);

OAI211xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_242),
.B(n_259),
.C(n_267),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_251),
.B1(n_222),
.B2(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_266),
.B1(n_261),
.B2(n_265),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.Y(n_271)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_212),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_259),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_268),
.B(n_263),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_266),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_271),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_277),
.A2(n_278),
.B(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_276),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_275),
.Y(n_281)
);


endmodule