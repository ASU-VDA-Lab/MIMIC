module fake_ibex_899_n_3152 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3152);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3152;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2846;
wire n_2685;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_2723;
wire n_1616;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2585;
wire n_2220;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_768;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_3104;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_1488;
wire n_849;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2148;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2961;
wire n_2996;
wire n_2704;
wire n_2770;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_683;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_219),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_242),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_93),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_277),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_591),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_118),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_34),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_537),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_604),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_221),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_239),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_57),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_274),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_401),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_410),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_431),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_64),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_185),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_69),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_530),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_267),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_296),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_391),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_251),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_153),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_130),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_91),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_340),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_7),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_92),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_96),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_96),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_337),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_177),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_39),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_433),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_80),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_373),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_259),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_339),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_68),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_62),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_192),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_540),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_314),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_216),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_119),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_404),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_344),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_603),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_566),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_319),
.Y(n_660)
);

CKINVDCx14_ASAP7_75t_R g661 ( 
.A(n_536),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_167),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_492),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_567),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_342),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_506),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_255),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_222),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_6),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_598),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_57),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_90),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_491),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_549),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_237),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_436),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_181),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_399),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_504),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_480),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_485),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_232),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_40),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_551),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_568),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_495),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_453),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_547),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_4),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_157),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_394),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_556),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_356),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_358),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_387),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_332),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_33),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_440),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_534),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_462),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_484),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_468),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_571),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_3),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_249),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_162),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_430),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_97),
.B(n_157),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_517),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_461),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_97),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_392),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_217),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_518),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_526),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_53),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_102),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_353),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_295),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_563),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_133),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_487),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_532),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_10),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_140),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_130),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_387),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_581),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_91),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_192),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_449),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_273),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_590),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_469),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_496),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_413),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_318),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_499),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_87),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_481),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_137),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_510),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_488),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_152),
.Y(n_745)
);

BUFx2_ASAP7_75t_SL g746 ( 
.A(n_15),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_369),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_76),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_423),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_502),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_278),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_327),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_281),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_538),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_323),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_336),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_391),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_334),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_490),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_399),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_217),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_412),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_543),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_521),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_225),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_298),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_80),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_561),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_489),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_284),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_106),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_535),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_122),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_364),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_13),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_493),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_427),
.B(n_560),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_40),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_334),
.Y(n_779)
);

CKINVDCx14_ASAP7_75t_R g780 ( 
.A(n_397),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_586),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_56),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_141),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_444),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_100),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_170),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_358),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_443),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_204),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_524),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_383),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_425),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_113),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_115),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_459),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_68),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_113),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_1),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_486),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_354),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_36),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_515),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_327),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_357),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_280),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_270),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_450),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_114),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_441),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_463),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_109),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_120),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_328),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_262),
.Y(n_814)
);

BUFx10_ASAP7_75t_L g815 ( 
.A(n_291),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_122),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_595),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_44),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_267),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_305),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_197),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_58),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_188),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_79),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_201),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_70),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_509),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_225),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_174),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_180),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_92),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_305),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_185),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_67),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_308),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_82),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_352),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_458),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_542),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_447),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_72),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_264),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_364),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_268),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_85),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_248),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_3),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_550),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_193),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_376),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_501),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_254),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_12),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_541),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_600),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_37),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_131),
.Y(n_857)
);

BUFx10_ASAP7_75t_L g858 ( 
.A(n_149),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_351),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_211),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_400),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_88),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_478),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_572),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_297),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_432),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_257),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_580),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_152),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_520),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_89),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_215),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_18),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_331),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_308),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_148),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_513),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_466),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_287),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_454),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_607),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_389),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_245),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_163),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_465),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_188),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_451),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_55),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_589),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_564),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_467),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_240),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_426),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_511),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_103),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_577),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_143),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_383),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_309),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_414),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_531),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_328),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_148),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_585),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_392),
.Y(n_905)
);

INVx4_ASAP7_75t_R g906 ( 
.A(n_187),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_318),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_232),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_66),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_177),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_322),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_38),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_405),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_39),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_220),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_592),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_199),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_161),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_601),
.Y(n_919)
);

BUFx5_ASAP7_75t_L g920 ( 
.A(n_47),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_324),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_546),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_311),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_52),
.Y(n_924)
);

INVx4_ASAP7_75t_R g925 ( 
.A(n_374),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_151),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_275),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_396),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_278),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_10),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_359),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_584),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_338),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_108),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_448),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_428),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_45),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_253),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_516),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_346),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_120),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_602),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_325),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_544),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_174),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_319),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_311),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_229),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_429),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_36),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_236),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_61),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_479),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_299),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_482),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_165),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_72),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_271),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_250),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_241),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_361),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_452),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_295),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_525),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_261),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_155),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_71),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_539),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_271),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_406),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_32),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_69),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_762),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_624),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_679),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_612),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_708),
.B(n_870),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_658),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_741),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_889),
.B(n_0),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_658),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_920),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_658),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_624),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_780),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_624),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_920),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_780),
.B(n_0),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_920),
.Y(n_989)
);

INVx5_ASAP7_75t_L g990 ( 
.A(n_658),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_612),
.B(n_621),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_741),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_942),
.B(n_1),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_644),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_679),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_795),
.Y(n_996)
);

BUFx8_ASAP7_75t_SL g997 ( 
.A(n_625),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_920),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_631),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_621),
.B(n_2),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_920),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_668),
.B(n_2),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_758),
.B(n_4),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_672),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_614),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_758),
.B(n_5),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_794),
.B(n_5),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_672),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_679),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_803),
.B(n_6),
.Y(n_1010)
);

BUFx8_ASAP7_75t_L g1011 ( 
.A(n_961),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_613),
.Y(n_1012)
);

BUFx12f_ASAP7_75t_L g1013 ( 
.A(n_697),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_920),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_795),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_697),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_644),
.B(n_7),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_971),
.B(n_8),
.Y(n_1018)
);

AOI22x1_ASAP7_75t_SL g1019 ( 
.A1(n_625),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_826),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_917),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_917),
.B(n_826),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_853),
.Y(n_1023)
);

OAI22x1_ASAP7_75t_SL g1024 ( 
.A1(n_692),
.A2(n_13),
.B1(n_9),
.B2(n_12),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_821),
.B(n_14),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_614),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_614),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_853),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_947),
.B(n_14),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_739),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_701),
.A2(n_407),
.B(n_403),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_614),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_617),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_701),
.A2(n_409),
.B(n_408),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_671),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_R g1036 ( 
.A1(n_692),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_962),
.B(n_411),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_636),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_825),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_697),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_947),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_671),
.B(n_19),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_743),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_636),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_739),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_636),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_609),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_739),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_646),
.B(n_20),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_636),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_739),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_775),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_648),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_739),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_646),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_628),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_648),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_650),
.B(n_21),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_711),
.A2(n_416),
.B(n_415),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_743),
.B(n_21),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_648),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_650),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_815),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_815),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_648),
.Y(n_1065)
);

BUFx8_ASAP7_75t_L g1066 ( 
.A(n_788),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_824),
.B(n_835),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_962),
.B(n_417),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_788),
.B(n_22),
.Y(n_1069)
);

BUFx8_ASAP7_75t_SL g1070 ( 
.A(n_775),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_801),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_609),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_841),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_841),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_815),
.Y(n_1075)
);

INVxp33_ASAP7_75t_SL g1076 ( 
.A(n_639),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_850),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_801),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_801),
.Y(n_1079)
);

AOI22x1_ASAP7_75t_SL g1080 ( 
.A1(n_793),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_739),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_711),
.A2(n_419),
.B(n_418),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_938),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_639),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_850),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_724),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_801),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_874),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1006),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_1047),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1020),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_1076),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_978),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_985),
.B(n_661),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_L g1095 ( 
.A(n_974),
.B(n_984),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_1076),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1007),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_978),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_985),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_977),
.B(n_894),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_994),
.B(n_922),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_974),
.B(n_640),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1007),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_997),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_978),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_997),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_1052),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1052),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_1070),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_1070),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_974),
.B(n_640),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_995),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_979),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_975),
.B(n_610),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1013),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_981),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1072),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_1084),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1016),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1064),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1075),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_991),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_1011),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_975),
.B(n_661),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1077),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1085),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1011),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_991),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_999),
.Y(n_1129)
);

AND3x2_ASAP7_75t_L g1130 ( 
.A(n_999),
.B(n_911),
.C(n_778),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1049),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1012),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_R g1133 ( 
.A(n_1025),
.B(n_641),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1049),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1058),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_973),
.B(n_641),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1033),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1056),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1058),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1056),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1066),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_988),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_1009),
.B(n_659),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1023),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1066),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_974),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_1004),
.Y(n_1147)
);

AND3x2_ASAP7_75t_L g1148 ( 
.A(n_1036),
.B(n_787),
.C(n_760),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1004),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_979),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_984),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_984),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1008),
.B(n_858),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1008),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1028),
.B(n_858),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1023),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1028),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_986),
.B(n_1041),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

NOR2xp67_ASAP7_75t_L g1160 ( 
.A(n_986),
.B(n_922),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1009),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1040),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1040),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_1022),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1022),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1063),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1041),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1029),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1019),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1037),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1080),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_996),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1002),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1024),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1010),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_994),
.B(n_964),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1037),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1029),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_R g1179 ( 
.A(n_1018),
.B(n_642),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_976),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_980),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1039),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1030),
.A2(n_790),
.B(n_724),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1039),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_989),
.A2(n_866),
.B(n_790),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1021),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1015),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1067),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_993),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_993),
.Y(n_1190)
);

AND2x6_ASAP7_75t_L g1191 ( 
.A(n_1017),
.B(n_866),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_R g1192 ( 
.A(n_1037),
.B(n_659),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1017),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1069),
.Y(n_1194)
);

CKINVDCx16_ASAP7_75t_R g1195 ( 
.A(n_1037),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1069),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_994),
.B(n_964),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1067),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1042),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1000),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_982),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1042),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1060),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_987),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1000),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1060),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_L g1207 ( 
.A(n_1035),
.B(n_813),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1003),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1035),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1035),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_R g1211 ( 
.A(n_1037),
.B(n_664),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1086),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1035),
.B(n_643),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1043),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1043),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1055),
.B(n_858),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1043),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1043),
.B(n_623),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1062),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_998),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_R g1221 ( 
.A(n_1068),
.B(n_664),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_R g1222 ( 
.A(n_1068),
.B(n_693),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1073),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1074),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1083),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1068),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1068),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1068),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1001),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1045),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_R g1231 ( 
.A(n_1059),
.B(n_643),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_998),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1014),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1014),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1059),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1048),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1048),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1051),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1051),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1054),
.A2(n_647),
.B1(n_649),
.B2(n_645),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1081),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1031),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_990),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_990),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_990),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1005),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1005),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1005),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_R g1249 ( 
.A(n_1026),
.B(n_693),
.Y(n_1249)
);

NAND2xp33_ASAP7_75t_R g1250 ( 
.A(n_1034),
.B(n_645),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1026),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1082),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1026),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1027),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1027),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1027),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1032),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1032),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1032),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1038),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1038),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1038),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_981),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1044),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1044),
.B(n_647),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1044),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1046),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1046),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1046),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1050),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1050),
.Y(n_1271)
);

NOR2xp67_ASAP7_75t_L g1272 ( 
.A(n_1050),
.B(n_652),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1053),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1053),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1208),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1212),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1205),
.B(n_916),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1165),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1170),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1200),
.A2(n_936),
.B1(n_735),
.B2(n_651),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1165),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1144),
.B(n_663),
.Y(n_1282)
);

NAND2xp33_ASAP7_75t_L g1283 ( 
.A(n_1226),
.B(n_675),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1199),
.B(n_677),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1202),
.B(n_682),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1216),
.B(n_709),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_L g1287 ( 
.A(n_1217),
.B(n_420),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1149),
.A2(n_615),
.B1(n_622),
.B2(n_611),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1203),
.B(n_685),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1206),
.B(n_686),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1156),
.B(n_687),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1150),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1147),
.B(n_688),
.Y(n_1293)
);

XOR2xp5_ASAP7_75t_L g1294 ( 
.A(n_1123),
.B(n_796),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1181),
.B(n_699),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1179),
.B(n_653),
.C(n_651),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1122),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1159),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1122),
.B(n_935),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1195),
.B(n_700),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1153),
.B(n_703),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1128),
.B(n_970),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1180),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_L g1304 ( 
.A(n_1227),
.B(n_715),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1155),
.B(n_1158),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_L g1306 ( 
.A(n_1228),
.B(n_716),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1154),
.A2(n_630),
.B1(n_632),
.B2(n_627),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1100),
.B(n_1132),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1167),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1172),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1137),
.B(n_749),
.Y(n_1311)
);

BUFx5_ASAP7_75t_L g1312 ( 
.A(n_1170),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1138),
.B(n_750),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1140),
.B(n_1177),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1117),
.Y(n_1315)
);

CKINVDCx16_ASAP7_75t_R g1316 ( 
.A(n_1143),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1164),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1177),
.B(n_754),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1231),
.B(n_666),
.C(n_656),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1191),
.B(n_759),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1161),
.B(n_768),
.Y(n_1321)
);

NAND2xp33_ASAP7_75t_L g1322 ( 
.A(n_1192),
.B(n_769),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1162),
.B(n_781),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1187),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1179),
.B(n_910),
.C(n_653),
.Y(n_1325)
);

BUFx8_ASAP7_75t_L g1326 ( 
.A(n_1173),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1089),
.A2(n_657),
.B(n_662),
.C(n_654),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1163),
.B(n_799),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1141),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1157),
.B(n_807),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1188),
.B(n_809),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1193),
.B(n_817),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1223),
.B(n_1224),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1186),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1188),
.B(n_838),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1118),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1164),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1166),
.B(n_839),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1242),
.A2(n_1252),
.B(n_1097),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1198),
.B(n_854),
.Y(n_1340)
);

AO221x1_ASAP7_75t_L g1341 ( 
.A1(n_1143),
.A2(n_811),
.B1(n_861),
.B2(n_800),
.C(n_793),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1194),
.B(n_855),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1225),
.B(n_863),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1091),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1183),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1196),
.B(n_864),
.Y(n_1346)
);

BUFx8_ASAP7_75t_L g1347 ( 
.A(n_1114),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1124),
.B(n_878),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1114),
.B(n_887),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1124),
.B(n_891),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1236),
.B(n_893),
.Y(n_1351)
);

INVx5_ASAP7_75t_L g1352 ( 
.A(n_1103),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1168),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1237),
.B(n_896),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1239),
.B(n_900),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1192),
.B(n_904),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1168),
.B(n_932),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1136),
.B(n_921),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1146),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1178),
.B(n_939),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1232),
.B(n_1230),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1131),
.B(n_746),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1211),
.B(n_944),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1134),
.B(n_616),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1189),
.A2(n_915),
.B1(n_918),
.B2(n_910),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1145),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1135),
.B(n_918),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1092),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1265),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1096),
.B(n_921),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1133),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1139),
.B(n_669),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1219),
.Y(n_1373)
);

AND2x6_ASAP7_75t_SL g1374 ( 
.A(n_1110),
.B(n_811),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1133),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1190),
.B(n_674),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1183),
.Y(n_1377)
);

BUFx5_ASAP7_75t_L g1378 ( 
.A(n_1238),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1221),
.B(n_680),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1183),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1102),
.B(n_681),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1231),
.B(n_1250),
.C(n_1235),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1222),
.B(n_689),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1175),
.B(n_930),
.C(n_926),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1253),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1185),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1160),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1112),
.B(n_1115),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1111),
.B(n_702),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1176),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1197),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1213),
.B(n_966),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1207),
.B(n_966),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1119),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_1169),
.B(n_843),
.C(n_831),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1263),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1222),
.B(n_704),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1094),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1148),
.B(n_1095),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1151),
.B(n_1152),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1171),
.B(n_914),
.C(n_888),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1218),
.B(n_710),
.Y(n_1402)
);

OAI21xp33_ASAP7_75t_L g1403 ( 
.A1(n_1241),
.A2(n_1234),
.B(n_1233),
.Y(n_1403)
);

INVxp33_ASAP7_75t_L g1404 ( 
.A(n_1249),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1249),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1220),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1101),
.B(n_721),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1130),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1093),
.Y(n_1409)
);

INVxp33_ASAP7_75t_L g1410 ( 
.A(n_1094),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1101),
.B(n_723),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1272),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1209),
.B(n_1210),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1214),
.B(n_1215),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1229),
.B(n_1201),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1142),
.B(n_729),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1270),
.B(n_421),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1127),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1204),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1182),
.A2(n_676),
.B1(n_678),
.B2(n_673),
.C(n_670),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1243),
.B(n_732),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1247),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1248),
.Y(n_1423)
);

NOR3xp33_ASAP7_75t_L g1424 ( 
.A(n_1174),
.B(n_1106),
.C(n_1104),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1244),
.B(n_618),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1245),
.B(n_619),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1251),
.Y(n_1427)
);

INVxp33_ASAP7_75t_L g1428 ( 
.A(n_1099),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1254),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1255),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1120),
.B(n_734),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1121),
.B(n_736),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1263),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1125),
.B(n_737),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1250),
.B(n_626),
.C(n_620),
.Y(n_1435)
);

NOR3xp33_ASAP7_75t_L g1436 ( 
.A(n_1107),
.B(n_1109),
.C(n_1108),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1256),
.B(n_629),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1126),
.B(n_633),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1184),
.B(n_744),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1257),
.B(n_924),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1258),
.B(n_634),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1260),
.A2(n_690),
.B1(n_691),
.B2(n_684),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1262),
.B(n_635),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1264),
.B(n_763),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1268),
.B(n_764),
.Y(n_1445)
);

INVxp33_ASAP7_75t_L g1446 ( 
.A(n_1246),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1271),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1274),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1266),
.B(n_772),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1269),
.B(n_637),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1273),
.B(n_776),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1259),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_1261),
.B(n_655),
.C(n_638),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1267),
.B(n_660),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1093),
.Y(n_1455)
);

NOR3xp33_ASAP7_75t_L g1456 ( 
.A(n_1093),
.B(n_951),
.C(n_927),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1093),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1098),
.B(n_792),
.C(n_784),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1098),
.B(n_802),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1098),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1098),
.B(n_810),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1105),
.Y(n_1462)
);

INVxp67_ASAP7_75t_SL g1463 ( 
.A(n_1105),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1105),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1116),
.B(n_694),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1116),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1116),
.Y(n_1467)
);

BUFx5_ASAP7_75t_L g1468 ( 
.A(n_1170),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1205),
.B(n_665),
.Y(n_1469)
);

NOR3xp33_ASAP7_75t_L g1470 ( 
.A(n_1240),
.B(n_967),
.C(n_957),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1113),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1113),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1205),
.B(n_827),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1205),
.B(n_667),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1208),
.B(n_683),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1205),
.B(n_840),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1205),
.B(n_848),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_SL g1478 ( 
.A(n_1149),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1200),
.B(n_422),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1181),
.B(n_698),
.C(n_695),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1205),
.B(n_851),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1129),
.B(n_972),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1181),
.B(n_707),
.C(n_706),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1205),
.B(n_696),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1208),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1205),
.B(n_868),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1208),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1205),
.B(n_877),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1205),
.B(n_880),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1118),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1205),
.B(n_881),
.Y(n_1491)
);

INVx5_ASAP7_75t_L g1492 ( 
.A(n_1188),
.Y(n_1492)
);

AO221x1_ASAP7_75t_L g1493 ( 
.A1(n_1090),
.A2(n_867),
.B1(n_872),
.B2(n_865),
.C(n_861),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1208),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1208),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1208),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1208),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1205),
.B(n_885),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1090),
.B(n_705),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1205),
.B(n_890),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1205),
.B(n_717),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1208),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1113),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1164),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1164),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1205),
.B(n_919),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1090),
.B(n_712),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1205),
.B(n_949),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1208),
.B(n_718),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1167),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1327),
.A2(n_714),
.B(n_720),
.C(n_713),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1275),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1378),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1485),
.B(n_719),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1487),
.B(n_726),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1382),
.A2(n_872),
.B1(n_875),
.B2(n_867),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1490),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1333),
.B(n_875),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_899),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1347),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1317),
.B(n_1337),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1494),
.B(n_727),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1280),
.A2(n_937),
.B1(n_948),
.B2(n_899),
.Y(n_1523)
);

INVx5_ASAP7_75t_L g1524 ( 
.A(n_1465),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1347),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1499),
.B(n_728),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1374),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1495),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1496),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1326),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1497),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1502),
.Y(n_1532)
);

AO21x1_ASAP7_75t_L g1533 ( 
.A1(n_1339),
.A2(n_968),
.B(n_955),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_R g1534 ( 
.A(n_1368),
.B(n_730),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_731),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1308),
.B(n_733),
.Y(n_1536)
);

O2A1O1Ixp5_ASAP7_75t_L g1537 ( 
.A1(n_1402),
.A2(n_913),
.B(n_953),
.C(n_901),
.Y(n_1537)
);

BUFx4f_ASAP7_75t_L g1538 ( 
.A(n_1507),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1324),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1361),
.B(n_738),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1305),
.B(n_745),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1326),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1303),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1315),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1277),
.B(n_747),
.Y(n_1545)
);

NOR2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1329),
.B(n_761),
.Y(n_1546)
);

AO22x1_ASAP7_75t_L g1547 ( 
.A1(n_1309),
.A2(n_752),
.B1(n_755),
.B2(n_751),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1319),
.A2(n_725),
.B1(n_740),
.B2(n_722),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1374),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1469),
.B(n_756),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1334),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1474),
.B(n_757),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1499),
.B(n_767),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1353),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1501),
.B(n_773),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1447),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1377),
.A2(n_1380),
.B(n_1386),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1476),
.B(n_774),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1373),
.Y(n_1559)
);

NOR2x2_ASAP7_75t_L g1560 ( 
.A(n_1294),
.B(n_906),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1297),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1482),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1280),
.B(n_779),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1279),
.B(n_785),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1336),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1488),
.B(n_789),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1279),
.B(n_791),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1278),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1504),
.B(n_798),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1281),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1505),
.Y(n_1571)
);

NOR2x2_ASAP7_75t_L g1572 ( 
.A(n_1362),
.B(n_925),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1510),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1345),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1370),
.B(n_805),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1418),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1369),
.Y(n_1577)
);

NOR2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1366),
.B(n_965),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1344),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1352),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1489),
.B(n_804),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1447),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1352),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1319),
.A2(n_748),
.B1(n_753),
.B2(n_742),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1492),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1440),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1292),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_SL g1588 ( 
.A(n_1316),
.B(n_819),
.C(n_812),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1298),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1491),
.B(n_820),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1492),
.Y(n_1591)
);

NAND2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1447),
.B(n_765),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1398),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1362),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1492),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1359),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1479),
.A2(n_770),
.B(n_771),
.C(n_766),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1506),
.A2(n_782),
.B1(n_786),
.B2(n_783),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1366),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1310),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1508),
.A2(n_797),
.B1(n_808),
.B2(n_806),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1358),
.B(n_1439),
.Y(n_1602)
);

BUFx4f_ASAP7_75t_L g1603 ( 
.A(n_1399),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1415),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1345),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1475),
.B(n_823),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1385),
.Y(n_1607)
);

INVx3_ASAP7_75t_SL g1608 ( 
.A(n_1399),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1362),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_1465),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1286),
.B(n_814),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1286),
.B(n_816),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1367),
.Y(n_1613)
);

AO22x1_ASAP7_75t_L g1614 ( 
.A1(n_1410),
.A2(n_830),
.B1(n_832),
.B2(n_829),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1448),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1509),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1408),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_L g1618 ( 
.A(n_1312),
.B(n_833),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1371),
.B(n_837),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1365),
.B(n_842),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1276),
.B(n_818),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1416),
.B(n_844),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1470),
.A2(n_822),
.B1(n_834),
.B2(n_828),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1394),
.B(n_836),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1471),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1388),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1364),
.B(n_847),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1478),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1472),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1338),
.B(n_869),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1375),
.B(n_873),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1384),
.B(n_876),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1503),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1296),
.B(n_883),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1372),
.B(n_1285),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1387),
.Y(n_1637)
);

AND2x6_ASAP7_75t_SL g1638 ( 
.A(n_1399),
.B(n_845),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1438),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1376),
.B(n_892),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1478),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1405),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1428),
.A2(n_898),
.B1(n_902),
.B2(n_897),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1435),
.A2(n_846),
.B1(n_852),
.B2(n_849),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1406),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1454),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1345),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1390),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1391),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1423),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1450),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1473),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1480),
.B(n_856),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1477),
.B(n_907),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1481),
.B(n_908),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1288),
.A2(n_857),
.B1(n_860),
.B2(n_859),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1486),
.B(n_931),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1498),
.B(n_933),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1381),
.A2(n_862),
.B1(n_879),
.B2(n_871),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1483),
.B(n_882),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1340),
.B(n_940),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1419),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1500),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1359),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1330),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1396),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1325),
.A2(n_895),
.B1(n_903),
.B2(n_886),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1295),
.B(n_943),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1456),
.A2(n_909),
.B1(n_912),
.B2(n_905),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1301),
.B(n_950),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1396),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1403),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1389),
.A2(n_928),
.B1(n_929),
.B2(n_923),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1307),
.B(n_956),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1351),
.B(n_958),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1403),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1396),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1407),
.B(n_963),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1343),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1420),
.B(n_934),
.Y(n_1680)
);

INVx5_ASAP7_75t_L g1681 ( 
.A(n_1433),
.Y(n_1681)
);

INVx6_ASAP7_75t_L g1682 ( 
.A(n_1409),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1433),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1433),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1427),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1411),
.B(n_941),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_SL g1687 ( 
.A(n_1395),
.B(n_946),
.C(n_945),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1421),
.B(n_952),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1493),
.A2(n_960),
.B1(n_969),
.B2(n_959),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1354),
.B(n_777),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1457),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1357),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1430),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1442),
.A2(n_884),
.B1(n_954),
.B2(n_874),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1393),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1413),
.B(n_874),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1320),
.A2(n_983),
.B(n_981),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1442),
.B(n_874),
.Y(n_1698)
);

AND2x6_ASAP7_75t_L g1699 ( 
.A(n_1422),
.B(n_884),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_SL g1700 ( 
.A(n_1401),
.B(n_24),
.C(n_25),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1412),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_1284),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1432),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1392),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1331),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1335),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1453),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1355),
.B(n_884),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1341),
.A2(n_954),
.B1(n_1061),
.B2(n_1057),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1429),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1299),
.B(n_954),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1291),
.B(n_954),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1379),
.A2(n_1057),
.B1(n_1065),
.B2(n_1061),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1302),
.B(n_1293),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1282),
.B(n_25),
.Y(n_1715)
);

CKINVDCx14_ASAP7_75t_R g1716 ( 
.A(n_1321),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1360),
.B(n_26),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1383),
.A2(n_1057),
.B1(n_1065),
.B2(n_1061),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1449),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1409),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1437),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1332),
.B(n_1065),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_SL g1723 ( 
.A(n_1431),
.B(n_26),
.C(n_27),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1451),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1409),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1323),
.B(n_27),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1328),
.B(n_28),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1349),
.B(n_28),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1459),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1441),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1461),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1425),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1426),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1313),
.B(n_29),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1404),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1452),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1434),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1342),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1443),
.Y(n_1739)
);

NAND2x1p5_ASAP7_75t_L g1740 ( 
.A(n_1300),
.B(n_1414),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1287),
.A2(n_983),
.B(n_424),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1397),
.A2(n_1078),
.B1(n_1079),
.B2(n_1071),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1458),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1322),
.A2(n_1078),
.B1(n_1079),
.B2(n_1071),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1444),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_R g1746 ( 
.A(n_1283),
.B(n_1304),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1445),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1460),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1458),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1287),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1346),
.B(n_29),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1311),
.B(n_1079),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1436),
.B(n_30),
.C(n_31),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1356),
.B(n_30),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1400),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_R g1756 ( 
.A(n_1348),
.B(n_1087),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1363),
.A2(n_1088),
.B1(n_1087),
.B2(n_34),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1318),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1350),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1314),
.Y(n_1760)
);

BUFx4f_ASAP7_75t_L g1761 ( 
.A(n_1424),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1306),
.B(n_31),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1462),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1417),
.B(n_35),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_SL g1765 ( 
.A(n_1446),
.B(n_35),
.Y(n_1765)
);

BUFx12f_ASAP7_75t_L g1766 ( 
.A(n_1468),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1468),
.B(n_37),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1463),
.B(n_38),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1455),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1466),
.B(n_41),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1467),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1464),
.B(n_42),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1382),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1347),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1333),
.B(n_46),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1275),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1512),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1577),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1635),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1694),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1528),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1604),
.B(n_49),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1538),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1714),
.A2(n_435),
.B(n_434),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1616),
.B(n_50),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1616),
.B(n_51),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1523),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1694),
.A2(n_1597),
.B(n_1511),
.C(n_1656),
.Y(n_1788)
);

O2A1O1Ixp5_ASAP7_75t_L g1789 ( 
.A1(n_1690),
.A2(n_438),
.B(n_439),
.C(n_437),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1562),
.B(n_58),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1534),
.Y(n_1791)
);

XNOR2xp5_ASAP7_75t_L g1792 ( 
.A(n_1523),
.B(n_59),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1529),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1610),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1531),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1562),
.B(n_59),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1602),
.B(n_60),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1532),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1709),
.B(n_62),
.C(n_63),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1519),
.B(n_63),
.Y(n_1800)
);

BUFx8_ASAP7_75t_L g1801 ( 
.A(n_1520),
.Y(n_1801)
);

AND2x4_ASAP7_75t_SL g1802 ( 
.A(n_1624),
.B(n_64),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1704),
.A2(n_71),
.B(n_65),
.C(n_67),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1574),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1518),
.B(n_73),
.Y(n_1805)
);

CKINVDCx20_ASAP7_75t_R g1806 ( 
.A(n_1576),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1573),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1586),
.B(n_74),
.Y(n_1808)
);

NOR2xp67_ASAP7_75t_SL g1809 ( 
.A(n_1524),
.B(n_1774),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1776),
.B(n_75),
.Y(n_1810)
);

O2A1O1Ixp5_ASAP7_75t_L g1811 ( 
.A1(n_1533),
.A2(n_445),
.B(n_446),
.C(n_442),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1544),
.B(n_77),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1563),
.B(n_78),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1689),
.B(n_1753),
.C(n_1687),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1689),
.A2(n_82),
.B1(n_78),
.B2(n_81),
.Y(n_1815)
);

CKINVDCx8_ASAP7_75t_R g1816 ( 
.A(n_1638),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1613),
.B(n_81),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1705),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1526),
.B(n_86),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1543),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1551),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1527),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1706),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1559),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1517),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1524),
.Y(n_1826)
);

A2O1A1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1715),
.A2(n_98),
.B(n_94),
.C(n_95),
.Y(n_1827)
);

BUFx8_ASAP7_75t_L g1828 ( 
.A(n_1525),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1733),
.B(n_94),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1610),
.A2(n_99),
.B1(n_95),
.B2(n_98),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1538),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1615),
.B(n_100),
.Y(n_1832)
);

CKINVDCx14_ASAP7_75t_R g1833 ( 
.A(n_1603),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1730),
.B(n_101),
.Y(n_1834)
);

BUFx4f_ASAP7_75t_L g1835 ( 
.A(n_1608),
.Y(n_1835)
);

NOR3xp33_ASAP7_75t_SL g1836 ( 
.A(n_1593),
.B(n_101),
.C(n_102),
.Y(n_1836)
);

NOR2xp67_ASAP7_75t_SL g1837 ( 
.A(n_1641),
.B(n_103),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1549),
.Y(n_1838)
);

A2O1A1Ixp33_ASAP7_75t_SL g1839 ( 
.A1(n_1536),
.A2(n_456),
.B(n_457),
.C(n_455),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1565),
.B(n_104),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1553),
.B(n_104),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_R g1842 ( 
.A(n_1603),
.B(n_105),
.Y(n_1842)
);

AO21x2_ASAP7_75t_L g1843 ( 
.A1(n_1741),
.A2(n_464),
.B(n_460),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1665),
.B(n_106),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1539),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1557),
.A2(n_471),
.B(n_470),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1574),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1622),
.B(n_107),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1561),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1639),
.B(n_107),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1645),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1574),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1692),
.A2(n_473),
.B(n_472),
.Y(n_1853)
);

OR2x6_ASAP7_75t_SL g1854 ( 
.A(n_1703),
.B(n_110),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1651),
.A2(n_114),
.B(n_111),
.C(n_112),
.Y(n_1855)
);

INVx8_ASAP7_75t_L g1856 ( 
.A(n_1624),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1522),
.A2(n_475),
.B(n_474),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1521),
.B(n_115),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1568),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1522),
.A2(n_477),
.B(n_476),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1570),
.Y(n_1861)
);

NOR3xp33_ASAP7_75t_SL g1862 ( 
.A(n_1700),
.B(n_116),
.C(n_117),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1579),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1530),
.Y(n_1864)
);

CKINVDCx11_ASAP7_75t_R g1865 ( 
.A(n_1638),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1624),
.Y(n_1866)
);

NAND2xp33_ASAP7_75t_L g1867 ( 
.A(n_1605),
.B(n_483),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1556),
.Y(n_1868)
);

BUFx12f_ASAP7_75t_L g1869 ( 
.A(n_1542),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1588),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1662),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1730),
.B(n_116),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1680),
.B(n_1516),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1710),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1739),
.B(n_121),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1521),
.B(n_123),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1775),
.A2(n_1724),
.B(n_1719),
.C(n_1646),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1516),
.B(n_123),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_R g1879 ( 
.A(n_1716),
.B(n_124),
.Y(n_1879)
);

O2A1O1Ixp5_ASAP7_75t_L g1880 ( 
.A1(n_1728),
.A2(n_497),
.B(n_498),
.C(n_494),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1582),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1606),
.A2(n_503),
.B(n_500),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1592),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1592),
.B(n_125),
.Y(n_1884)
);

A2O1A1Ixp33_ASAP7_75t_SL g1885 ( 
.A1(n_1670),
.A2(n_507),
.B(n_508),
.C(n_505),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1594),
.B(n_126),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1739),
.B(n_1652),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1663),
.B(n_127),
.Y(n_1888)
);

AOI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1611),
.A2(n_1612),
.B1(n_1623),
.B2(n_1688),
.C(n_1575),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1695),
.A2(n_131),
.B(n_128),
.C(n_129),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1599),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1609),
.B(n_129),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1546),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1571),
.B(n_132),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1679),
.B(n_133),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1541),
.B(n_134),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1702),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_SL g1898 ( 
.A(n_1605),
.B(n_1647),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1755),
.B(n_135),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1732),
.B(n_136),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1554),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1643),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1535),
.B(n_138),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1771),
.A2(n_514),
.B(n_512),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1626),
.B(n_139),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1721),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1759),
.B(n_140),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1605),
.Y(n_1908)
);

NOR3xp33_ASAP7_75t_L g1909 ( 
.A(n_1614),
.B(n_141),
.C(n_142),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1698),
.B(n_142),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1620),
.B(n_143),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1766),
.Y(n_1912)
);

AO221x1_ASAP7_75t_L g1913 ( 
.A1(n_1643),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.C(n_147),
.Y(n_1913)
);

OAI21xp33_ASAP7_75t_L g1914 ( 
.A1(n_1598),
.A2(n_1601),
.B(n_1659),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1621),
.B(n_144),
.Y(n_1915)
);

OAI21xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1764),
.A2(n_149),
.B(n_150),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1737),
.B(n_150),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_SL g1918 ( 
.A(n_1738),
.B(n_151),
.C(n_153),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1621),
.B(n_154),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1598),
.B(n_154),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1601),
.B(n_155),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1764),
.A2(n_159),
.B1(n_156),
.B2(n_158),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1550),
.B(n_158),
.Y(n_1923)
);

INVx4_ASAP7_75t_L g1924 ( 
.A(n_1720),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_SL g1925 ( 
.A1(n_1768),
.A2(n_522),
.B(n_523),
.C(n_519),
.Y(n_1925)
);

BUFx4f_ASAP7_75t_L g1926 ( 
.A(n_1764),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1659),
.B(n_160),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1625),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1628),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1629),
.Y(n_1930)
);

O2A1O1Ixp33_ASAP7_75t_SL g1931 ( 
.A1(n_1767),
.A2(n_528),
.B(n_529),
.C(n_527),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1729),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_1932)
);

O2A1O1Ixp33_ASAP7_75t_L g1933 ( 
.A1(n_1686),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1578),
.B(n_166),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1587),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1673),
.B(n_167),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1650),
.B(n_168),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_SL g1938 ( 
.A(n_1773),
.B(n_168),
.C(n_169),
.Y(n_1938)
);

INVx4_ASAP7_75t_L g1939 ( 
.A(n_1720),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1552),
.B(n_169),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1589),
.Y(n_1941)
);

BUFx4f_ASAP7_75t_L g1942 ( 
.A(n_1740),
.Y(n_1942)
);

A2O1A1Ixp33_ASAP7_75t_L g1943 ( 
.A1(n_1731),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1673),
.B(n_1548),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1633),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1555),
.B(n_172),
.Y(n_1946)
);

CKINVDCx16_ASAP7_75t_R g1947 ( 
.A(n_1746),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1693),
.B(n_173),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1584),
.B(n_175),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1672),
.A2(n_178),
.B1(n_175),
.B2(n_176),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1676),
.A2(n_179),
.B1(n_176),
.B2(n_178),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1674),
.B(n_179),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1720),
.B(n_1681),
.Y(n_1953)
);

AND2x6_ASAP7_75t_L g1954 ( 
.A(n_1647),
.B(n_1513),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1773),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1584),
.B(n_182),
.Y(n_1956)
);

O2A1O1Ixp33_ASAP7_75t_L g1957 ( 
.A1(n_1558),
.A2(n_186),
.B(n_183),
.C(n_184),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1661),
.B(n_183),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1674),
.B(n_184),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1607),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1640),
.B(n_186),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1697),
.A2(n_548),
.B(n_545),
.Y(n_1962)
);

BUFx12f_ASAP7_75t_L g1963 ( 
.A(n_1617),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1653),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1630),
.B(n_191),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1685),
.B(n_193),
.Y(n_1966)
);

O2A1O1Ixp5_ASAP7_75t_L g1967 ( 
.A1(n_1708),
.A2(n_553),
.B(n_554),
.C(n_552),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1736),
.A2(n_557),
.B(n_555),
.Y(n_1968)
);

O2A1O1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1566),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_1969)
);

INVx3_ASAP7_75t_SL g1970 ( 
.A(n_1572),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1547),
.B(n_195),
.Y(n_1971)
);

INVx4_ASAP7_75t_L g1972 ( 
.A(n_1681),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1667),
.B(n_196),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1747),
.B(n_198),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1691),
.B(n_198),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1745),
.B(n_199),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1545),
.A2(n_559),
.B(n_558),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1725),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1769),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1514),
.B(n_202),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1515),
.B(n_203),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1540),
.B(n_203),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1668),
.B(n_204),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1769),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1600),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1644),
.B(n_205),
.Y(n_1986)
);

A2O1A1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1717),
.A2(n_1765),
.B(n_1537),
.C(n_1734),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1712),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1696),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1590),
.B(n_206),
.Y(n_1991)
);

AO32x1_ASAP7_75t_L g1992 ( 
.A1(n_1757),
.A2(n_207),
.A3(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_1992)
);

INVx3_ASAP7_75t_L g1993 ( 
.A(n_1725),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1696),
.B(n_208),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1726),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1685),
.B(n_212),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1682),
.Y(n_1997)
);

AOI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1741),
.A2(n_565),
.B(n_562),
.Y(n_1998)
);

AND2x6_ASAP7_75t_L g1999 ( 
.A(n_1647),
.B(n_213),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1678),
.A2(n_1669),
.B1(n_1740),
.B2(n_1727),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1682),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1684),
.B(n_213),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1618),
.A2(n_570),
.B(n_569),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1683),
.B(n_214),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1701),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1678),
.A2(n_574),
.B(n_573),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1632),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_2007)
);

NOR2xp67_ASAP7_75t_L g2008 ( 
.A(n_1735),
.B(n_218),
.Y(n_2008)
);

OA21x2_ASAP7_75t_L g2009 ( 
.A1(n_1770),
.A2(n_576),
.B(n_575),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1684),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1637),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1653),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1648),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1649),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1761),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1660),
.A2(n_1634),
.B1(n_1707),
.B2(n_1627),
.Y(n_2016)
);

CKINVDCx20_ASAP7_75t_R g2017 ( 
.A(n_1761),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1754),
.Y(n_2018)
);

BUFx6f_ASAP7_75t_L g2019 ( 
.A(n_1748),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1711),
.A2(n_579),
.B(n_578),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1569),
.B(n_1654),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1642),
.B(n_222),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1660),
.B(n_223),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1655),
.B(n_223),
.Y(n_2024)
);

INVx4_ASAP7_75t_L g2025 ( 
.A(n_1683),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1751),
.Y(n_2026)
);

O2A1O1Ixp33_ASAP7_75t_SL g2027 ( 
.A1(n_1762),
.A2(n_608),
.B(n_606),
.C(n_605),
.Y(n_2027)
);

O2A1O1Ixp33_ASAP7_75t_L g2028 ( 
.A1(n_1675),
.A2(n_224),
.B(n_226),
.C(n_227),
.Y(n_2028)
);

O2A1O1Ixp33_ASAP7_75t_L g2029 ( 
.A1(n_1657),
.A2(n_226),
.B(n_228),
.C(n_229),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1760),
.B(n_228),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1743),
.A2(n_583),
.B(n_582),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1758),
.Y(n_2032)
);

O2A1O1Ixp33_ASAP7_75t_SL g2033 ( 
.A1(n_1772),
.A2(n_599),
.B(n_597),
.C(n_596),
.Y(n_2033)
);

OR2x6_ASAP7_75t_L g2034 ( 
.A(n_1752),
.B(n_230),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1580),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1596),
.B(n_1664),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1658),
.B(n_230),
.Y(n_2037)
);

INVxp67_ASAP7_75t_L g2038 ( 
.A(n_1756),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1723),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_R g2040 ( 
.A(n_1699),
.B(n_1583),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1619),
.B(n_231),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1585),
.Y(n_2042)
);

AOI21xp33_ASAP7_75t_L g2043 ( 
.A1(n_1591),
.A2(n_1595),
.B(n_1631),
.Y(n_2043)
);

OAI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1749),
.A2(n_231),
.B(n_233),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1564),
.B(n_1567),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1722),
.B(n_234),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1666),
.B(n_235),
.Y(n_2047)
);

A2O1A1Ixp33_ASAP7_75t_L g2048 ( 
.A1(n_1713),
.A2(n_235),
.B(n_236),
.C(n_237),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1671),
.B(n_238),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1677),
.B(n_238),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1744),
.B(n_239),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1560),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1699),
.B(n_241),
.Y(n_2053)
);

AOI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1763),
.A2(n_588),
.B(n_587),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1699),
.B(n_242),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1763),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1699),
.B(n_243),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1744),
.B(n_243),
.Y(n_2058)
);

INVx5_ASAP7_75t_L g2059 ( 
.A(n_1742),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1718),
.Y(n_2060)
);

AOI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_1718),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1604),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_2062)
);

OR2x6_ASAP7_75t_L g2063 ( 
.A(n_1520),
.B(n_247),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1577),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1604),
.B(n_248),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1604),
.B(n_249),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1512),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1604),
.B(n_250),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1604),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1604),
.B(n_252),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1512),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1562),
.B(n_256),
.Y(n_2072)
);

BUFx4f_ASAP7_75t_L g2073 ( 
.A(n_1608),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1764),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1764),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_1610),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1636),
.A2(n_593),
.B(n_594),
.Y(n_2077)
);

A2O1A1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_1635),
.A2(n_263),
.B(n_265),
.C(n_266),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1604),
.B(n_265),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1512),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1562),
.B(n_266),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1524),
.B(n_269),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1604),
.B(n_269),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1577),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1764),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1604),
.B(n_276),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1764),
.A2(n_277),
.B1(n_279),
.B2(n_282),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1604),
.B(n_279),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1604),
.B(n_282),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1604),
.B(n_283),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1635),
.A2(n_285),
.B(n_286),
.C(n_287),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1577),
.B(n_288),
.Y(n_2092)
);

O2A1O1Ixp33_ASAP7_75t_L g2093 ( 
.A1(n_1635),
.A2(n_288),
.B(n_289),
.C(n_290),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1512),
.Y(n_2094)
);

INVx2_ASAP7_75t_SL g2095 ( 
.A(n_1538),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_L g2096 ( 
.A1(n_1635),
.A2(n_291),
.B(n_292),
.C(n_293),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1534),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_1636),
.A2(n_292),
.B(n_293),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1562),
.B(n_294),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1574),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1604),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_2101)
);

OAI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_1516),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1534),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1577),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1577),
.B(n_303),
.Y(n_2105)
);

AOI21x1_ASAP7_75t_L g2106 ( 
.A1(n_1750),
.A2(n_304),
.B(n_306),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1577),
.Y(n_2107)
);

INVx2_ASAP7_75t_SL g2108 ( 
.A(n_1538),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1604),
.B(n_306),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1562),
.B(n_307),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1604),
.B(n_307),
.Y(n_2111)
);

O2A1O1Ixp33_ASAP7_75t_L g2112 ( 
.A1(n_1635),
.A2(n_309),
.B(n_310),
.C(n_312),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1512),
.Y(n_2113)
);

NAND2x1p5_ASAP7_75t_L g2114 ( 
.A(n_1524),
.B(n_313),
.Y(n_2114)
);

BUFx10_ASAP7_75t_L g2115 ( 
.A(n_1802),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1778),
.Y(n_2116)
);

INVxp67_ASAP7_75t_SL g2117 ( 
.A(n_1926),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_1801),
.Y(n_2118)
);

BUFx2_ASAP7_75t_L g2119 ( 
.A(n_1806),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1820),
.B(n_314),
.Y(n_2120)
);

NAND2x1p5_ASAP7_75t_L g2121 ( 
.A(n_1926),
.B(n_315),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_1804),
.Y(n_2122)
);

NAND2x1p5_ASAP7_75t_L g2123 ( 
.A(n_1826),
.B(n_315),
.Y(n_2123)
);

BUFx12f_ASAP7_75t_L g2124 ( 
.A(n_1801),
.Y(n_2124)
);

AOI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_1914),
.A2(n_316),
.B1(n_317),
.B2(n_320),
.Y(n_2125)
);

OR2x6_ASAP7_75t_SL g2126 ( 
.A(n_1791),
.B(n_316),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_1828),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1821),
.B(n_402),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_SL g2129 ( 
.A(n_2063),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1856),
.Y(n_2130)
);

BUFx3_ASAP7_75t_L g2131 ( 
.A(n_1828),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_1998),
.A2(n_320),
.B(n_321),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2064),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1924),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_1845),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_1847),
.Y(n_2136)
);

INVx4_ASAP7_75t_L g2137 ( 
.A(n_1856),
.Y(n_2137)
);

BUFx2_ASAP7_75t_SL g2138 ( 
.A(n_1783),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1873),
.B(n_326),
.Y(n_2139)
);

BUFx2_ASAP7_75t_L g2140 ( 
.A(n_1856),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_2019),
.Y(n_2141)
);

OAI21x1_ASAP7_75t_L g2142 ( 
.A1(n_1846),
.A2(n_326),
.B(n_329),
.Y(n_2142)
);

INVx1_ASAP7_75t_SL g2143 ( 
.A(n_1825),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_2044),
.B(n_330),
.Y(n_2144)
);

INVx5_ASAP7_75t_L g2145 ( 
.A(n_1999),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2034),
.Y(n_2146)
);

INVx5_ASAP7_75t_L g2147 ( 
.A(n_1999),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_1924),
.Y(n_2148)
);

OAI21x1_ASAP7_75t_L g2149 ( 
.A1(n_1880),
.A2(n_333),
.B(n_335),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2084),
.Y(n_2150)
);

INVx6_ASAP7_75t_SL g2151 ( 
.A(n_2034),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_SL g2152 ( 
.A1(n_2074),
.A2(n_336),
.B(n_338),
.Y(n_2152)
);

AOI22x1_ASAP7_75t_L g2153 ( 
.A1(n_2006),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_2153)
);

AO21x2_ASAP7_75t_L g2154 ( 
.A1(n_1938),
.A2(n_341),
.B(n_343),
.Y(n_2154)
);

CKINVDCx14_ASAP7_75t_R g2155 ( 
.A(n_1833),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2104),
.Y(n_2156)
);

INVx4_ASAP7_75t_L g2157 ( 
.A(n_1835),
.Y(n_2157)
);

AO21x2_ASAP7_75t_L g2158 ( 
.A1(n_1987),
.A2(n_345),
.B(n_346),
.Y(n_2158)
);

BUFx12f_ASAP7_75t_L g2159 ( 
.A(n_1865),
.Y(n_2159)
);

INVx4_ASAP7_75t_L g2160 ( 
.A(n_1835),
.Y(n_2160)
);

OAI21x1_ASAP7_75t_L g2161 ( 
.A1(n_2031),
.A2(n_345),
.B(n_347),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2107),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1944),
.B(n_347),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_1939),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_SL g2165 ( 
.A1(n_1787),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_2165)
);

BUFx2_ASAP7_75t_R g2166 ( 
.A(n_1822),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_1990),
.B(n_348),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_2034),
.Y(n_2168)
);

BUFx3_ASAP7_75t_L g2169 ( 
.A(n_2019),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_1877),
.A2(n_349),
.B(n_350),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1866),
.B(n_351),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2073),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_2019),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_2009),
.A2(n_355),
.B(n_356),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_SL g2175 ( 
.A(n_2073),
.B(n_359),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1781),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1939),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1852),
.Y(n_2178)
);

NAND2x1p5_ASAP7_75t_L g2179 ( 
.A(n_1826),
.B(n_360),
.Y(n_2179)
);

OAI21x1_ASAP7_75t_L g2180 ( 
.A1(n_2054),
.A2(n_360),
.B(n_361),
.Y(n_2180)
);

INVx5_ASAP7_75t_L g2181 ( 
.A(n_1999),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1906),
.B(n_362),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1889),
.B(n_363),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_1852),
.Y(n_2184)
);

INVxp67_ASAP7_75t_SL g2185 ( 
.A(n_1908),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_1831),
.Y(n_2186)
);

INVx6_ASAP7_75t_L g2187 ( 
.A(n_1972),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1908),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1795),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_1912),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_2003),
.A2(n_363),
.B(n_365),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1908),
.Y(n_2192)
);

AO21x2_ASAP7_75t_L g2193 ( 
.A1(n_1925),
.A2(n_365),
.B(n_366),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1794),
.B(n_402),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1798),
.Y(n_2195)
);

BUFx2_ASAP7_75t_SL g2196 ( 
.A(n_2095),
.Y(n_2196)
);

BUFx2_ASAP7_75t_L g2197 ( 
.A(n_1807),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_2097),
.Y(n_2198)
);

OAI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_1788),
.A2(n_366),
.B(n_367),
.Y(n_2199)
);

INVxp67_ASAP7_75t_SL g2200 ( 
.A(n_2100),
.Y(n_2200)
);

INVx1_ASAP7_75t_SL g2201 ( 
.A(n_1900),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1887),
.B(n_367),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_2025),
.Y(n_2203)
);

NAND2x1p5_ASAP7_75t_L g2204 ( 
.A(n_1809),
.B(n_2025),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_L g2205 ( 
.A1(n_1811),
.A2(n_2020),
.B(n_1784),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_1857),
.A2(n_368),
.B(n_369),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_1860),
.A2(n_368),
.B(n_370),
.Y(n_2207)
);

INVx4_ASAP7_75t_L g2208 ( 
.A(n_1869),
.Y(n_2208)
);

BUFx3_ASAP7_75t_L g2209 ( 
.A(n_1912),
.Y(n_2209)
);

NAND2x1p5_ASAP7_75t_L g2210 ( 
.A(n_2076),
.B(n_370),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_1952),
.A2(n_371),
.B(n_372),
.Y(n_2211)
);

INVx5_ASAP7_75t_L g2212 ( 
.A(n_1999),
.Y(n_2212)
);

AOI21x1_ASAP7_75t_L g2213 ( 
.A1(n_2106),
.A2(n_371),
.B(n_372),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1868),
.Y(n_2214)
);

OAI21x1_ASAP7_75t_SL g2215 ( 
.A1(n_2074),
.A2(n_375),
.B(n_376),
.Y(n_2215)
);

AOI22x1_ASAP7_75t_L g2216 ( 
.A1(n_1882),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_2216)
);

INVx4_ASAP7_75t_L g2217 ( 
.A(n_2063),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1777),
.Y(n_2218)
);

OAI21x1_ASAP7_75t_L g2219 ( 
.A1(n_1977),
.A2(n_378),
.B(n_379),
.Y(n_2219)
);

AO21x2_ASAP7_75t_L g2220 ( 
.A1(n_1839),
.A2(n_380),
.B(n_381),
.Y(n_2220)
);

INVx8_ASAP7_75t_L g2221 ( 
.A(n_2063),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2076),
.B(n_400),
.Y(n_2222)
);

OAI21x1_ASAP7_75t_L g2223 ( 
.A1(n_2010),
.A2(n_380),
.B(n_381),
.Y(n_2223)
);

AOI22xp33_ASAP7_75t_L g2224 ( 
.A1(n_1814),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_2224)
);

BUFx2_ASAP7_75t_SL g2225 ( 
.A(n_2108),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1793),
.Y(n_2226)
);

INVx1_ASAP7_75t_SL g2227 ( 
.A(n_1900),
.Y(n_2227)
);

INVx1_ASAP7_75t_SL g2228 ( 
.A(n_1937),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_1942),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_1881),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1997),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_1937),
.Y(n_2232)
);

AO21x2_ASAP7_75t_L g2233 ( 
.A1(n_1885),
.A2(n_382),
.B(n_384),
.Y(n_2233)
);

AO21x2_ASAP7_75t_L g2234 ( 
.A1(n_1843),
.A2(n_385),
.B(n_386),
.Y(n_2234)
);

OAI21x1_ASAP7_75t_L g2235 ( 
.A1(n_1968),
.A2(n_386),
.B(n_388),
.Y(n_2235)
);

INVx3_ASAP7_75t_L g2236 ( 
.A(n_1978),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1874),
.B(n_388),
.Y(n_2237)
);

OAI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_1959),
.A2(n_389),
.B(n_390),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1851),
.Y(n_2239)
);

INVx4_ASAP7_75t_SL g2240 ( 
.A(n_1954),
.Y(n_2240)
);

OAI21x1_ASAP7_75t_L g2241 ( 
.A1(n_1962),
.A2(n_390),
.B(n_393),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_2000),
.B(n_393),
.Y(n_2242)
);

OAI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_2016),
.A2(n_395),
.B(n_396),
.Y(n_2243)
);

OAI21x1_ASAP7_75t_SL g2244 ( 
.A1(n_2075),
.A2(n_397),
.B(n_398),
.Y(n_2244)
);

INVx4_ASAP7_75t_L g2245 ( 
.A(n_1864),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_1991),
.A2(n_1961),
.B(n_1782),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2067),
.Y(n_2247)
);

BUFx2_ASAP7_75t_SL g2248 ( 
.A(n_1816),
.Y(n_2248)
);

CKINVDCx11_ASAP7_75t_R g2249 ( 
.A(n_1854),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1813),
.B(n_2026),
.Y(n_2250)
);

INVx4_ASAP7_75t_L g2251 ( 
.A(n_2114),
.Y(n_2251)
);

CKINVDCx6p67_ASAP7_75t_R g2252 ( 
.A(n_1970),
.Y(n_2252)
);

BUFx2_ASAP7_75t_R g2253 ( 
.A(n_1838),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2071),
.Y(n_2254)
);

INVxp33_ASAP7_75t_L g2255 ( 
.A(n_1844),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_2021),
.B(n_1819),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_1797),
.B(n_1911),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2080),
.Y(n_2258)
);

NAND2x1p5_ASAP7_75t_L g2259 ( 
.A(n_1942),
.B(n_1978),
.Y(n_2259)
);

INVxp67_ASAP7_75t_L g2260 ( 
.A(n_1829),
.Y(n_2260)
);

AO21x2_ASAP7_75t_L g2261 ( 
.A1(n_1843),
.A2(n_1799),
.B(n_2049),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2094),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_1966),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_1954),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2113),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1824),
.Y(n_2266)
);

NAND2x1p5_ASAP7_75t_L g2267 ( 
.A(n_1993),
.B(n_1829),
.Y(n_2267)
);

INVxp67_ASAP7_75t_SL g2268 ( 
.A(n_2092),
.Y(n_2268)
);

OA21x2_ASAP7_75t_L g2269 ( 
.A1(n_1799),
.A2(n_1789),
.B(n_2077),
.Y(n_2269)
);

BUFx3_ASAP7_75t_L g2270 ( 
.A(n_1954),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1863),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1928),
.Y(n_2272)
);

AO21x2_ASAP7_75t_L g2273 ( 
.A1(n_2050),
.A2(n_2033),
.B(n_1931),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1930),
.Y(n_2274)
);

OR2x4_ASAP7_75t_L g2275 ( 
.A(n_1971),
.B(n_1840),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_1898),
.A2(n_1896),
.B(n_1980),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1871),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1945),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_2056),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_SL g2280 ( 
.A1(n_2075),
.A2(n_2087),
.B(n_2085),
.Y(n_2280)
);

AO21x2_ASAP7_75t_L g2281 ( 
.A1(n_2027),
.A2(n_2046),
.B(n_2002),
.Y(n_2281)
);

INVx6_ASAP7_75t_L g2282 ( 
.A(n_1963),
.Y(n_2282)
);

OAI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2065),
.A2(n_2068),
.B(n_2066),
.Y(n_2283)
);

BUFx10_ASAP7_75t_L g2284 ( 
.A(n_1934),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_1808),
.B(n_2099),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_1800),
.B(n_1989),
.Y(n_2286)
);

OAI21x1_ASAP7_75t_L g2287 ( 
.A1(n_1967),
.A2(n_1904),
.B(n_1853),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1849),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_1993),
.Y(n_2289)
);

NAND2x1p5_ASAP7_75t_L g2290 ( 
.A(n_2092),
.B(n_2105),
.Y(n_2290)
);

BUFx2_ASAP7_75t_L g2291 ( 
.A(n_1842),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1859),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1935),
.Y(n_2293)
);

INVx1_ASAP7_75t_SL g2294 ( 
.A(n_1948),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1861),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_1954),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_2056),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_1988),
.B(n_2015),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2070),
.A2(n_2083),
.B(n_2079),
.Y(n_2299)
);

INVx2_ASAP7_75t_SL g2300 ( 
.A(n_1948),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1941),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2105),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2110),
.B(n_1947),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2086),
.A2(n_2089),
.B(n_2088),
.Y(n_2304)
);

INVx6_ASAP7_75t_SL g2305 ( 
.A(n_1966),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_2056),
.Y(n_2306)
);

OR2x6_ASAP7_75t_L g2307 ( 
.A(n_2114),
.B(n_2052),
.Y(n_2307)
);

CKINVDCx20_ASAP7_75t_R g2308 ( 
.A(n_2103),
.Y(n_2308)
);

INVx4_ASAP7_75t_L g2309 ( 
.A(n_2004),
.Y(n_2309)
);

INVx5_ASAP7_75t_L g2310 ( 
.A(n_1886),
.Y(n_2310)
);

BUFx3_ASAP7_75t_L g2311 ( 
.A(n_1891),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1901),
.Y(n_2312)
);

BUFx2_ASAP7_75t_R g2313 ( 
.A(n_1870),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1985),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_1796),
.B(n_1883),
.Y(n_2315)
);

BUFx2_ASAP7_75t_L g2316 ( 
.A(n_1929),
.Y(n_2316)
);

NAND2x1p5_ASAP7_75t_L g2317 ( 
.A(n_1953),
.B(n_1994),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_2036),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_1893),
.Y(n_2319)
);

OAI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2090),
.A2(n_2111),
.B(n_2109),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1903),
.B(n_1848),
.Y(n_2321)
);

OA21x2_ASAP7_75t_L g2322 ( 
.A1(n_2078),
.A2(n_2096),
.B(n_1943),
.Y(n_2322)
);

BUFx2_ASAP7_75t_SL g2323 ( 
.A(n_1934),
.Y(n_2323)
);

NAND2x1p5_ASAP7_75t_L g2324 ( 
.A(n_1907),
.B(n_1886),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_1792),
.B(n_1878),
.Y(n_2325)
);

BUFx2_ASAP7_75t_SL g2326 ( 
.A(n_2017),
.Y(n_2326)
);

OAI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_1817),
.A2(n_1940),
.B(n_1923),
.Y(n_2327)
);

INVx4_ASAP7_75t_L g2328 ( 
.A(n_1892),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_2036),
.Y(n_2329)
);

NAND2x1p5_ASAP7_75t_L g2330 ( 
.A(n_1907),
.B(n_1892),
.Y(n_2330)
);

INVx3_ASAP7_75t_SL g2331 ( 
.A(n_2039),
.Y(n_2331)
);

OA21x2_ASAP7_75t_L g2332 ( 
.A1(n_1932),
.A2(n_1823),
.B(n_1818),
.Y(n_2332)
);

BUFx2_ASAP7_75t_R g2333 ( 
.A(n_2060),
.Y(n_2333)
);

AO21x2_ASAP7_75t_L g2334 ( 
.A1(n_1810),
.A2(n_1867),
.B(n_1910),
.Y(n_2334)
);

CKINVDCx16_ASAP7_75t_R g2335 ( 
.A(n_1879),
.Y(n_2335)
);

AO21x2_ASAP7_75t_L g2336 ( 
.A1(n_1981),
.A2(n_1888),
.B(n_2098),
.Y(n_2336)
);

INVx1_ASAP7_75t_SL g2337 ( 
.A(n_2045),
.Y(n_2337)
);

INVx1_ASAP7_75t_SL g2338 ( 
.A(n_1960),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2011),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2005),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_2040),
.Y(n_2341)
);

AO21x2_ASAP7_75t_L g2342 ( 
.A1(n_1976),
.A2(n_2058),
.B(n_2051),
.Y(n_2342)
);

AO21x2_ASAP7_75t_L g2343 ( 
.A1(n_1890),
.A2(n_1803),
.B(n_2048),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2013),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_1841),
.B(n_1946),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2014),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2032),
.Y(n_2347)
);

BUFx3_ASAP7_75t_L g2348 ( 
.A(n_2001),
.Y(n_2348)
);

OR2x6_ASAP7_75t_L g2349 ( 
.A(n_2038),
.B(n_1815),
.Y(n_2349)
);

INVx3_ASAP7_75t_L g2350 ( 
.A(n_2035),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1950),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_2042),
.B(n_1958),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1950),
.Y(n_2353)
);

INVx1_ASAP7_75t_SL g2354 ( 
.A(n_1915),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_1919),
.Y(n_2355)
);

OAI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_1785),
.A2(n_1786),
.B(n_2024),
.Y(n_2356)
);

OAI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2037),
.A2(n_1834),
.B(n_1872),
.Y(n_2357)
);

AOI22x1_ASAP7_75t_L g2358 ( 
.A1(n_2018),
.A2(n_1965),
.B1(n_2057),
.B2(n_1916),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2059),
.Y(n_2359)
);

AO21x2_ASAP7_75t_L g2360 ( 
.A1(n_1827),
.A2(n_1855),
.B(n_1884),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1951),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_1805),
.B(n_1895),
.Y(n_2362)
);

INVxp67_ASAP7_75t_SL g2363 ( 
.A(n_1979),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1951),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2059),
.Y(n_2365)
);

OAI21x1_ASAP7_75t_L g2366 ( 
.A1(n_1779),
.A2(n_2091),
.B(n_2112),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1927),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2059),
.Y(n_2368)
);

OA21x2_ASAP7_75t_L g2369 ( 
.A1(n_1949),
.A2(n_1956),
.B(n_2055),
.Y(n_2369)
);

INVx3_ASAP7_75t_SL g2370 ( 
.A(n_1858),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1920),
.Y(n_2371)
);

HB1xp67_ASAP7_75t_L g2372 ( 
.A(n_1996),
.Y(n_2372)
);

INVx5_ASAP7_75t_L g2373 ( 
.A(n_1922),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1921),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_1790),
.B(n_2072),
.Y(n_2375)
);

HB1xp67_ASAP7_75t_L g2376 ( 
.A(n_1875),
.Y(n_2376)
);

BUFx3_ASAP7_75t_L g2377 ( 
.A(n_1850),
.Y(n_2377)
);

HB1xp67_ASAP7_75t_L g2378 ( 
.A(n_1979),
.Y(n_2378)
);

OA21x2_ASAP7_75t_L g2379 ( 
.A1(n_2053),
.A2(n_2061),
.B(n_2047),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_1812),
.B(n_2081),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1936),
.Y(n_2381)
);

AO21x2_ASAP7_75t_L g2382 ( 
.A1(n_1975),
.A2(n_2008),
.B(n_2023),
.Y(n_2382)
);

OAI21x1_ASAP7_75t_L g2383 ( 
.A1(n_2093),
.A2(n_2082),
.B(n_1933),
.Y(n_2383)
);

INVx4_ASAP7_75t_L g2384 ( 
.A(n_1837),
.Y(n_2384)
);

AO21x2_ASAP7_75t_L g2385 ( 
.A1(n_1984),
.A2(n_1909),
.B(n_1957),
.Y(n_2385)
);

AO21x2_ASAP7_75t_L g2386 ( 
.A1(n_1984),
.A2(n_1969),
.B(n_1913),
.Y(n_2386)
);

BUFx3_ASAP7_75t_L g2387 ( 
.A(n_1973),
.Y(n_2387)
);

AO21x2_ASAP7_75t_L g2388 ( 
.A1(n_1995),
.A2(n_2029),
.B(n_2102),
.Y(n_2388)
);

OAI21x1_ASAP7_75t_L g2389 ( 
.A1(n_2028),
.A2(n_2030),
.B(n_1780),
.Y(n_2389)
);

INVxp67_ASAP7_75t_SL g2390 ( 
.A(n_1995),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1986),
.Y(n_2391)
);

AO21x2_ASAP7_75t_L g2392 ( 
.A1(n_1899),
.A2(n_1876),
.B(n_1832),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_1992),
.Y(n_2393)
);

BUFx2_ASAP7_75t_L g2394 ( 
.A(n_1918),
.Y(n_2394)
);

CKINVDCx20_ASAP7_75t_R g2395 ( 
.A(n_1815),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2043),
.Y(n_2396)
);

AOI21x1_ASAP7_75t_L g2397 ( 
.A1(n_1905),
.A2(n_2022),
.B(n_1894),
.Y(n_2397)
);

CKINVDCx20_ASAP7_75t_R g2398 ( 
.A(n_1836),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_1974),
.B(n_1983),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2062),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_1982),
.Y(n_2401)
);

AOI22x1_ASAP7_75t_L g2402 ( 
.A1(n_1862),
.A2(n_1992),
.B1(n_1955),
.B2(n_2041),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_1917),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2069),
.Y(n_2404)
);

BUFx8_ASAP7_75t_SL g2405 ( 
.A(n_1830),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2101),
.Y(n_2406)
);

BUFx2_ASAP7_75t_L g2407 ( 
.A(n_1897),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_1902),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_1992),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2116),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2124),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2133),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2339),
.Y(n_2413)
);

INVx1_ASAP7_75t_SL g2414 ( 
.A(n_2228),
.Y(n_2414)
);

BUFx2_ASAP7_75t_L g2415 ( 
.A(n_2151),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2150),
.Y(n_2416)
);

INVxp67_ASAP7_75t_SL g2417 ( 
.A(n_2290),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2156),
.Y(n_2418)
);

CKINVDCx20_ASAP7_75t_R g2419 ( 
.A(n_2124),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2344),
.Y(n_2420)
);

HB1xp67_ASAP7_75t_L g2421 ( 
.A(n_2143),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_2118),
.Y(n_2422)
);

OAI21xp33_ASAP7_75t_SL g2423 ( 
.A1(n_2268),
.A2(n_2390),
.B(n_2144),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2162),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2176),
.Y(n_2425)
);

AO21x1_ASAP7_75t_L g2426 ( 
.A1(n_2144),
.A2(n_2007),
.B(n_2012),
.Y(n_2426)
);

CKINVDCx20_ASAP7_75t_R g2427 ( 
.A(n_2155),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_2309),
.Y(n_2428)
);

AOI22xp33_ASAP7_75t_L g2429 ( 
.A1(n_2280),
.A2(n_1964),
.B1(n_2407),
.B2(n_2378),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2325),
.B(n_2256),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2256),
.B(n_2167),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2351),
.B(n_2353),
.Y(n_2432)
);

AOI21x1_ASAP7_75t_L g2433 ( 
.A1(n_2276),
.A2(n_2174),
.B(n_2393),
.Y(n_2433)
);

OR2x6_ASAP7_75t_L g2434 ( 
.A(n_2221),
.B(n_2267),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2349),
.B(n_2275),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2268),
.A2(n_2378),
.B1(n_2363),
.B2(n_2151),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2189),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2118),
.Y(n_2438)
);

OAI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2395),
.A2(n_2349),
.B1(n_2175),
.B2(n_2221),
.Y(n_2439)
);

INVx3_ASAP7_75t_L g2440 ( 
.A(n_2309),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_2127),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2218),
.B(n_2226),
.Y(n_2442)
);

OAI21x1_ASAP7_75t_L g2443 ( 
.A1(n_2149),
.A2(n_2205),
.B(n_2287),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2195),
.Y(n_2444)
);

NAND2x1p5_ASAP7_75t_L g2445 ( 
.A(n_2145),
.B(n_2147),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2288),
.Y(n_2446)
);

BUFx2_ASAP7_75t_R g2447 ( 
.A(n_2127),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2292),
.Y(n_2448)
);

INVx2_ASAP7_75t_SL g2449 ( 
.A(n_2131),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2295),
.Y(n_2450)
);

CKINVDCx20_ASAP7_75t_R g2451 ( 
.A(n_2155),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2117),
.B(n_2145),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_L g2453 ( 
.A1(n_2363),
.A2(n_2408),
.B1(n_2345),
.B2(n_2405),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_SL g2454 ( 
.A1(n_2395),
.A2(n_2221),
.B1(n_2129),
.B2(n_2217),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2361),
.B(n_2364),
.Y(n_2455)
);

INVx4_ASAP7_75t_L g2456 ( 
.A(n_2131),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2312),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2340),
.Y(n_2458)
);

HB1xp67_ASAP7_75t_L g2459 ( 
.A(n_2197),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2266),
.Y(n_2460)
);

BUFx2_ASAP7_75t_R g2461 ( 
.A(n_2248),
.Y(n_2461)
);

OAI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2349),
.A2(n_2151),
.B1(n_2217),
.B2(n_2324),
.Y(n_2462)
);

BUFx4_ASAP7_75t_SL g2463 ( 
.A(n_2308),
.Y(n_2463)
);

AOI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_2408),
.A2(n_2345),
.B1(n_2405),
.B2(n_2257),
.Y(n_2464)
);

AOI22xp33_ASAP7_75t_L g2465 ( 
.A1(n_2257),
.A2(n_2129),
.B1(n_2401),
.B2(n_2362),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2232),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2401),
.A2(n_2362),
.B1(n_2380),
.B2(n_2394),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2271),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2272),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2274),
.Y(n_2470)
);

BUFx4f_ASAP7_75t_SL g2471 ( 
.A(n_2159),
.Y(n_2471)
);

INVx2_ASAP7_75t_SL g2472 ( 
.A(n_2282),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2278),
.Y(n_2473)
);

OAI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_2324),
.A2(n_2330),
.B1(n_2310),
.B2(n_2291),
.Y(n_2474)
);

AOI22xp33_ASAP7_75t_SL g2475 ( 
.A1(n_2146),
.A2(n_2168),
.B1(n_2323),
.B2(n_2328),
.Y(n_2475)
);

OA21x2_ASAP7_75t_L g2476 ( 
.A1(n_2393),
.A2(n_2409),
.B(n_2132),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2239),
.Y(n_2477)
);

BUFx12f_ASAP7_75t_L g2478 ( 
.A(n_2208),
.Y(n_2478)
);

NAND2x1p5_ASAP7_75t_L g2479 ( 
.A(n_2145),
.B(n_2147),
.Y(n_2479)
);

CKINVDCx14_ASAP7_75t_R g2480 ( 
.A(n_2249),
.Y(n_2480)
);

INVx1_ASAP7_75t_SL g2481 ( 
.A(n_2294),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2247),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2254),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2371),
.B(n_2374),
.Y(n_2484)
);

BUFx2_ASAP7_75t_R g2485 ( 
.A(n_2198),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2258),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_2305),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2139),
.B(n_2262),
.Y(n_2488)
);

AOI22xp33_ASAP7_75t_SL g2489 ( 
.A1(n_2146),
.A2(n_2168),
.B1(n_2328),
.B2(n_2117),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2265),
.B(n_2346),
.Y(n_2490)
);

INVx6_ASAP7_75t_L g2491 ( 
.A(n_2208),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2347),
.Y(n_2492)
);

BUFx2_ASAP7_75t_SL g2493 ( 
.A(n_2157),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2347),
.Y(n_2494)
);

AOI222xp33_ASAP7_75t_L g2495 ( 
.A1(n_2249),
.A2(n_2250),
.B1(n_2390),
.B2(n_2302),
.C1(n_2260),
.C2(n_2159),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2166),
.Y(n_2496)
);

BUFx12f_ASAP7_75t_L g2497 ( 
.A(n_2157),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2346),
.B(n_2337),
.Y(n_2498)
);

INVx6_ASAP7_75t_L g2499 ( 
.A(n_2160),
.Y(n_2499)
);

INVx6_ASAP7_75t_L g2500 ( 
.A(n_2160),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_2253),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2120),
.Y(n_2502)
);

AOI22xp33_ASAP7_75t_L g2503 ( 
.A1(n_2380),
.A2(n_2399),
.B1(n_2250),
.B2(n_2375),
.Y(n_2503)
);

BUFx10_ASAP7_75t_L g2504 ( 
.A(n_2282),
.Y(n_2504)
);

NAND2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2147),
.B(n_2181),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2267),
.Y(n_2506)
);

BUFx2_ASAP7_75t_SL g2507 ( 
.A(n_2137),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2128),
.Y(n_2508)
);

BUFx3_ASAP7_75t_L g2509 ( 
.A(n_2135),
.Y(n_2509)
);

INVx6_ASAP7_75t_L g2510 ( 
.A(n_2137),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_SL g2511 ( 
.A1(n_2358),
.A2(n_2330),
.B1(n_2310),
.B2(n_2263),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2398),
.A2(n_2242),
.B1(n_2183),
.B2(n_2406),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2128),
.Y(n_2513)
);

INVx1_ASAP7_75t_SL g2514 ( 
.A(n_2201),
.Y(n_2514)
);

INVx4_ASAP7_75t_L g2515 ( 
.A(n_2147),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2182),
.B(n_2227),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2403),
.A2(n_2372),
.B1(n_2404),
.B2(n_2400),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2371),
.B(n_2374),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2310),
.A2(n_2260),
.B1(n_2302),
.B2(n_2181),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2237),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2403),
.A2(n_2387),
.B1(n_2402),
.B2(n_2255),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2277),
.Y(n_2522)
);

AND2x4_ASAP7_75t_L g2523 ( 
.A(n_2181),
.B(n_2212),
.Y(n_2523)
);

BUFx4_ASAP7_75t_SL g2524 ( 
.A(n_2308),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2251),
.Y(n_2525)
);

OAI21x1_ASAP7_75t_SL g2526 ( 
.A1(n_2251),
.A2(n_2215),
.B(n_2152),
.Y(n_2526)
);

INVxp67_ASAP7_75t_SL g2527 ( 
.A(n_2263),
.Y(n_2527)
);

NAND2x1p5_ASAP7_75t_L g2528 ( 
.A(n_2181),
.B(n_2212),
.Y(n_2528)
);

BUFx3_ASAP7_75t_L g2529 ( 
.A(n_2135),
.Y(n_2529)
);

BUFx4f_ASAP7_75t_SL g2530 ( 
.A(n_2252),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2381),
.B(n_2367),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2293),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_2285),
.B(n_2130),
.Y(n_2533)
);

AOI21x1_ASAP7_75t_L g2534 ( 
.A1(n_2269),
.A2(n_2199),
.B(n_2213),
.Y(n_2534)
);

AOI22xp33_ASAP7_75t_L g2535 ( 
.A1(n_2387),
.A2(n_2255),
.B1(n_2377),
.B2(n_2242),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2301),
.Y(n_2536)
);

AOI21x1_ASAP7_75t_L g2537 ( 
.A1(n_2269),
.A2(n_2376),
.B(n_2369),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2301),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2377),
.A2(n_2373),
.B1(n_2398),
.B2(n_2386),
.Y(n_2539)
);

OAI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_2310),
.A2(n_2212),
.B1(n_2305),
.B2(n_2275),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2314),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2198),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2314),
.Y(n_2543)
);

AOI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2373),
.A2(n_2386),
.B1(n_2307),
.B2(n_2355),
.Y(n_2544)
);

INVx6_ASAP7_75t_L g2545 ( 
.A(n_2282),
.Y(n_2545)
);

AO21x2_ASAP7_75t_L g2546 ( 
.A1(n_2261),
.A2(n_2158),
.B(n_2234),
.Y(n_2546)
);

CKINVDCx20_ASAP7_75t_R g2547 ( 
.A(n_2119),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2259),
.Y(n_2548)
);

CKINVDCx11_ASAP7_75t_R g2549 ( 
.A(n_2126),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2381),
.B(n_2391),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2210),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2212),
.A2(n_2305),
.B1(n_2125),
.B2(n_2165),
.Y(n_2552)
);

AOI22xp33_ASAP7_75t_L g2553 ( 
.A1(n_2373),
.A2(n_2307),
.B1(n_2355),
.B2(n_2327),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2214),
.Y(n_2554)
);

BUFx10_ASAP7_75t_L g2555 ( 
.A(n_2172),
.Y(n_2555)
);

HB1xp67_ASAP7_75t_L g2556 ( 
.A(n_2140),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2204),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2210),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2187),
.Y(n_2559)
);

AOI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2273),
.A2(n_2261),
.B(n_2283),
.Y(n_2560)
);

INVx2_ASAP7_75t_SL g2561 ( 
.A(n_2115),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2350),
.Y(n_2562)
);

OAI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2121),
.A2(n_2335),
.B1(n_2307),
.B2(n_2370),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_2373),
.A2(n_2246),
.B1(n_2370),
.B2(n_2165),
.Y(n_2564)
);

BUFx2_ASAP7_75t_L g2565 ( 
.A(n_2204),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2171),
.B(n_2121),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_SL g2567 ( 
.A1(n_2244),
.A2(n_2123),
.B1(n_2179),
.B2(n_2284),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2391),
.B(n_2163),
.Y(n_2568)
);

CKINVDCx20_ASAP7_75t_R g2569 ( 
.A(n_2316),
.Y(n_2569)
);

INVx6_ASAP7_75t_L g2570 ( 
.A(n_2115),
.Y(n_2570)
);

AND2x6_ASAP7_75t_L g2571 ( 
.A(n_2359),
.B(n_2368),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2303),
.B(n_2333),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2194),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2194),
.Y(n_2574)
);

NAND2x1p5_ASAP7_75t_L g2575 ( 
.A(n_2203),
.B(n_2229),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2223),
.Y(n_2576)
);

NAND2x1p5_ASAP7_75t_L g2577 ( 
.A(n_2203),
.B(n_2264),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2300),
.B(n_2284),
.Y(n_2578)
);

OAI22xp33_ASAP7_75t_L g2579 ( 
.A1(n_2123),
.A2(n_2179),
.B1(n_2321),
.B2(n_2341),
.Y(n_2579)
);

AO21x1_ASAP7_75t_L g2580 ( 
.A1(n_2170),
.A2(n_2243),
.B(n_2222),
.Y(n_2580)
);

AO21x1_ASAP7_75t_L g2581 ( 
.A1(n_2170),
.A2(n_2222),
.B(n_2211),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2222),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2298),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2298),
.Y(n_2584)
);

INVx4_ASAP7_75t_L g2585 ( 
.A(n_2245),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2385),
.A2(n_2388),
.B1(n_2286),
.B2(n_2352),
.Y(n_2586)
);

CKINVDCx11_ASAP7_75t_R g2587 ( 
.A(n_2331),
.Y(n_2587)
);

BUFx2_ASAP7_75t_SL g2588 ( 
.A(n_2245),
.Y(n_2588)
);

OAI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2125),
.A2(n_2224),
.B1(n_2238),
.B2(n_2202),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2264),
.Y(n_2590)
);

AOI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2352),
.A2(n_2392),
.B1(n_2384),
.B2(n_2202),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2214),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_SL g2593 ( 
.A1(n_2138),
.A2(n_2384),
.B1(n_2153),
.B2(n_2216),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2338),
.Y(n_2594)
);

INVx2_ASAP7_75t_SL g2595 ( 
.A(n_2187),
.Y(n_2595)
);

AOI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_2352),
.A2(n_2392),
.B1(n_2354),
.B2(n_2356),
.Y(n_2596)
);

NAND2x1p5_ASAP7_75t_L g2597 ( 
.A(n_2270),
.B(n_2230),
.Y(n_2597)
);

OA21x2_ASAP7_75t_L g2598 ( 
.A1(n_2142),
.A2(n_2366),
.B(n_2206),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2190),
.Y(n_2599)
);

NAND2x1p5_ASAP7_75t_L g2600 ( 
.A(n_2190),
.B(n_2209),
.Y(n_2600)
);

INVxp67_ASAP7_75t_SL g2601 ( 
.A(n_2359),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2430),
.B(n_2311),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2421),
.Y(n_2603)
);

CKINVDCx16_ASAP7_75t_R g2604 ( 
.A(n_2419),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2459),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2431),
.B(n_2396),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2410),
.Y(n_2607)
);

OR2x6_ASAP7_75t_L g2608 ( 
.A(n_2507),
.B(n_2326),
.Y(n_2608)
);

O2A1O1Ixp33_ASAP7_75t_L g2609 ( 
.A1(n_2563),
.A2(n_2357),
.B(n_2315),
.C(n_2320),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2463),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_R g2611 ( 
.A(n_2427),
.B(n_2341),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2533),
.B(n_2186),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2488),
.B(n_2396),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_2504),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2412),
.Y(n_2615)
);

OR2x6_ASAP7_75t_L g2616 ( 
.A(n_2588),
.B(n_2493),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_R g2617 ( 
.A(n_2451),
.B(n_2480),
.Y(n_2617)
);

AOI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2503),
.A2(n_2224),
.B1(n_2299),
.B2(n_2304),
.C(n_2319),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2416),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2498),
.Y(n_2620)
);

AND2x4_ASAP7_75t_L g2621 ( 
.A(n_2434),
.B(n_2240),
.Y(n_2621)
);

AND2x4_ASAP7_75t_L g2622 ( 
.A(n_2434),
.B(n_2240),
.Y(n_2622)
);

OAI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2439),
.A2(n_2187),
.B1(n_2317),
.B2(n_2365),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_L g2624 ( 
.A1(n_2552),
.A2(n_2382),
.B1(n_2360),
.B2(n_2322),
.Y(n_2624)
);

NAND2x1_ASAP7_75t_L g2625 ( 
.A(n_2515),
.B(n_2359),
.Y(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2552),
.A2(n_2382),
.B1(n_2360),
.B2(n_2322),
.Y(n_2626)
);

BUFx4f_ASAP7_75t_L g2627 ( 
.A(n_2478),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2429),
.B(n_2318),
.Y(n_2628)
);

CKINVDCx16_ASAP7_75t_R g2629 ( 
.A(n_2569),
.Y(n_2629)
);

AND2x4_ASAP7_75t_L g2630 ( 
.A(n_2434),
.B(n_2452),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2418),
.B(n_2318),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2524),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2516),
.B(n_2490),
.Y(n_2633)
);

OR2x2_ASAP7_75t_L g2634 ( 
.A(n_2442),
.B(n_2148),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2530),
.Y(n_2635)
);

AO31x2_ASAP7_75t_L g2636 ( 
.A1(n_2560),
.A2(n_2234),
.A3(n_2158),
.B(n_2273),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2424),
.Y(n_2637)
);

NAND3xp33_ASAP7_75t_L g2638 ( 
.A(n_2495),
.B(n_2332),
.C(n_2348),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2471),
.Y(n_2639)
);

O2A1O1Ixp33_ASAP7_75t_L g2640 ( 
.A1(n_2579),
.A2(n_2331),
.B(n_2317),
.C(n_2348),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_R g2641 ( 
.A(n_2438),
.B(n_2148),
.Y(n_2641)
);

NOR3xp33_ASAP7_75t_SL g2642 ( 
.A(n_2496),
.B(n_2313),
.C(n_2196),
.Y(n_2642)
);

NAND2xp33_ASAP7_75t_R g2643 ( 
.A(n_2501),
.B(n_2177),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2509),
.B(n_2177),
.Y(n_2644)
);

INVxp67_ASAP7_75t_L g2645 ( 
.A(n_2556),
.Y(n_2645)
);

AO32x2_ASAP7_75t_L g2646 ( 
.A1(n_2436),
.A2(n_2369),
.A3(n_2154),
.B1(n_2365),
.B2(n_2343),
.Y(n_2646)
);

OR2x6_ASAP7_75t_L g2647 ( 
.A(n_2411),
.B(n_2225),
.Y(n_2647)
);

INVx2_ASAP7_75t_SL g2648 ( 
.A(n_2504),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2495),
.A2(n_2564),
.B1(n_2589),
.B2(n_2435),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2425),
.B(n_2329),
.Y(n_2650)
);

OR2x6_ASAP7_75t_L g2651 ( 
.A(n_2422),
.B(n_2231),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2437),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2594),
.B(n_2134),
.Y(n_2653)
);

AND2x2_ASAP7_75t_SL g2654 ( 
.A(n_2422),
.B(n_2368),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2587),
.Y(n_2655)
);

OAI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2589),
.A2(n_2383),
.B(n_2593),
.Y(n_2656)
);

AND2x6_ASAP7_75t_L g2657 ( 
.A(n_2523),
.B(n_2368),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2453),
.A2(n_2134),
.B1(n_2164),
.B2(n_2289),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2464),
.A2(n_2164),
.B1(n_2236),
.B2(n_2289),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_R g2660 ( 
.A(n_2542),
.B(n_2231),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2510),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2444),
.B(n_2329),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2413),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2446),
.B(n_2154),
.Y(n_2664)
);

OAI21xp5_ASAP7_75t_SL g2665 ( 
.A1(n_2454),
.A2(n_2296),
.B(n_2368),
.Y(n_2665)
);

NOR3xp33_ASAP7_75t_SL g2666 ( 
.A(n_2462),
.B(n_2122),
.C(n_2200),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_2549),
.Y(n_2667)
);

OAI21xp5_ASAP7_75t_SL g2668 ( 
.A1(n_2454),
.A2(n_2397),
.B(n_2236),
.Y(n_2668)
);

CKINVDCx20_ASAP7_75t_R g2669 ( 
.A(n_2547),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2485),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2529),
.B(n_2173),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2448),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2554),
.B(n_2173),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2441),
.B(n_2169),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2441),
.B(n_2141),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_2485),
.Y(n_2676)
);

CKINVDCx8_ASAP7_75t_R g2677 ( 
.A(n_2557),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2450),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2447),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2447),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2456),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2456),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2420),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2457),
.Y(n_2684)
);

BUFx6f_ASAP7_75t_L g2685 ( 
.A(n_2510),
.Y(n_2685)
);

AND2x2_ASAP7_75t_SL g2686 ( 
.A(n_2585),
.B(n_2240),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2452),
.B(n_2141),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2458),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2460),
.B(n_2336),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2567),
.B(n_2192),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_R g2691 ( 
.A(n_2497),
.B(n_2169),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2468),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2469),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_2491),
.Y(n_2694)
);

OR2x2_ASAP7_75t_L g2695 ( 
.A(n_2492),
.B(n_2122),
.Y(n_2695)
);

BUFx4f_ASAP7_75t_SL g2696 ( 
.A(n_2585),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2592),
.B(n_2185),
.Y(n_2697)
);

CKINVDCx11_ASAP7_75t_R g2698 ( 
.A(n_2555),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2470),
.B(n_2379),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2473),
.B(n_2379),
.Y(n_2700)
);

NAND2xp33_ASAP7_75t_SL g2701 ( 
.A(n_2582),
.B(n_2540),
.Y(n_2701)
);

INVxp67_ASAP7_75t_L g2702 ( 
.A(n_2449),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2494),
.B(n_2185),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_2482),
.B(n_2136),
.Y(n_2704)
);

CKINVDCx16_ASAP7_75t_R g2705 ( 
.A(n_2555),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2483),
.Y(n_2706)
);

BUFx8_ASAP7_75t_SL g2707 ( 
.A(n_2415),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2486),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2491),
.B(n_2389),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2531),
.Y(n_2710)
);

INVx3_ASAP7_75t_L g2711 ( 
.A(n_2499),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_R g2712 ( 
.A(n_2548),
.B(n_2136),
.Y(n_2712)
);

NAND2xp33_ASAP7_75t_SL g2713 ( 
.A(n_2540),
.B(n_2136),
.Y(n_2713)
);

CKINVDCx14_ASAP7_75t_R g2714 ( 
.A(n_2545),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_2565),
.Y(n_2715)
);

HB1xp67_ASAP7_75t_L g2716 ( 
.A(n_2414),
.Y(n_2716)
);

XNOR2xp5_ASAP7_75t_L g2717 ( 
.A(n_2472),
.B(n_2241),
.Y(n_2717)
);

CKINVDCx16_ASAP7_75t_R g2718 ( 
.A(n_2461),
.Y(n_2718)
);

NAND4xp25_ASAP7_75t_SL g2719 ( 
.A(n_2465),
.B(n_2553),
.C(n_2475),
.D(n_2535),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2467),
.B(n_2207),
.Y(n_2720)
);

O2A1O1Ixp33_ASAP7_75t_L g2721 ( 
.A1(n_2520),
.A2(n_2342),
.B(n_2193),
.C(n_2233),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2466),
.Y(n_2722)
);

AND2x4_ASAP7_75t_L g2723 ( 
.A(n_2428),
.B(n_2192),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2522),
.Y(n_2724)
);

O2A1O1Ixp33_ASAP7_75t_SL g2725 ( 
.A1(n_2474),
.A2(n_2207),
.B(n_2206),
.C(n_2219),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2512),
.B(n_2517),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2532),
.Y(n_2727)
);

INVxp67_ASAP7_75t_L g2728 ( 
.A(n_2561),
.Y(n_2728)
);

AO31x2_ASAP7_75t_L g2729 ( 
.A1(n_2580),
.A2(n_2193),
.A3(n_2233),
.B(n_2220),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2566),
.B(n_2180),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2545),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2466),
.B(n_2235),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_2461),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2536),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2512),
.B(n_2342),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2538),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2570),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_R g2738 ( 
.A(n_2548),
.B(n_2192),
.Y(n_2738)
);

OAI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2489),
.A2(n_2192),
.B1(n_2178),
.B2(n_2184),
.Y(n_2739)
);

NOR3xp33_ASAP7_75t_SL g2740 ( 
.A(n_2572),
.B(n_2191),
.C(n_2161),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_2570),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2481),
.B(n_2514),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2499),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2500),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2432),
.B(n_2334),
.Y(n_2745)
);

AOI21xp33_ASAP7_75t_L g2746 ( 
.A1(n_2591),
.A2(n_2281),
.B(n_2184),
.Y(n_2746)
);

NAND2xp33_ASAP7_75t_R g2747 ( 
.A(n_2428),
.B(n_2440),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2455),
.B(n_2481),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2500),
.Y(n_2749)
);

NAND3xp33_ASAP7_75t_SL g2750 ( 
.A(n_2575),
.B(n_2178),
.C(n_2184),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2514),
.B(n_2178),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2527),
.B(n_2188),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2455),
.B(n_2188),
.Y(n_2753)
);

O2A1O1Ixp33_ASAP7_75t_SL g2754 ( 
.A1(n_2551),
.A2(n_2188),
.B(n_2279),
.C(n_2297),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2440),
.B(n_2306),
.Y(n_2755)
);

INVx5_ASAP7_75t_L g2756 ( 
.A(n_2525),
.Y(n_2756)
);

NAND2xp33_ASAP7_75t_SL g2757 ( 
.A(n_2525),
.B(n_2306),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2595),
.B(n_2306),
.Y(n_2758)
);

CKINVDCx16_ASAP7_75t_R g2759 ( 
.A(n_2578),
.Y(n_2759)
);

OR2x6_ASAP7_75t_L g2760 ( 
.A(n_2600),
.B(n_2597),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2543),
.Y(n_2761)
);

OAI21xp33_ASAP7_75t_L g2762 ( 
.A1(n_2423),
.A2(n_2586),
.B(n_2596),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2559),
.Y(n_2763)
);

HB1xp67_ASAP7_75t_L g2764 ( 
.A(n_2681),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2607),
.Y(n_2765)
);

OAI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2616),
.A2(n_2558),
.B1(n_2511),
.B2(n_2417),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2615),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2619),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2620),
.B(n_2633),
.Y(n_2769)
);

INVx2_ASAP7_75t_R g2770 ( 
.A(n_2756),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2663),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2637),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2716),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2699),
.B(n_2546),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2683),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2652),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2700),
.B(n_2546),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2672),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2710),
.B(n_2706),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2602),
.B(n_2583),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2708),
.B(n_2568),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2689),
.B(n_2537),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2678),
.Y(n_2783)
);

HB1xp67_ASAP7_75t_L g2784 ( 
.A(n_2722),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2720),
.B(n_2624),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2626),
.B(n_2476),
.Y(n_2786)
);

OR2x2_ASAP7_75t_L g2787 ( 
.A(n_2605),
.B(n_2484),
.Y(n_2787)
);

CKINVDCx16_ASAP7_75t_R g2788 ( 
.A(n_2604),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2684),
.B(n_2476),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2688),
.B(n_2692),
.Y(n_2790)
);

AND2x4_ASAP7_75t_SL g2791 ( 
.A(n_2616),
.B(n_2523),
.Y(n_2791)
);

INVxp33_ASAP7_75t_L g2792 ( 
.A(n_2712),
.Y(n_2792)
);

BUFx6f_ASAP7_75t_L g2793 ( 
.A(n_2682),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2693),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2606),
.B(n_2735),
.Y(n_2795)
);

INVx3_ASAP7_75t_L g2796 ( 
.A(n_2723),
.Y(n_2796)
);

NOR2x1_ASAP7_75t_L g2797 ( 
.A(n_2608),
.B(n_2647),
.Y(n_2797)
);

BUFx6f_ASAP7_75t_L g2798 ( 
.A(n_2686),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2745),
.B(n_2423),
.Y(n_2799)
);

AND2x2_ASAP7_75t_SL g2800 ( 
.A(n_2654),
.B(n_2515),
.Y(n_2800)
);

OR2x2_ASAP7_75t_L g2801 ( 
.A(n_2759),
.B(n_2484),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2726),
.B(n_2599),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2603),
.Y(n_2803)
);

BUFx3_ASAP7_75t_L g2804 ( 
.A(n_2696),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2742),
.B(n_2518),
.Y(n_2805)
);

INVx3_ASAP7_75t_L g2806 ( 
.A(n_2755),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2747),
.Y(n_2807)
);

BUFx2_ASAP7_75t_L g2808 ( 
.A(n_2641),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2730),
.B(n_2613),
.Y(n_2809)
);

INVxp67_ASAP7_75t_L g2810 ( 
.A(n_2651),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2724),
.B(n_2727),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2651),
.Y(n_2812)
);

CKINVDCx14_ASAP7_75t_R g2813 ( 
.A(n_2617),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2734),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2736),
.Y(n_2815)
);

INVx3_ASAP7_75t_L g2816 ( 
.A(n_2755),
.Y(n_2816)
);

OR2x2_ASAP7_75t_L g2817 ( 
.A(n_2748),
.B(n_2550),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2761),
.B(n_2433),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2753),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2664),
.B(n_2502),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2732),
.B(n_2508),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2653),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2646),
.B(n_2513),
.Y(n_2823)
);

AND2x4_ASAP7_75t_L g2824 ( 
.A(n_2751),
.B(n_2709),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2695),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2666),
.B(n_2656),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2625),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2645),
.B(n_2562),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2634),
.B(n_2559),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2703),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2657),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2631),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2650),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2662),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2704),
.Y(n_2835)
);

NOR2x1p5_ASAP7_75t_L g2836 ( 
.A(n_2679),
.B(n_2590),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2636),
.B(n_2573),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2762),
.B(n_2574),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2612),
.B(n_2541),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2649),
.B(n_2477),
.Y(n_2840)
);

INVxp67_ASAP7_75t_L g2841 ( 
.A(n_2647),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2618),
.A2(n_2581),
.B1(n_2426),
.B2(n_2584),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2763),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2697),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2715),
.Y(n_2845)
);

BUFx2_ASAP7_75t_L g2846 ( 
.A(n_2608),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2657),
.Y(n_2847)
);

BUFx2_ASAP7_75t_SL g2848 ( 
.A(n_2677),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2752),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2729),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2657),
.Y(n_2851)
);

BUFx2_ASAP7_75t_L g2852 ( 
.A(n_2738),
.Y(n_2852)
);

NOR3xp33_ASAP7_75t_L g2853 ( 
.A(n_2797),
.B(n_2638),
.C(n_2609),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2809),
.B(n_2746),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2789),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2764),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2830),
.B(n_2628),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2809),
.B(n_2729),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2795),
.B(n_2729),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2790),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2789),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2790),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2765),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2767),
.Y(n_2864)
);

OR2x2_ASAP7_75t_L g2865 ( 
.A(n_2769),
.B(n_2629),
.Y(n_2865)
);

NAND3xp33_ASAP7_75t_L g2866 ( 
.A(n_2842),
.B(n_2784),
.C(n_2773),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2768),
.Y(n_2867)
);

INVxp67_ASAP7_75t_SL g2868 ( 
.A(n_2801),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2818),
.Y(n_2869)
);

NAND3xp33_ASAP7_75t_L g2870 ( 
.A(n_2842),
.B(n_2740),
.C(n_2521),
.Y(n_2870)
);

OR2x2_ASAP7_75t_L g2871 ( 
.A(n_2825),
.B(n_2705),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2795),
.B(n_2598),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2772),
.Y(n_2873)
);

HB1xp67_ASAP7_75t_L g2874 ( 
.A(n_2771),
.Y(n_2874)
);

OR2x2_ASAP7_75t_L g2875 ( 
.A(n_2825),
.B(n_2702),
.Y(n_2875)
);

OR2x2_ASAP7_75t_L g2876 ( 
.A(n_2849),
.B(n_2719),
.Y(n_2876)
);

AND2x4_ASAP7_75t_SL g2877 ( 
.A(n_2798),
.B(n_2630),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2821),
.B(n_2598),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2776),
.Y(n_2879)
);

NAND3xp33_ASAP7_75t_L g2880 ( 
.A(n_2826),
.B(n_2668),
.C(n_2539),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2818),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_R g2882 ( 
.A(n_2813),
.B(n_2718),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2778),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2799),
.B(n_2576),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2783),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2799),
.B(n_2534),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2771),
.Y(n_2887)
);

OR2x2_ASAP7_75t_L g2888 ( 
.A(n_2805),
.B(n_2644),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2794),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2814),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2774),
.B(n_2721),
.Y(n_2891)
);

OR2x2_ASAP7_75t_L g2892 ( 
.A(n_2805),
.B(n_2648),
.Y(n_2892)
);

OR2x2_ASAP7_75t_L g2893 ( 
.A(n_2787),
.B(n_2728),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2802),
.B(n_2717),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2774),
.B(n_2544),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2802),
.B(n_2623),
.Y(n_2896)
);

AND2x4_ASAP7_75t_L g2897 ( 
.A(n_2824),
.B(n_2690),
.Y(n_2897)
);

OR2x2_ASAP7_75t_L g2898 ( 
.A(n_2844),
.B(n_2630),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2815),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2811),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2775),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2803),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2779),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2832),
.B(n_2671),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2833),
.B(n_2673),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2777),
.B(n_2511),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2777),
.B(n_2443),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2858),
.B(n_2785),
.Y(n_2908)
);

HB1xp67_ASAP7_75t_L g2909 ( 
.A(n_2856),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2877),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2858),
.B(n_2822),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2872),
.B(n_2785),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2872),
.B(n_2782),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_2877),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2874),
.Y(n_2915)
);

AND2x4_ASAP7_75t_L g2916 ( 
.A(n_2897),
.B(n_2824),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2874),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2855),
.B(n_2819),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2886),
.B(n_2782),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2901),
.Y(n_2920)
);

AOI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2853),
.A2(n_2826),
.B1(n_2840),
.B2(n_2766),
.Y(n_2921)
);

AND2x2_ASAP7_75t_L g2922 ( 
.A(n_2886),
.B(n_2786),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2856),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2859),
.B(n_2834),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2869),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2901),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2854),
.B(n_2786),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2859),
.B(n_2835),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2854),
.B(n_2823),
.Y(n_2929)
);

HB1xp67_ASAP7_75t_L g2930 ( 
.A(n_2888),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2865),
.B(n_2788),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2869),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2900),
.B(n_2813),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2860),
.B(n_2820),
.Y(n_2934)
);

INVxp67_ASAP7_75t_L g2935 ( 
.A(n_2868),
.Y(n_2935)
);

INVx1_ASAP7_75t_SL g2936 ( 
.A(n_2882),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2907),
.B(n_2823),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2862),
.B(n_2820),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2903),
.B(n_2838),
.Y(n_2939)
);

INVx2_ASAP7_75t_SL g2940 ( 
.A(n_2882),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2861),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2907),
.B(n_2824),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2881),
.B(n_2857),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2878),
.B(n_2837),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2878),
.B(n_2837),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2861),
.B(n_2843),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2887),
.Y(n_2947)
);

AND2x4_ASAP7_75t_L g2948 ( 
.A(n_2897),
.B(n_2807),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2902),
.B(n_2838),
.Y(n_2949)
);

HB1xp67_ASAP7_75t_L g2950 ( 
.A(n_2892),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2887),
.Y(n_2951)
);

OR2x2_ASAP7_75t_L g2952 ( 
.A(n_2875),
.B(n_2817),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2921),
.A2(n_2880),
.B1(n_2826),
.B2(n_2876),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2919),
.B(n_2897),
.Y(n_2954)
);

HB1xp67_ASAP7_75t_L g2955 ( 
.A(n_2923),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2908),
.B(n_2891),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2909),
.Y(n_2957)
);

OAI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2940),
.A2(n_2896),
.B1(n_2798),
.B2(n_2866),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2919),
.B(n_2884),
.Y(n_2959)
);

A2O1A1Ixp33_ASAP7_75t_L g2960 ( 
.A1(n_2940),
.A2(n_2808),
.B(n_2846),
.C(n_2791),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2925),
.Y(n_2961)
);

NAND2x1p5_ASAP7_75t_L g2962 ( 
.A(n_2936),
.B(n_2804),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2925),
.Y(n_2963)
);

HB1xp67_ASAP7_75t_L g2964 ( 
.A(n_2923),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2908),
.A2(n_2876),
.B1(n_2870),
.B2(n_2894),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2912),
.B(n_2891),
.Y(n_2966)
);

NAND3xp33_ASAP7_75t_L g2967 ( 
.A(n_2935),
.B(n_2845),
.C(n_2871),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2939),
.A2(n_2927),
.B1(n_2948),
.B2(n_2922),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2930),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2942),
.B(n_2884),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2952),
.Y(n_2971)
);

XNOR2x2_ASAP7_75t_L g2972 ( 
.A(n_2933),
.B(n_2893),
.Y(n_2972)
);

OAI31xp33_ASAP7_75t_L g2973 ( 
.A1(n_2931),
.A2(n_2804),
.A3(n_2791),
.B(n_2836),
.Y(n_2973)
);

OR2x6_ASAP7_75t_L g2974 ( 
.A(n_2910),
.B(n_2848),
.Y(n_2974)
);

A2O1A1Ixp33_ASAP7_75t_L g2975 ( 
.A1(n_2948),
.A2(n_2812),
.B(n_2841),
.C(n_2640),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2912),
.B(n_2895),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2952),
.Y(n_2977)
);

OA222x2_ASAP7_75t_L g2978 ( 
.A1(n_2946),
.A2(n_2812),
.B1(n_2851),
.B2(n_2831),
.C1(n_2898),
.C2(n_2810),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2947),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2932),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2947),
.Y(n_2981)
);

XNOR2xp5_ASAP7_75t_L g2982 ( 
.A(n_2950),
.B(n_2655),
.Y(n_2982)
);

INVx2_ASAP7_75t_SL g2983 ( 
.A(n_2946),
.Y(n_2983)
);

HB1xp67_ASAP7_75t_L g2984 ( 
.A(n_2915),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2942),
.B(n_2913),
.Y(n_2985)
);

OAI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2910),
.A2(n_2798),
.B1(n_2792),
.B2(n_2793),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2951),
.Y(n_2987)
);

INVxp67_ASAP7_75t_L g2988 ( 
.A(n_2915),
.Y(n_2988)
);

AND2x2_ASAP7_75t_SL g2989 ( 
.A(n_2948),
.B(n_2800),
.Y(n_2989)
);

INVx1_ASAP7_75t_SL g2990 ( 
.A(n_2914),
.Y(n_2990)
);

INVx2_ASAP7_75t_SL g2991 ( 
.A(n_2914),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2949),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2913),
.B(n_2895),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2943),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2957),
.Y(n_2995)
);

INVxp67_ASAP7_75t_SL g2996 ( 
.A(n_2955),
.Y(n_2996)
);

NAND3xp33_ASAP7_75t_SL g2997 ( 
.A(n_2975),
.B(n_2680),
.C(n_2669),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2961),
.Y(n_2998)
);

NAND4xp75_ASAP7_75t_L g2999 ( 
.A(n_2973),
.B(n_2642),
.C(n_2800),
.D(n_2927),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2969),
.Y(n_3000)
);

A2O1A1Ixp33_ASAP7_75t_L g3001 ( 
.A1(n_2960),
.A2(n_2627),
.B(n_2670),
.C(n_2676),
.Y(n_3001)
);

NAND2x1p5_ASAP7_75t_L g3002 ( 
.A(n_2989),
.B(n_2793),
.Y(n_3002)
);

OAI21xp5_ASAP7_75t_L g3003 ( 
.A1(n_2960),
.A2(n_2975),
.B(n_2953),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2974),
.A2(n_2916),
.B1(n_2924),
.B2(n_2798),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2989),
.A2(n_2713),
.B(n_2916),
.Y(n_3005)
);

HB1xp67_ASAP7_75t_L g3006 ( 
.A(n_2955),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2971),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2978),
.B(n_2922),
.Y(n_3008)
);

INVxp67_ASAP7_75t_L g3009 ( 
.A(n_2974),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2977),
.Y(n_3010)
);

AOI22xp33_ASAP7_75t_L g3011 ( 
.A1(n_2972),
.A2(n_2965),
.B1(n_2974),
.B2(n_2967),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2994),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2984),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2984),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2992),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2964),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2964),
.Y(n_3017)
);

INVx3_ASAP7_75t_L g3018 ( 
.A(n_2962),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2988),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2988),
.Y(n_3020)
);

INVxp67_ASAP7_75t_SL g3021 ( 
.A(n_2962),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_3006),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_3009),
.B(n_2954),
.Y(n_3023)
);

OAI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_3001),
.A2(n_2958),
.B(n_2982),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2997),
.A2(n_2958),
.B1(n_2990),
.B2(n_2991),
.Y(n_3025)
);

NOR2x1_ASAP7_75t_L g3026 ( 
.A(n_3001),
.B(n_2986),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_3012),
.B(n_2993),
.Y(n_3027)
);

NOR2x1_ASAP7_75t_L g3028 ( 
.A(n_3018),
.B(n_2986),
.Y(n_3028)
);

AOI211xp5_ASAP7_75t_L g3029 ( 
.A1(n_3003),
.A2(n_2667),
.B(n_2733),
.C(n_2610),
.Y(n_3029)
);

OAI221xp5_ASAP7_75t_L g3030 ( 
.A1(n_3011),
.A2(n_2968),
.B1(n_2956),
.B2(n_2966),
.C(n_2983),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_3021),
.B(n_2985),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_3006),
.Y(n_3032)
);

AOI211x1_ASAP7_75t_L g3033 ( 
.A1(n_3008),
.A2(n_2976),
.B(n_2929),
.C(n_2937),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_3015),
.B(n_2929),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2995),
.B(n_2959),
.Y(n_3035)
);

AOI211xp5_ASAP7_75t_L g3036 ( 
.A1(n_3004),
.A2(n_2632),
.B(n_2792),
.C(n_2793),
.Y(n_3036)
);

AOI221xp5_ASAP7_75t_L g3037 ( 
.A1(n_3011),
.A2(n_2911),
.B1(n_2885),
.B2(n_2883),
.C(n_2879),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_3018),
.B(n_2793),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_3000),
.B(n_2944),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_3019),
.B(n_2944),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_3020),
.Y(n_3041)
);

AOI211xp5_ASAP7_75t_L g3042 ( 
.A1(n_3005),
.A2(n_2665),
.B(n_2694),
.C(n_2611),
.Y(n_3042)
);

NOR2x1_ASAP7_75t_L g3043 ( 
.A(n_3018),
.B(n_2614),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2999),
.A2(n_2916),
.B1(n_2906),
.B2(n_2905),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_3020),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2996),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_3016),
.Y(n_3047)
);

AOI221xp5_ASAP7_75t_L g3048 ( 
.A1(n_3017),
.A2(n_2873),
.B1(n_2889),
.B2(n_2890),
.C(n_2863),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_3002),
.B(n_2970),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_3046),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_3022),
.Y(n_3051)
);

NAND3xp33_ASAP7_75t_SL g3052 ( 
.A(n_3024),
.B(n_3002),
.C(n_2660),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_3030),
.B(n_3007),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_3031),
.Y(n_3054)
);

INVx3_ASAP7_75t_L g3055 ( 
.A(n_3023),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_3026),
.B(n_3013),
.Y(n_3056)
);

OR2x2_ASAP7_75t_L g3057 ( 
.A(n_3034),
.B(n_3014),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_SL g3058 ( 
.A(n_3043),
.B(n_2635),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_3037),
.B(n_3010),
.Y(n_3059)
);

NAND2x1_ASAP7_75t_L g3060 ( 
.A(n_3028),
.B(n_2998),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_3032),
.Y(n_3061)
);

XNOR2xp5_ASAP7_75t_L g3062 ( 
.A(n_3029),
.B(n_2639),
.Y(n_3062)
);

OAI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_3024),
.A2(n_2714),
.B(n_2998),
.Y(n_3063)
);

NOR3x1_ASAP7_75t_L g3064 ( 
.A(n_3041),
.B(n_2487),
.C(n_2847),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_3034),
.B(n_3045),
.Y(n_3065)
);

OAI21xp5_ASAP7_75t_SL g3066 ( 
.A1(n_3025),
.A2(n_2852),
.B(n_2851),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_3038),
.A2(n_2741),
.B(n_2737),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_3036),
.B(n_2961),
.Y(n_3068)
);

OR2x2_ASAP7_75t_L g3069 ( 
.A(n_3047),
.B(n_2928),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3035),
.Y(n_3070)
);

AOI211xp5_ASAP7_75t_L g3071 ( 
.A1(n_3052),
.A2(n_3042),
.B(n_3044),
.C(n_3049),
.Y(n_3071)
);

OAI211xp5_ASAP7_75t_SL g3072 ( 
.A1(n_3063),
.A2(n_2698),
.B(n_3048),
.C(n_3040),
.Y(n_3072)
);

AOI22x1_ASAP7_75t_L g3073 ( 
.A1(n_3056),
.A2(n_2743),
.B1(n_2744),
.B2(n_2749),
.Y(n_3073)
);

NOR2x1_ASAP7_75t_L g3074 ( 
.A(n_3060),
.B(n_3062),
.Y(n_3074)
);

NAND3xp33_ASAP7_75t_L g3075 ( 
.A(n_3050),
.B(n_3033),
.C(n_3027),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_3058),
.A2(n_3039),
.B(n_2757),
.Y(n_3076)
);

AOI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_3066),
.A2(n_2828),
.B(n_2701),
.Y(n_3077)
);

OAI211xp5_ASAP7_75t_SL g3078 ( 
.A1(n_3055),
.A2(n_2711),
.B(n_2904),
.C(n_2675),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3054),
.Y(n_3079)
);

AO22x1_ASAP7_75t_L g3080 ( 
.A1(n_3064),
.A2(n_2756),
.B1(n_2621),
.B2(n_2622),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_3067),
.A2(n_2760),
.B(n_2725),
.Y(n_3081)
);

AO22x2_ASAP7_75t_L g3082 ( 
.A1(n_3051),
.A2(n_3061),
.B1(n_3055),
.B2(n_3070),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_3053),
.A2(n_2760),
.B(n_2963),
.Y(n_3083)
);

NOR2x1_ASAP7_75t_SL g3084 ( 
.A(n_3068),
.B(n_2661),
.Y(n_3084)
);

NOR2x1_ASAP7_75t_L g3085 ( 
.A(n_3059),
.B(n_2661),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_3064),
.B(n_2937),
.Y(n_3086)
);

AND4x1_ASAP7_75t_L g3087 ( 
.A(n_3065),
.B(n_2707),
.C(n_2643),
.D(n_2691),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_3079),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3082),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_3082),
.B(n_3057),
.Y(n_3090)
);

NAND4xp75_ASAP7_75t_L g3091 ( 
.A(n_3074),
.B(n_2840),
.C(n_2945),
.D(n_2906),
.Y(n_3091)
);

OAI21x1_ASAP7_75t_SL g3092 ( 
.A1(n_3084),
.A2(n_3069),
.B(n_2526),
.Y(n_3092)
);

NAND4xp25_ASAP7_75t_L g3093 ( 
.A(n_3071),
.B(n_2621),
.C(n_2622),
.D(n_2831),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_3086),
.B(n_2945),
.Y(n_3094)
);

NAND4xp75_ASAP7_75t_L g3095 ( 
.A(n_3085),
.B(n_2920),
.C(n_2926),
.D(n_2917),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_3076),
.A2(n_2731),
.B(n_2658),
.Y(n_3096)
);

OAI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_3083),
.A2(n_3075),
.B(n_3077),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_3073),
.A2(n_2731),
.B(n_2659),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_3072),
.A2(n_2980),
.B(n_2963),
.Y(n_3099)
);

OAI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_3081),
.A2(n_2519),
.B(n_2739),
.Y(n_3100)
);

OAI221xp5_ASAP7_75t_SL g3101 ( 
.A1(n_3087),
.A2(n_2851),
.B1(n_2831),
.B2(n_2839),
.C(n_2829),
.Y(n_3101)
);

OAI21xp5_ASAP7_75t_SL g3102 ( 
.A1(n_3078),
.A2(n_2685),
.B(n_2528),
.Y(n_3102)
);

OAI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_3091),
.A2(n_3080),
.B1(n_2980),
.B2(n_2926),
.Y(n_3103)
);

INVxp33_ASAP7_75t_L g3104 ( 
.A(n_3088),
.Y(n_3104)
);

NOR2x1p5_ASAP7_75t_L g3105 ( 
.A(n_3093),
.B(n_2685),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_3089),
.Y(n_3106)
);

AO211x2_ASAP7_75t_L g3107 ( 
.A1(n_3097),
.A2(n_2920),
.B(n_2917),
.C(n_2899),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_3093),
.A2(n_2867),
.B1(n_2864),
.B2(n_2938),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3090),
.B(n_3094),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3096),
.Y(n_3110)
);

INVx2_ASAP7_75t_SL g3111 ( 
.A(n_3092),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_3098),
.A2(n_2934),
.B1(n_2519),
.B2(n_2979),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_3095),
.Y(n_3113)
);

OR2x2_ASAP7_75t_L g3114 ( 
.A(n_3099),
.B(n_3101),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_3105),
.Y(n_3115)
);

NOR2x1p5_ASAP7_75t_L g3116 ( 
.A(n_3110),
.B(n_3102),
.Y(n_3116)
);

NAND3xp33_ASAP7_75t_SL g3117 ( 
.A(n_3106),
.B(n_3100),
.C(n_2600),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_3112),
.B(n_2981),
.Y(n_3118)
);

AOI221xp5_ASAP7_75t_L g3119 ( 
.A1(n_3104),
.A2(n_2987),
.B1(n_2781),
.B2(n_2941),
.C(n_2506),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_3114),
.B(n_2827),
.Y(n_3120)
);

AOI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_3109),
.A2(n_2756),
.B1(n_2827),
.B2(n_2687),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_3111),
.Y(n_3122)
);

INVx2_ASAP7_75t_SL g3123 ( 
.A(n_3113),
.Y(n_3123)
);

INVx1_ASAP7_75t_SL g3124 ( 
.A(n_3108),
.Y(n_3124)
);

NOR3xp33_ASAP7_75t_L g3125 ( 
.A(n_3103),
.B(n_2750),
.C(n_2590),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_3107),
.A2(n_2674),
.B(n_2597),
.Y(n_3126)
);

NOR3x1_ASAP7_75t_L g3127 ( 
.A(n_3111),
.B(n_2941),
.C(n_2918),
.Y(n_3127)
);

HB1xp67_ASAP7_75t_L g3128 ( 
.A(n_3123),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_3122),
.Y(n_3129)
);

NOR2xp67_ASAP7_75t_L g3130 ( 
.A(n_3115),
.B(n_2827),
.Y(n_3130)
);

BUFx12f_ASAP7_75t_L g3131 ( 
.A(n_3116),
.Y(n_3131)
);

NOR4xp25_ASAP7_75t_SL g3132 ( 
.A(n_3119),
.B(n_2754),
.C(n_2770),
.D(n_2601),
.Y(n_3132)
);

BUFx2_ASAP7_75t_L g3133 ( 
.A(n_3121),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_3124),
.Y(n_3134)
);

AOI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_3129),
.A2(n_3120),
.B1(n_3117),
.B2(n_3125),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3128),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_3131),
.A2(n_3118),
.B1(n_3126),
.B2(n_3127),
.Y(n_3137)
);

INVxp67_ASAP7_75t_SL g3138 ( 
.A(n_3128),
.Y(n_3138)
);

INVxp67_ASAP7_75t_L g3139 ( 
.A(n_3134),
.Y(n_3139)
);

AOI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_3139),
.A2(n_3133),
.B1(n_3130),
.B2(n_3132),
.Y(n_3140)
);

AOI22xp5_ASAP7_75t_L g3141 ( 
.A1(n_3138),
.A2(n_2479),
.B1(n_2505),
.B2(n_2528),
.Y(n_3141)
);

NOR2xp67_ASAP7_75t_L g3142 ( 
.A(n_3136),
.B(n_3137),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_3135),
.B(n_2850),
.Y(n_3143)
);

INVx4_ASAP7_75t_L g3144 ( 
.A(n_3136),
.Y(n_3144)
);

CKINVDCx5p33_ASAP7_75t_R g3145 ( 
.A(n_3144),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_3140),
.A2(n_2505),
.B1(n_2479),
.B2(n_2445),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_3142),
.B(n_2780),
.Y(n_3147)
);

OAI222xp33_ASAP7_75t_L g3148 ( 
.A1(n_3145),
.A2(n_3143),
.B1(n_3141),
.B2(n_2445),
.C1(n_2506),
.C2(n_2577),
.Y(n_3148)
);

OAI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_3148),
.A2(n_3147),
.B(n_3146),
.Y(n_3149)
);

AOI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_3149),
.A2(n_2571),
.B1(n_2687),
.B2(n_2758),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_3150),
.B(n_2770),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_3151),
.A2(n_2816),
.B1(n_2796),
.B2(n_2806),
.Y(n_3152)
);


endmodule