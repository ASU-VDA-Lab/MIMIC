module fake_jpeg_18636_n_65 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_24),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_38),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_4),
.B(n_6),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_47),
.B(n_49),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_8),
.B2(n_10),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_7),
.B(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_53),
.B(n_50),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_56),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_21),
.Y(n_65)
);


endmodule