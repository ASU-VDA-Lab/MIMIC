module fake_netlist_6_20_n_1899 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1899);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1899;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_18),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_91),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_0),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_17),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_167),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_89),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_72),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_17),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_139),
.Y(n_197)
);

BUFx2_ASAP7_75t_SL g198 ( 
.A(n_92),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_74),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_46),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_137),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_14),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_55),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_46),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_3),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_62),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_77),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_144),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_8),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_126),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_31),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_27),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_80),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_70),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_33),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_27),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_147),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_98),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_94),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_115),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_60),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_26),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_82),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_65),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_71),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_60),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_138),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_96),
.Y(n_246)
);

BUFx2_ASAP7_75t_SL g247 ( 
.A(n_162),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_22),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_34),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_15),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_146),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_160),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_78),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_148),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_108),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_54),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_140),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_42),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_33),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_56),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_18),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_13),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_124),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_88),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_57),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_76),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_15),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_16),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_83),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_19),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_154),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_47),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_129),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_119),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_62),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_32),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_32),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_127),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_112),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_153),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_136),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_73),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_30),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_4),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_110),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_85),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_9),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_133),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_21),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_172),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_161),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_47),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_102),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_158),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_58),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_132),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_63),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_10),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_100),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_16),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_12),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_67),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_159),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_81),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_25),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_125),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_87),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_131),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_111),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_134),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_177),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_122),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_23),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_150),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_14),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_25),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_1),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_103),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_149),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_49),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_55),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_130),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_40),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_176),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_43),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_9),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_8),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_54),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_51),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_101),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_50),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_151),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_6),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_52),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_36),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_34),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_43),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_93),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_51),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_66),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_0),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_128),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_121),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_168),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_99),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_175),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_48),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_155),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_170),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_36),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_23),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_181),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_163),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_7),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_12),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_56),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_219),
.B(n_1),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_185),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_224),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_275),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_226),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_219),
.B(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_195),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_195),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_227),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_231),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_260),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_292),
.B(n_2),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_275),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_232),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_233),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_307),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_241),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_243),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_254),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_364),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_275),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_240),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_195),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_245),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_192),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_184),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_195),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_195),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_200),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_214),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_200),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_200),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_249),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_200),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_200),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_252),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_283),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_255),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_332),
.B(n_3),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_362),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_362),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_256),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_257),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_292),
.B(n_4),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_186),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_235),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_246),
.B(n_5),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_258),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_235),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_262),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_273),
.B(n_5),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_203),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_264),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_270),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_203),
.Y(n_436)
);

BUFx6f_ASAP7_75t_SL g437 ( 
.A(n_193),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_188),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_193),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_274),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_246),
.B(n_6),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_288),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_274),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_290),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_286),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_206),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_296),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_309),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_286),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_193),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_216),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_217),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_220),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_229),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_312),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_184),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_316),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_319),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_199),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_187),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_187),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_323),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_324),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_244),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_269),
.B(n_7),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_325),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_373),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_374),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_376),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_410),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_380),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_283),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_381),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_385),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_283),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_386),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_283),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_399),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_388),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_389),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_403),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_403),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_394),
.B(n_269),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_401),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_387),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_398),
.B(n_189),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_372),
.B(n_354),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_377),
.B(n_283),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

AND2x2_ASAP7_75t_SL g508 ( 
.A(n_423),
.B(n_360),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_439),
.B(n_223),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_408),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_408),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_395),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_414),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_391),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_439),
.B(n_223),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_375),
.B(n_360),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_404),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_384),
.B(n_273),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_414),
.B(n_205),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_418),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_409),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_420),
.A2(n_268),
.B(n_259),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_415),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_431),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_411),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g532 ( 
.A(n_434),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_421),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_435),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_416),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_444),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_448),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_424),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_455),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_442),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_438),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_508),
.B(n_392),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_501),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_536),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_504),
.B(n_503),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_478),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_303),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_522),
.B(n_457),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_508),
.A2(n_465),
.B1(n_383),
.B2(n_417),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

BUFx4f_ASAP7_75t_L g555 ( 
.A(n_532),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_508),
.B(n_303),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g557 ( 
.A(n_504),
.B(n_422),
.C(n_450),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_498),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_503),
.B(n_397),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_478),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_506),
.A2(n_328),
.B1(n_284),
.B2(n_298),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_518),
.B(n_520),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_496),
.B(n_303),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_518),
.B(n_520),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_328),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_412),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_520),
.B(n_461),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_496),
.B(n_458),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_462),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_470),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_496),
.B(n_303),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_467),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_500),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_198),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_523),
.B(n_450),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_490),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_496),
.B(n_463),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_538),
.B(n_390),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_496),
.B(n_459),
.Y(n_582)
);

OAI22x1_ASAP7_75t_L g583 ( 
.A1(n_509),
.A2(n_370),
.B1(n_194),
.B2(n_348),
.Y(n_583)
);

BUFx4f_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_478),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_521),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_476),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_521),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_521),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_469),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_487),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_506),
.B(n_436),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_487),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_490),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_506),
.B(n_303),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_506),
.B(n_222),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_469),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_506),
.A2(n_335),
.B1(n_369),
.B2(n_365),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_516),
.B(n_530),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_521),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_487),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_472),
.Y(n_603)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_527),
.B(n_367),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_523),
.B(n_433),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_521),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_494),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_230),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_501),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_506),
.B(n_347),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_493),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_493),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_468),
.B(n_438),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_483),
.B(n_367),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_536),
.B(n_440),
.Y(n_615)
);

INVx4_ASAP7_75t_SL g616 ( 
.A(n_476),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_493),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_533),
.B(n_447),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_506),
.B(n_483),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_468),
.B(n_367),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_499),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_471),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_533),
.B(n_466),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_483),
.B(n_367),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_471),
.Y(n_625)
);

BUFx4f_ASAP7_75t_L g626 ( 
.A(n_527),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_480),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_492),
.B(n_419),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_506),
.B(n_368),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_527),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_483),
.B(n_337),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_517),
.B(n_437),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_527),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_488),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_489),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_475),
.B(n_367),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_499),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_469),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_477),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_492),
.B(n_440),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_509),
.B(n_437),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_479),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_469),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_507),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_507),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_R g649 ( 
.A(n_482),
.B(n_354),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_486),
.B(n_443),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_473),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_473),
.B(n_247),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_491),
.B(n_513),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_473),
.B(n_218),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_473),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_519),
.B(n_437),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_526),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_511),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_534),
.A2(n_352),
.B1(n_346),
.B2(n_343),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_514),
.B(n_234),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_495),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_528),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_494),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_514),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_524),
.B(n_238),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_494),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_529),
.B(n_194),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_443),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_540),
.B(n_445),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_524),
.B(n_525),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_494),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_541),
.B(n_445),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_543),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_525),
.B(n_242),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_531),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_531),
.B(n_446),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_534),
.A2(n_350),
.B1(n_310),
.B2(n_277),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_534),
.B(n_446),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_485),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_545),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_545),
.B(n_253),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_545),
.B(n_449),
.C(n_228),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_485),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_495),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_485),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_494),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_494),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_545),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_545),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_485),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_545),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_515),
.B(n_474),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_505),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_545),
.B(n_272),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_549),
.B(n_546),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_554),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_559),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_586),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_560),
.B(n_301),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_563),
.B(n_515),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_563),
.B(n_515),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_559),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_588),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_563),
.B(n_566),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_SL g706 ( 
.A(n_568),
.B(n_276),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_556),
.A2(n_329),
.B1(n_355),
.B2(n_322),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_564),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_657),
.B(n_449),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_560),
.B(n_305),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_601),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_564),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_570),
.B(n_189),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_570),
.B(n_237),
.C(n_225),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_572),
.B(n_190),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_563),
.A2(n_197),
.B1(n_196),
.B2(n_191),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_584),
.B(n_282),
.Y(n_718)
);

AOI221xp5_ASAP7_75t_L g719 ( 
.A1(n_583),
.A2(n_278),
.B1(n_351),
.B2(n_221),
.C(n_212),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_572),
.B(n_190),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_563),
.B(n_474),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_584),
.B(n_287),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_605),
.B(n_451),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_566),
.B(n_474),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_626),
.B(n_289),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_615),
.B(n_451),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_591),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_558),
.B(n_452),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_606),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_SL g730 ( 
.A(n_555),
.B(n_642),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_566),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_591),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_593),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_566),
.A2(n_202),
.B1(n_208),
.B2(n_209),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_566),
.A2(n_202),
.B1(n_208),
.B2(n_209),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_626),
.B(n_297),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_582),
.B(n_505),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_628),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_593),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_548),
.B(n_539),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_585),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_553),
.A2(n_358),
.B1(n_210),
.B2(n_213),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_619),
.A2(n_502),
.B(n_497),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_552),
.B(n_542),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_550),
.B(n_505),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_550),
.B(n_505),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_561),
.B(n_505),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_561),
.B(n_505),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_668),
.B(n_210),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_668),
.B(n_213),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_669),
.B(n_215),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_618),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_694),
.B(n_300),
.Y(n_753)
);

O2A1O1Ixp5_ASAP7_75t_L g754 ( 
.A1(n_556),
.A2(n_334),
.B(n_333),
.C(n_326),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_631),
.A2(n_634),
.B(n_604),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_553),
.A2(n_327),
.B1(n_306),
.B2(n_315),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_571),
.B(n_302),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_672),
.B(n_215),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_631),
.A2(n_320),
.B1(n_304),
.B2(n_317),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_643),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_580),
.B(n_537),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_650),
.B(n_279),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_622),
.B(n_537),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_602),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_551),
.B(n_279),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_625),
.B(n_497),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_627),
.B(n_497),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_638),
.B(n_281),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_629),
.B(n_502),
.Y(n_769)
);

BUFx12f_ASAP7_75t_SL g770 ( 
.A(n_569),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_638),
.B(n_281),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_644),
.A2(n_358),
.B1(n_339),
.B2(n_345),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_602),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_579),
.B(n_544),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_594),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_694),
.B(n_339),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_604),
.B(n_345),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_510),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_621),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_637),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_644),
.A2(n_359),
.B1(n_361),
.B2(n_363),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_592),
.A2(n_512),
.B(n_510),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_647),
.B(n_512),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_611),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_599),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_648),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_680),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_633),
.A2(n_464),
.B(n_454),
.C(n_453),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_581),
.B(n_353),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_581),
.B(n_235),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_634),
.B(n_353),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_611),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_598),
.A2(n_359),
.B1(n_357),
.B2(n_361),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_596),
.B(n_357),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_658),
.B(n_481),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_664),
.Y(n_796)
);

AOI22x1_ASAP7_75t_L g797 ( 
.A1(n_651),
.A2(n_363),
.B1(n_464),
.B2(n_454),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_SL g798 ( 
.A1(n_576),
.A2(n_204),
.B1(n_236),
.B2(n_285),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_612),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_547),
.B(n_341),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_633),
.B(n_239),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_675),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_562),
.A2(n_223),
.B1(n_481),
.B2(n_476),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_578),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_562),
.A2(n_481),
.B1(n_476),
.B2(n_201),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_613),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_612),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_598),
.A2(n_610),
.B1(n_608),
.B2(n_630),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_576),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_614),
.A2(n_481),
.B(n_476),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_656),
.B(n_248),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_632),
.A2(n_313),
.B1(n_294),
.B2(n_280),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_656),
.B(n_250),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_551),
.B(n_481),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_613),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_609),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_670),
.B(n_251),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_682),
.B(n_613),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_551),
.B(n_476),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_577),
.B(n_261),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_676),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_551),
.B(n_481),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_624),
.A2(n_293),
.B1(n_295),
.B2(n_263),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_568),
.B(n_265),
.Y(n_824)
);

OAI22x1_ASAP7_75t_SL g825 ( 
.A1(n_575),
.A2(n_370),
.B1(n_221),
.B2(n_212),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_676),
.Y(n_826)
);

OAI221xp5_ASAP7_75t_L g827 ( 
.A1(n_659),
.A2(n_677),
.B1(n_674),
.B2(n_665),
.C(n_660),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_551),
.B(n_476),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_557),
.B(n_481),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_617),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_618),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_679),
.B(n_481),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_577),
.B(n_266),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_577),
.B(n_683),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_685),
.B(n_481),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_624),
.A2(n_201),
.B1(n_207),
.B2(n_211),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_617),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_676),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_640),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_690),
.B(n_267),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_640),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_661),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_639),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_568),
.B(n_271),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_667),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_568),
.B(n_291),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_565),
.A2(n_430),
.B(n_429),
.C(n_428),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_661),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_590),
.B(n_597),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_684),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_590),
.B(n_597),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_565),
.A2(n_207),
.B1(n_211),
.B2(n_278),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_678),
.B(n_426),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_573),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_641),
.B(n_299),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_574),
.A2(n_430),
.B(n_429),
.C(n_428),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_641),
.B(n_308),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_649),
.B(n_336),
.C(n_311),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_587),
.B(n_636),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_678),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_649),
.A2(n_314),
.B1(n_318),
.B2(n_321),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_755),
.A2(n_808),
.B(n_696),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_696),
.B(n_653),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_737),
.A2(n_595),
.B(n_680),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_700),
.B(n_653),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_700),
.A2(n_623),
.B1(n_673),
.B2(n_642),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_779),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_718),
.A2(n_574),
.B(n_692),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_730),
.B(n_662),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_718),
.A2(n_725),
.B(n_722),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_711),
.B(n_646),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_756),
.A2(n_623),
.B1(n_673),
.B2(n_662),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_761),
.A2(n_595),
.B(n_691),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_646),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_777),
.A2(n_681),
.B(n_654),
.C(n_652),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_722),
.A2(n_736),
.B(n_725),
.Y(n_876)
);

AND2x6_ASAP7_75t_SL g877 ( 
.A(n_774),
.B(n_567),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_860),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_736),
.A2(n_691),
.B(n_689),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_705),
.A2(n_689),
.B(n_663),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_701),
.B(n_555),
.Y(n_881)
);

NOR2x1_ASAP7_75t_L g882 ( 
.A(n_715),
.B(n_569),
.Y(n_882)
);

AOI21x1_ASAP7_75t_L g883 ( 
.A1(n_721),
.A2(n_724),
.B(n_832),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_780),
.B(n_569),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_745),
.A2(n_671),
.B(n_663),
.Y(n_885)
);

OR2x2_ASAP7_75t_SL g886 ( 
.A(n_858),
.B(n_600),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_746),
.A2(n_671),
.B(n_666),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_806),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_716),
.B(n_714),
.Y(n_889)
);

NOR2x1_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_567),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_716),
.A2(n_655),
.B(n_659),
.C(n_677),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_747),
.A2(n_666),
.B(n_587),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_787),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_714),
.A2(n_678),
.B(n_681),
.C(n_687),
.Y(n_894)
);

BUFx8_ASAP7_75t_L g895 ( 
.A(n_809),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_752),
.B(n_603),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_791),
.A2(n_684),
.B(n_687),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_791),
.A2(n_636),
.B(n_587),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_816),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_768),
.A2(n_771),
.B(n_801),
.C(n_817),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_748),
.A2(n_587),
.B(n_636),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_817),
.B(n_599),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_702),
.A2(n_636),
.B(n_686),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_699),
.B(n_693),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_SL g905 ( 
.A(n_801),
.B(n_575),
.C(n_351),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_704),
.B(n_693),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_849),
.A2(n_693),
.B(n_686),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_851),
.A2(n_693),
.B(n_686),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_777),
.A2(n_567),
.B1(n_330),
.B2(n_331),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_738),
.B(n_603),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_785),
.A2(n_686),
.B(n_599),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_710),
.B(n_599),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_843),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_815),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_759),
.A2(n_607),
.B1(n_340),
.B2(n_348),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_743),
.A2(n_753),
.B(n_782),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_787),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_785),
.A2(n_607),
.B(n_688),
.Y(n_918)
);

INVxp33_ASAP7_75t_SL g919 ( 
.A(n_798),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_786),
.B(n_616),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_728),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_831),
.B(n_603),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_859),
.A2(n_607),
.B(n_688),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_859),
.A2(n_607),
.B(n_688),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_855),
.A2(n_616),
.B(n_427),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_857),
.A2(n_757),
.B(n_795),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_812),
.B(n_280),
.C(n_340),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_763),
.A2(n_620),
.B(n_349),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_728),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_776),
.A2(n_349),
.B(n_356),
.C(n_341),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_712),
.B(n_645),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_821),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_729),
.B(n_645),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_835),
.A2(n_620),
.B(n_356),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_796),
.B(n_802),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_760),
.B(n_573),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_826),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_789),
.B(n_620),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_789),
.B(n_620),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_768),
.B(n_620),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_804),
.B(n_13),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_762),
.B(n_20),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_707),
.A2(n_75),
.B1(n_182),
.B2(n_180),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_753),
.A2(n_342),
.B1(n_341),
.B2(n_26),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_838),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_818),
.A2(n_68),
.B(n_178),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_818),
.A2(n_64),
.B(n_174),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_762),
.A2(n_342),
.B(n_22),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_720),
.B(n_20),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_853),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_818),
.A2(n_767),
.B(n_766),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_769),
.A2(n_84),
.B(n_156),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_719),
.B(n_750),
.C(n_749),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_771),
.B(n_29),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_723),
.B(n_30),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_741),
.B(n_31),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_775),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_717),
.A2(n_90),
.B1(n_145),
.B2(n_141),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_811),
.B(n_342),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_776),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_778),
.A2(n_123),
.B(n_118),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_853),
.B(n_113),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_787),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_852),
.A2(n_742),
.B(n_836),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_SL g965 ( 
.A(n_787),
.B(n_38),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_800),
.B(n_39),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_728),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_811),
.A2(n_39),
.B(n_41),
.C(n_42),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_827),
.A2(n_44),
.B(n_45),
.C(n_48),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_853),
.B(n_44),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_783),
.A2(n_95),
.B(n_114),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_726),
.B(n_52),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_794),
.A2(n_105),
.B(n_107),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_794),
.A2(n_53),
.B(n_59),
.C(n_61),
.Y(n_974)
);

NOR2xp67_ASAP7_75t_L g975 ( 
.A(n_854),
.B(n_106),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_847),
.A2(n_53),
.B(n_61),
.C(n_63),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_790),
.B(n_751),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_731),
.A2(n_734),
.B1(n_735),
.B2(n_834),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_840),
.B(n_695),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_754),
.A2(n_697),
.B(n_698),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_709),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_703),
.A2(n_807),
.B(n_708),
.Y(n_982)
);

OAI321xp33_ASAP7_75t_L g983 ( 
.A1(n_772),
.A2(n_781),
.A3(n_861),
.B1(n_823),
.B2(n_820),
.C(n_833),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_740),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_708),
.A2(n_830),
.B(n_850),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_856),
.A2(n_788),
.B(n_829),
.C(n_793),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_758),
.A2(n_709),
.B1(n_845),
.B2(n_797),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_713),
.A2(n_850),
.B(n_727),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_713),
.A2(n_848),
.B(n_727),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_732),
.A2(n_848),
.B(n_733),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_732),
.A2(n_841),
.B(n_733),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_744),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_739),
.A2(n_799),
.B(n_764),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_764),
.B(n_830),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_820),
.B(n_833),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_813),
.B(n_837),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_773),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_784),
.A2(n_841),
.B(n_842),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_770),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_784),
.B(n_837),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_792),
.B(n_839),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_799),
.B(n_842),
.Y(n_1002)
);

AO21x1_ASAP7_75t_L g1003 ( 
.A1(n_824),
.A2(n_846),
.B(n_844),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_839),
.A2(n_765),
.B(n_828),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_805),
.B(n_810),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_814),
.B(n_819),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_822),
.B(n_803),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_706),
.B(n_825),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_695),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_700),
.A2(n_549),
.B(n_711),
.C(n_716),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_700),
.B(n_711),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_696),
.B(n_549),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_700),
.B(n_711),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_696),
.B(n_549),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_860),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_700),
.A2(n_549),
.B(n_711),
.C(n_716),
.Y(n_1018)
);

NOR2x1p5_ASAP7_75t_L g1019 ( 
.A(n_858),
.B(n_642),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_816),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_696),
.B(n_549),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_860),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_787),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_779),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_L g1029 ( 
.A(n_816),
.B(n_843),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_860),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_816),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_696),
.B(n_549),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_696),
.B(n_549),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_700),
.B(n_711),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_700),
.A2(n_549),
.B1(n_566),
.B2(n_563),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_696),
.B(n_549),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_700),
.A2(n_549),
.B(n_711),
.C(n_716),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_737),
.A2(n_761),
.B(n_619),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_696),
.B(n_549),
.Y(n_1041)
);

BUFx4f_ASAP7_75t_SL g1042 ( 
.A(n_1028),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_1012),
.A2(n_1036),
.B(n_1014),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1012),
.A2(n_1014),
.B(n_1036),
.C(n_1018),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_900),
.A2(n_1011),
.A3(n_1039),
.B(n_1003),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_889),
.A2(n_1015),
.B(n_1013),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_865),
.B(n_984),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_942),
.A2(n_866),
.B(n_944),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1021),
.B(n_1032),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_902),
.A2(n_876),
.B(n_870),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1009),
.A2(n_1022),
.B(n_1017),
.Y(n_1051)
);

OA22x2_ASAP7_75t_L g1052 ( 
.A1(n_964),
.A2(n_948),
.B1(n_872),
.B2(n_992),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1023),
.A2(n_1027),
.B(n_1024),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_883),
.A2(n_1004),
.B(n_880),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1033),
.A2(n_1041),
.B(n_1038),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_995),
.B(n_992),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_863),
.B(n_871),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_862),
.A2(n_1037),
.B(n_1005),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1007),
.A2(n_1040),
.B(n_1034),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_951),
.A2(n_1006),
.B(n_926),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_867),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_874),
.B(n_942),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_977),
.B(n_983),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_899),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_894),
.A2(n_954),
.A3(n_968),
.B(n_891),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_977),
.A2(n_978),
.B(n_949),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_878),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_873),
.A2(n_868),
.B(n_864),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_997),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_935),
.B(n_953),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_986),
.A2(n_916),
.B(n_979),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_950),
.B(n_962),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_913),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_953),
.B(n_869),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_938),
.A2(n_939),
.B(n_940),
.C(n_973),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_875),
.A2(n_897),
.B(n_991),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_944),
.A2(n_949),
.B1(n_927),
.B2(n_958),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_895),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_963),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1020),
.B(n_955),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_927),
.B(n_941),
.C(n_896),
.Y(n_1081)
);

AO21x1_ASAP7_75t_L g1082 ( 
.A1(n_969),
.A2(n_960),
.B(n_974),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_972),
.B(n_888),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_922),
.B1(n_981),
.B2(n_1035),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_922),
.A2(n_981),
.B1(n_1016),
.B2(n_1025),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_885),
.A2(n_887),
.B(n_879),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_972),
.B(n_914),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1030),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_SL g1089 ( 
.A1(n_946),
.A2(n_947),
.B(n_976),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_932),
.B(n_937),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_918),
.A2(n_903),
.B(n_923),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1031),
.Y(n_1092)
);

AO21x2_ASAP7_75t_L g1093 ( 
.A1(n_980),
.A2(n_907),
.B(n_908),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_SL g1094 ( 
.A1(n_970),
.A2(n_971),
.B(n_961),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_924),
.A2(n_898),
.B(n_892),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_881),
.A2(n_912),
.B(n_906),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_930),
.A2(n_959),
.B(n_1020),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_982),
.A2(n_998),
.B(n_985),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_963),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_945),
.B(n_996),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_905),
.B(n_933),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_966),
.B(n_962),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_987),
.A2(n_1019),
.B1(n_882),
.B2(n_884),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1002),
.B(n_956),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_881),
.A2(n_904),
.B(n_1001),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_989),
.A2(n_990),
.B(n_993),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_988),
.A2(n_911),
.B(n_994),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1010),
.B(n_931),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_941),
.A2(n_936),
.B(n_965),
.C(n_975),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1000),
.A2(n_925),
.B(n_901),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_893),
.B(n_1026),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_997),
.B(n_917),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_963),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_963),
.Y(n_1114)
);

OAI211xp5_ASAP7_75t_L g1115 ( 
.A1(n_921),
.A2(n_929),
.B(n_967),
.C(n_890),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_934),
.A2(n_928),
.B(n_920),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_917),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_936),
.B(n_893),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_909),
.A2(n_884),
.B(n_952),
.C(n_943),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_920),
.A2(n_915),
.B(n_1029),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_910),
.A2(n_1008),
.B(n_929),
.C(n_921),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_919),
.A2(n_957),
.B(n_981),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_981),
.B(n_1026),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1026),
.A2(n_999),
.B(n_886),
.Y(n_1124)
);

OAI22x1_ASAP7_75t_L g1125 ( 
.A1(n_877),
.A2(n_1012),
.B1(n_1036),
.B2(n_1014),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_895),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1026),
.A2(n_1040),
.B(n_1034),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_SL g1128 ( 
.A1(n_973),
.A2(n_1003),
.B(n_947),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1012),
.A2(n_1036),
.B(n_1014),
.C(n_1018),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1011),
.A2(n_1039),
.B(n_1018),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_883),
.A2(n_1004),
.B(n_880),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_997),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_883),
.A2(n_1004),
.B(n_880),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1139)
);

AO21x2_ASAP7_75t_L g1140 ( 
.A1(n_862),
.A2(n_900),
.B(n_916),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1031),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1011),
.A2(n_1039),
.B(n_1018),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_997),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1012),
.A2(n_1036),
.B(n_1014),
.C(n_1018),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_900),
.A2(n_1018),
.A3(n_1039),
.B(n_1011),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_867),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1012),
.A2(n_1036),
.B1(n_1014),
.B2(n_889),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_997),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_916),
.A2(n_883),
.B(n_876),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_889),
.A2(n_1011),
.B1(n_1039),
.B2(n_1018),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1028),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_883),
.A2(n_1004),
.B(n_880),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1012),
.A2(n_1014),
.B1(n_1036),
.B2(n_889),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_867),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1011),
.A2(n_1039),
.B(n_1018),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1011),
.A2(n_1039),
.B(n_1018),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_916),
.A2(n_883),
.B(n_876),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1011),
.A2(n_1039),
.B(n_1018),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_L g1170 ( 
.A1(n_902),
.A2(n_876),
.B(n_870),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_878),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_889),
.A2(n_1011),
.B1(n_1039),
.B2(n_1018),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_883),
.A2(n_1004),
.B(n_880),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_916),
.A2(n_883),
.B(n_876),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_916),
.A2(n_883),
.B(n_876),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1012),
.A2(n_1036),
.B(n_1014),
.C(n_1018),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_902),
.A2(n_876),
.B(n_870),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_900),
.B(n_889),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1011),
.A2(n_1039),
.B1(n_1018),
.B2(n_1012),
.C(n_1036),
.Y(n_1183)
);

AND3x2_ASAP7_75t_L g1184 ( 
.A(n_1012),
.B(n_1036),
.C(n_1014),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_900),
.B(n_889),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_SL g1186 ( 
.A1(n_973),
.A2(n_1003),
.B(n_947),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_889),
.A2(n_1011),
.B1(n_1039),
.B2(n_1018),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1012),
.A2(n_1036),
.B(n_1014),
.C(n_1018),
.Y(n_1188)
);

NAND2x1_ASAP7_75t_L g1189 ( 
.A(n_893),
.B(n_963),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1031),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1012),
.B(n_1036),
.C(n_1014),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1031),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1009),
.A2(n_1040),
.B(n_1034),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_999),
.B(n_816),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_867),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1042),
.Y(n_1198)
);

INVx3_ASAP7_75t_SL g1199 ( 
.A(n_1197),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1190),
.A2(n_1043),
.B(n_1148),
.C(n_1048),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1201)
);

BUFx12f_ASAP7_75t_L g1202 ( 
.A(n_1126),
.Y(n_1202)
);

BUFx10_ASAP7_75t_L g1203 ( 
.A(n_1197),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1192),
.B(n_1130),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1141),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1124),
.B(n_1196),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1141),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1208)
);

AND2x6_ASAP7_75t_L g1209 ( 
.A(n_1072),
.B(n_1063),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1088),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1051),
.A2(n_1134),
.B(n_1053),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1063),
.A2(n_1160),
.B1(n_1178),
.B2(n_1133),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1137),
.A2(n_1149),
.B(n_1139),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1181),
.B(n_1136),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1042),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1073),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1114),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1114),
.B(n_1189),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1047),
.B(n_1056),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1147),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1150),
.A2(n_1158),
.B(n_1152),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1191),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1160),
.B(n_1066),
.C(n_1129),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1072),
.B(n_1191),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1163),
.A2(n_1195),
.B(n_1194),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1135),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1092),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1172),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1168),
.B(n_1169),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1174),
.B(n_1046),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1114),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1161),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1131),
.A2(n_1166),
.B(n_1142),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1072),
.B(n_1193),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1157),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1044),
.B(n_1129),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1049),
.B(n_1044),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1103),
.B(n_1102),
.Y(n_1239)
);

INVx3_ASAP7_75t_SL g1240 ( 
.A(n_1078),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1114),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1079),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1060),
.A2(n_1059),
.B(n_1127),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1064),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1144),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_SL g1246 ( 
.A1(n_1145),
.A2(n_1188),
.B(n_1179),
.C(n_1182),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1078),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1071),
.A2(n_1182),
.B(n_1185),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1061),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1090),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1145),
.A2(n_1188),
.B(n_1179),
.C(n_1162),
.Y(n_1251)
);

BUFx4_ASAP7_75t_SL g1252 ( 
.A(n_1196),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1111),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1196),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1100),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1080),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1123),
.B(n_1120),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1125),
.B(n_1101),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1079),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1111),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1057),
.B(n_1062),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1101),
.B(n_1052),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1113),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1074),
.B(n_1113),
.Y(n_1264)
);

CKINVDCx6p67_ASAP7_75t_R g1265 ( 
.A(n_1074),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1122),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1153),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1099),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1077),
.A2(n_1173),
.B1(n_1187),
.B2(n_1156),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1185),
.A2(n_1076),
.B(n_1086),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1184),
.Y(n_1271)
);

NOR2x1_ASAP7_75t_SL g1272 ( 
.A(n_1118),
.B(n_1085),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1077),
.A2(n_1164),
.B1(n_1052),
.B2(n_1081),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1070),
.A2(n_1083),
.B1(n_1087),
.B2(n_1104),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1108),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1058),
.A2(n_1068),
.B(n_1140),
.Y(n_1276)
);

NOR2xp67_ASAP7_75t_L g1277 ( 
.A(n_1115),
.B(n_1117),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1140),
.A2(n_1095),
.B(n_1098),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1112),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1055),
.B(n_1183),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1099),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1082),
.A2(n_1184),
.B1(n_1097),
.B2(n_1089),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1146),
.B(n_1045),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1146),
.B(n_1045),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1146),
.B(n_1045),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1084),
.A2(n_1109),
.B1(n_1121),
.B2(n_1116),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1045),
.B(n_1109),
.Y(n_1287)
);

CKINVDCx16_ASAP7_75t_R g1288 ( 
.A(n_1121),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1096),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1065),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1065),
.B(n_1119),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1119),
.A2(n_1105),
.B1(n_1180),
.B2(n_1170),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1155),
.B(n_1165),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1155),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1176),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1075),
.A2(n_1106),
.B(n_1177),
.C(n_1176),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1094),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1128),
.B(n_1186),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1110),
.A2(n_1075),
.B(n_1091),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1093),
.A2(n_1132),
.B(n_1054),
.Y(n_1300)
);

CKINVDCx6p67_ASAP7_75t_R g1301 ( 
.A(n_1050),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1093),
.B(n_1107),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1138),
.Y(n_1303)
);

OR2x6_ASAP7_75t_SL g1304 ( 
.A(n_1159),
.B(n_1175),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1051),
.A2(n_1134),
.B(n_1053),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1044),
.A2(n_1018),
.B(n_1039),
.C(n_1011),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1067),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1047),
.B(n_1151),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1114),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1072),
.B(n_1141),
.Y(n_1311)
);

INVx3_ASAP7_75t_SL g1312 ( 
.A(n_1197),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1197),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1042),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1114),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1067),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1141),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1190),
.A2(n_919),
.B1(n_1014),
.B2(n_1012),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1042),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1072),
.B(n_1141),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1073),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1069),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1073),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1063),
.A2(n_1012),
.B(n_1036),
.C(n_1014),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1051),
.A2(n_1134),
.B(n_1053),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1192),
.B(n_779),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1051),
.A2(n_1134),
.B(n_1053),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1047),
.B(n_1151),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1047),
.B(n_1151),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1066),
.B(n_889),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1047),
.B(n_1151),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1190),
.A2(n_1012),
.B1(n_1036),
.B2(n_1014),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1114),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1066),
.B(n_889),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1114),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1073),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1190),
.B(n_1151),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1190),
.A2(n_1012),
.B1(n_1036),
.B2(n_1014),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1114),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1190),
.A2(n_1012),
.B1(n_1036),
.B2(n_1014),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1042),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1319),
.A2(n_1269),
.B1(n_1335),
.B2(n_1343),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1300),
.A2(n_1213),
.B(n_1211),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1247),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1284),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1262),
.B(n_1212),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1299),
.A2(n_1243),
.B(n_1278),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1335),
.A2(n_1343),
.B1(n_1341),
.B2(n_1239),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1299),
.A2(n_1243),
.B(n_1278),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1283),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1227),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1318),
.Y(n_1355)
);

BUFx2_ASAP7_75t_SL g1356 ( 
.A(n_1342),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1285),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1265),
.A2(n_1266),
.B1(n_1220),
.B2(n_1204),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1341),
.A2(n_1239),
.B1(n_1224),
.B2(n_1273),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1342),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1230),
.B(n_1309),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1212),
.B(n_1200),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1290),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1264),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1211),
.A2(n_1226),
.B(n_1222),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1247),
.Y(n_1366)
);

CKINVDCx14_ASAP7_75t_R g1367 ( 
.A(n_1313),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1267),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1264),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1323),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1342),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1209),
.Y(n_1372)
);

INVx11_ASAP7_75t_L g1373 ( 
.A(n_1233),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1322),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1258),
.A2(n_1237),
.B1(n_1209),
.B2(n_1286),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1215),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1276),
.A2(n_1292),
.B(n_1270),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1236),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1318),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1214),
.A2(n_1305),
.B1(n_1314),
.B2(n_1340),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1287),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1324),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1271),
.A2(n_1206),
.B1(n_1273),
.B2(n_1201),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1237),
.A2(n_1333),
.B1(n_1337),
.B2(n_1234),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1294),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1291),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1339),
.Y(n_1388)
);

AO21x1_ASAP7_75t_L g1389 ( 
.A1(n_1307),
.A2(n_1333),
.B(n_1337),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1339),
.Y(n_1390)
);

CKINVDCx6p67_ASAP7_75t_R g1391 ( 
.A(n_1199),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1276),
.A2(n_1270),
.B(n_1327),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1234),
.A2(n_1274),
.B1(n_1328),
.B2(n_1209),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1325),
.A2(n_1330),
.B1(n_1261),
.B2(n_1208),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1210),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1203),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1209),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1222),
.A2(n_1329),
.B(n_1306),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1229),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1226),
.A2(n_1306),
.B(n_1329),
.Y(n_1400)
);

CKINVDCx6p67_ASAP7_75t_R g1401 ( 
.A(n_1199),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1217),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1205),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1312),
.Y(n_1404)
);

CKINVDCx6p67_ASAP7_75t_R g1405 ( 
.A(n_1312),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1244),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1308),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1317),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1331),
.B(n_1332),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1295),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1295),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1209),
.A2(n_1282),
.B1(n_1231),
.B2(n_1206),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1216),
.Y(n_1413)
);

BUFx4_ASAP7_75t_R g1414 ( 
.A(n_1203),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1327),
.A2(n_1302),
.B(n_1248),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1320),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1200),
.A2(n_1250),
.B1(n_1282),
.B2(n_1275),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1334),
.B(n_1219),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1206),
.A2(n_1249),
.B1(n_1221),
.B2(n_1257),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1288),
.A2(n_1255),
.B1(n_1272),
.B2(n_1298),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1257),
.B(n_1297),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_SL g1422 ( 
.A1(n_1307),
.A2(n_1248),
.B(n_1238),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1256),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1242),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1257),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1280),
.A2(n_1254),
.B1(n_1235),
.B2(n_1277),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1281),
.Y(n_1427)
);

CKINVDCx6p67_ASAP7_75t_R g1428 ( 
.A(n_1240),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1326),
.B(n_1279),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1245),
.B(n_1251),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1289),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1293),
.A2(n_1218),
.B(n_1304),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1198),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1289),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1242),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1289),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1245),
.Y(n_1437)
);

INVx6_ASAP7_75t_L g1438 ( 
.A(n_1223),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1246),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1252),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1251),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1301),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1223),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1281),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1235),
.A2(n_1321),
.B1(n_1225),
.B2(n_1311),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1303),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1253),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1303),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1296),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1225),
.Y(n_1450)
);

OAI21xp33_ASAP7_75t_L g1451 ( 
.A1(n_1228),
.A2(n_1344),
.B(n_1315),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1242),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1252),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1296),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1232),
.B(n_1338),
.Y(n_1455)
);

AO21x1_ASAP7_75t_L g1456 ( 
.A1(n_1326),
.A2(n_1218),
.B(n_1241),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1259),
.Y(n_1457)
);

BUFx12f_ASAP7_75t_L g1458 ( 
.A(n_1320),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1259),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1232),
.B(n_1338),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1311),
.A2(n_1321),
.B1(n_1202),
.B2(n_1240),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1207),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1217),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1268),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1316),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1263),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1253),
.A2(n_1260),
.B1(n_1310),
.B2(n_1316),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1253),
.A2(n_1260),
.B1(n_1310),
.B2(n_1241),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1336),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1260),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1336),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1336),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1387),
.B(n_1336),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1387),
.B(n_1353),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1347),
.Y(n_1475)
);

NAND2x1_ASAP7_75t_L g1476 ( 
.A(n_1372),
.B(n_1397),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1421),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1386),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1406),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1382),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1410),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1353),
.B(n_1357),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1357),
.B(n_1349),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1400),
.A2(n_1398),
.B(n_1365),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1382),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1378),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1411),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1425),
.B(n_1421),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1425),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1421),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1349),
.B(n_1381),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1380),
.B(n_1394),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1348),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1363),
.Y(n_1494)
);

BUFx8_ASAP7_75t_L g1495 ( 
.A(n_1396),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1372),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1363),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1421),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1346),
.A2(n_1454),
.B(n_1449),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1372),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1409),
.B(n_1361),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1430),
.B(n_1385),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1423),
.B(n_1418),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1430),
.B(n_1362),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1398),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1415),
.A2(n_1377),
.B(n_1392),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1362),
.B(n_1364),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1395),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1364),
.B(n_1369),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1367),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1383),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1413),
.Y(n_1512)
);

BUFx4f_ASAP7_75t_L g1513 ( 
.A(n_1397),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1399),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1383),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1350),
.A2(n_1352),
.B(n_1415),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1432),
.A2(n_1422),
.B(n_1448),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1432),
.A2(n_1422),
.B(n_1448),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1390),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1389),
.B(n_1446),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1369),
.B(n_1437),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1429),
.B(n_1350),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1437),
.B(n_1359),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1417),
.B(n_1384),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1389),
.A2(n_1393),
.B(n_1412),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1374),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1407),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1427),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1441),
.B(n_1408),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1358),
.B(n_1388),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1347),
.Y(n_1532)
);

AO21x2_ASAP7_75t_L g1533 ( 
.A1(n_1350),
.A2(n_1352),
.B(n_1400),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1436),
.A2(n_1456),
.B(n_1439),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1356),
.B(n_1442),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1427),
.Y(n_1536)
);

BUFx2_ASAP7_75t_SL g1537 ( 
.A(n_1442),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1444),
.Y(n_1538)
);

AOI21xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1419),
.A2(n_1375),
.B(n_1440),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1352),
.A2(n_1431),
.B(n_1434),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1438),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1345),
.B(n_1351),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1355),
.Y(n_1544)
);

AOI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1466),
.A2(n_1457),
.B(n_1452),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1420),
.A2(n_1426),
.B(n_1451),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1413),
.B(n_1354),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1501),
.B(n_1462),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1524),
.A2(n_1428),
.B1(n_1461),
.B2(n_1450),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1483),
.B(n_1472),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1478),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1540),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1477),
.B(n_1470),
.Y(n_1553)
);

AO21x1_ASAP7_75t_L g1554 ( 
.A1(n_1492),
.A2(n_1472),
.B(n_1469),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1546),
.A2(n_1428),
.B1(n_1450),
.B2(n_1433),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1483),
.B(n_1502),
.Y(n_1556)
);

NAND2x1_ASAP7_75t_L g1557 ( 
.A(n_1535),
.B(n_1435),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1471),
.Y(n_1558)
);

NAND2x1_ASAP7_75t_L g1559 ( 
.A(n_1535),
.B(n_1435),
.Y(n_1559)
);

AO21x2_ASAP7_75t_L g1560 ( 
.A1(n_1484),
.A2(n_1471),
.B(n_1452),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1540),
.B(n_1463),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1543),
.A2(n_1433),
.B1(n_1453),
.B2(n_1464),
.C(n_1445),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1499),
.B(n_1463),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1499),
.B(n_1465),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1539),
.A2(n_1405),
.B1(n_1391),
.B2(n_1401),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1520),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1502),
.B(n_1460),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1522),
.B(n_1379),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1490),
.B(n_1498),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1522),
.B(n_1370),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1488),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1535),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1482),
.B(n_1368),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1525),
.A2(n_1366),
.B1(n_1404),
.B2(n_1440),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1520),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1489),
.B(n_1379),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1491),
.B(n_1460),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1491),
.B(n_1455),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1356),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1504),
.B(n_1455),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1488),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1504),
.B(n_1470),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1474),
.B(n_1447),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1503),
.B(n_1486),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1533),
.B(n_1402),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1531),
.A2(n_1405),
.B1(n_1391),
.B2(n_1401),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1507),
.B(n_1459),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1489),
.B(n_1355),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1556),
.B(n_1507),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1574),
.A2(n_1539),
.B1(n_1479),
.B2(n_1512),
.C(n_1537),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1555),
.A2(n_1520),
.B1(n_1535),
.B2(n_1488),
.C(n_1547),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1585),
.B(n_1488),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1574),
.A2(n_1513),
.B1(n_1488),
.B2(n_1537),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1554),
.A2(n_1513),
.B(n_1525),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1567),
.B(n_1527),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1585),
.B(n_1481),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1586),
.A2(n_1513),
.B1(n_1498),
.B2(n_1525),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1542),
.C(n_1476),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1480),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1577),
.B(n_1485),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1565),
.A2(n_1515),
.B1(n_1526),
.B2(n_1511),
.C(n_1519),
.Y(n_1601)
);

AOI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1554),
.A2(n_1523),
.B(n_1536),
.C(n_1538),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1586),
.A2(n_1523),
.B(n_1467),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1548),
.B(n_1414),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1549),
.A2(n_1513),
.B1(n_1525),
.B2(n_1468),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1521),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1521),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1529),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1584),
.B(n_1529),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1562),
.A2(n_1403),
.B1(n_1476),
.B2(n_1542),
.C(n_1544),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1551),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1550),
.B(n_1570),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1562),
.A2(n_1438),
.B1(n_1443),
.B2(n_1544),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1579),
.B(n_1496),
.Y(n_1614)
);

NAND4xp25_ASAP7_75t_L g1615 ( 
.A(n_1568),
.B(n_1541),
.C(n_1403),
.D(n_1528),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1550),
.B(n_1509),
.Y(n_1616)
);

OAI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1579),
.A2(n_1443),
.B1(n_1438),
.B2(n_1510),
.C(n_1500),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1552),
.A2(n_1506),
.B(n_1505),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1509),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1396),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1571),
.A2(n_1475),
.B1(n_1532),
.B2(n_1496),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1558),
.B(n_1487),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1573),
.B(n_1508),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1557),
.A2(n_1518),
.B(n_1517),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1573),
.B(n_1587),
.Y(n_1625)
);

AND2x2_ASAP7_75t_SL g1626 ( 
.A(n_1572),
.B(n_1493),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1552),
.B(n_1494),
.C(n_1497),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1587),
.B(n_1580),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1558),
.B(n_1487),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1558),
.B(n_1494),
.C(n_1497),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1561),
.B(n_1517),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1583),
.B(n_1514),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1557),
.A2(n_1518),
.B(n_1534),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1551),
.Y(n_1634)
);

OAI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1566),
.A2(n_1530),
.B(n_1473),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1559),
.A2(n_1533),
.B(n_1516),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1561),
.B(n_1576),
.C(n_1588),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1553),
.B(n_1496),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1611),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1611),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1634),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1626),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1626),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1634),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1618),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1622),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1592),
.B(n_1572),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1622),
.B(n_1561),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1637),
.B(n_1575),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1592),
.Y(n_1652)
);

INVx6_ASAP7_75t_L g1653 ( 
.A(n_1629),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1560),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1563),
.Y(n_1655)
);

CKINVDCx8_ASAP7_75t_R g1656 ( 
.A(n_1604),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1638),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1618),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1589),
.B(n_1563),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1632),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1630),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1619),
.B(n_1560),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1624),
.B(n_1572),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1625),
.B(n_1564),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_1609),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1627),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1623),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1618),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1614),
.B(n_1572),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1628),
.B(n_1564),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1599),
.B(n_1533),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_1594),
.B(n_1560),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1672),
.B(n_1608),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1639),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1672),
.B(n_1595),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1616),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1639),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1666),
.A2(n_1590),
.B(n_1673),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1672),
.B(n_1600),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1661),
.B(n_1606),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1640),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1652),
.B(n_1642),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1652),
.B(n_1571),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1652),
.B(n_1581),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1666),
.Y(n_1687)
);

OR3x2_ASAP7_75t_L g1688 ( 
.A(n_1651),
.B(n_1615),
.C(n_1495),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1656),
.B(n_1475),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1655),
.B(n_1607),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1660),
.B(n_1601),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1655),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1641),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1641),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1582),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1670),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1646),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1667),
.B(n_1671),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

AOI32xp33_ASAP7_75t_L g1702 ( 
.A1(n_1644),
.A2(n_1593),
.A3(n_1597),
.B1(n_1610),
.B2(n_1605),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1642),
.B(n_1581),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1642),
.B(n_1569),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1643),
.B(n_1569),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1646),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1646),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1643),
.B(n_1569),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1673),
.A2(n_1603),
.B(n_1591),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1648),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1648),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1643),
.B(n_1569),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1647),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1659),
.B(n_1633),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1692),
.B(n_1667),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1670),
.Y(n_1716)
);

NOR2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1690),
.B(n_1532),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1671),
.Y(n_1718)
);

AOI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1680),
.A2(n_1617),
.B(n_1663),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1720)
);

OAI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1709),
.A2(n_1651),
.B(n_1635),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1676),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1687),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1689),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1684),
.B(n_1704),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1693),
.B(n_1671),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1674),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1680),
.B(n_1656),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1676),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1674),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1682),
.B(n_1664),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1709),
.A2(n_1645),
.B(n_1644),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1674),
.Y(n_1734)
);

OAI21xp33_ASAP7_75t_L g1735 ( 
.A1(n_1702),
.A2(n_1651),
.B(n_1635),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1682),
.B(n_1664),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1679),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1679),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1683),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1683),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1684),
.B(n_1649),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1690),
.B(n_1664),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1681),
.B(n_1662),
.Y(n_1743)
);

AOI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1702),
.A2(n_1663),
.B(n_1621),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1698),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1691),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1691),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1704),
.B(n_1649),
.Y(n_1748)
);

AND2x2_ASAP7_75t_SL g1749 ( 
.A(n_1695),
.B(n_1645),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1695),
.B(n_1598),
.C(n_1613),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1700),
.B(n_1657),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_L g1752 ( 
.A(n_1701),
.B(n_1636),
.C(n_1656),
.Y(n_1752)
);

NOR2xp67_ASAP7_75t_L g1753 ( 
.A(n_1695),
.B(n_1657),
.Y(n_1753)
);

NAND2x1p5_ASAP7_75t_L g1754 ( 
.A(n_1695),
.B(n_1559),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1705),
.B(n_1663),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1705),
.B(n_1649),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1714),
.A2(n_1663),
.B(n_1669),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1722),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1749),
.B(n_1714),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1753),
.B(n_1663),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1729),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1737),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1738),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1749),
.B(n_1708),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1710),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1723),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1739),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1741),
.B(n_1708),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1728),
.B(n_1710),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1741),
.B(n_1712),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1724),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1754),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1728),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1727),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1740),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1748),
.B(n_1712),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1748),
.B(n_1703),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1742),
.B(n_1732),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1756),
.B(n_1703),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1745),
.Y(n_1781)
);

AO21x2_ASAP7_75t_L g1782 ( 
.A1(n_1733),
.A2(n_1752),
.B(n_1734),
.Y(n_1782)
);

NAND2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1717),
.B(n_1545),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1756),
.B(n_1685),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1731),
.Y(n_1785)
);

CKINVDCx16_ASAP7_75t_R g1786 ( 
.A(n_1725),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1719),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1746),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1731),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1754),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1721),
.B(n_1665),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1725),
.B(n_1685),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1735),
.B(n_1711),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1777),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1787),
.A2(n_1744),
.B1(n_1757),
.B2(n_1750),
.C(n_1716),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1772),
.B(n_1726),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1786),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1781),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1767),
.B(n_1747),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1786),
.A2(n_1688),
.B1(n_1755),
.B2(n_1669),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1787),
.A2(n_1688),
.B1(n_1751),
.B2(n_1755),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1767),
.B(n_1718),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1772),
.B(n_1736),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1781),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1774),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1777),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1791),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1774),
.A2(n_1754),
.B(n_1620),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1758),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1793),
.B(n_1694),
.Y(n_1810)
);

INVxp33_ASAP7_75t_L g1811 ( 
.A(n_1791),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1782),
.A2(n_1755),
.B1(n_1669),
.B2(n_1649),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1770),
.B(n_1657),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1793),
.A2(n_1743),
.B1(n_1730),
.B2(n_1720),
.C(n_1734),
.Y(n_1814)
);

AOI32xp33_ASAP7_75t_L g1815 ( 
.A1(n_1759),
.A2(n_1686),
.A3(n_1743),
.B1(n_1720),
.B2(n_1730),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1782),
.A2(n_1669),
.B(n_1681),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1758),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1759),
.Y(n_1818)
);

O2A1O1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1782),
.A2(n_1668),
.B(n_1713),
.C(n_1662),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1805),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1797),
.B(n_1765),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1818),
.B(n_1807),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1798),
.B(n_1770),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1795),
.B(n_1759),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1804),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1809),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1811),
.B(n_1792),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1796),
.B(n_1782),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1819),
.B(n_1773),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1803),
.B(n_1779),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1799),
.B(n_1782),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1794),
.B(n_1792),
.Y(n_1832)
);

NAND2x1_ASAP7_75t_L g1833 ( 
.A(n_1812),
.B(n_1773),
.Y(n_1833)
);

OAI21xp33_ASAP7_75t_L g1834 ( 
.A1(n_1815),
.A2(n_1765),
.B(n_1779),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1802),
.B(n_1779),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1806),
.B(n_1765),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1817),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_L g1838 ( 
.A(n_1801),
.B(n_1766),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1808),
.B(n_1777),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_L g1840 ( 
.A(n_1824),
.B(n_1799),
.C(n_1802),
.Y(n_1840)
);

AOI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1824),
.A2(n_1800),
.B(n_1814),
.C(n_1816),
.Y(n_1841)
);

AOI222xp33_ASAP7_75t_L g1842 ( 
.A1(n_1838),
.A2(n_1810),
.B1(n_1813),
.B2(n_1768),
.C1(n_1764),
.C2(n_1776),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1828),
.A2(n_1810),
.B1(n_1764),
.B2(n_1762),
.C(n_1776),
.Y(n_1843)
);

AOI211xp5_ASAP7_75t_L g1844 ( 
.A1(n_1828),
.A2(n_1790),
.B(n_1760),
.C(n_1762),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1834),
.A2(n_1831),
.B1(n_1829),
.B2(n_1823),
.C(n_1820),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1832),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1831),
.A2(n_1788),
.B1(n_1761),
.B2(n_1768),
.C(n_1790),
.Y(n_1847)
);

AOI322xp5_ASAP7_75t_L g1848 ( 
.A1(n_1822),
.A2(n_1792),
.A3(n_1784),
.B1(n_1788),
.B2(n_1761),
.C1(n_1766),
.C2(n_1789),
.Y(n_1848)
);

O2A1O1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1829),
.A2(n_1789),
.B(n_1790),
.C(n_1783),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_L g1850 ( 
.A(n_1821),
.B(n_1773),
.C(n_1763),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1827),
.B(n_1778),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1839),
.B(n_1778),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1833),
.A2(n_1773),
.B(n_1760),
.Y(n_1853)
);

NOR3x1_ASAP7_75t_L g1854 ( 
.A(n_1850),
.B(n_1846),
.C(n_1852),
.Y(n_1854)
);

NOR4xp75_ASAP7_75t_L g1855 ( 
.A(n_1851),
.B(n_1836),
.C(n_1830),
.D(n_1825),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1840),
.A2(n_1835),
.B1(n_1773),
.B2(n_1760),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1845),
.B(n_1826),
.Y(n_1857)
);

NOR3xp33_ASAP7_75t_L g1858 ( 
.A(n_1841),
.B(n_1847),
.C(n_1843),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1848),
.B(n_1778),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1844),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1853),
.Y(n_1861)
);

NOR2x1_ASAP7_75t_L g1862 ( 
.A(n_1849),
.B(n_1837),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1842),
.Y(n_1863)
);

AOI211x1_ASAP7_75t_L g1864 ( 
.A1(n_1850),
.A2(n_1784),
.B(n_1780),
.C(n_1769),
.Y(n_1864)
);

NOR4xp25_ASAP7_75t_L g1865 ( 
.A(n_1845),
.B(n_1763),
.C(n_1785),
.D(n_1775),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_SL g1866 ( 
.A(n_1855),
.B(n_1376),
.C(n_1783),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1858),
.A2(n_1857),
.B1(n_1863),
.B2(n_1865),
.C(n_1856),
.Y(n_1867)
);

NOR3xp33_ASAP7_75t_L g1868 ( 
.A(n_1860),
.B(n_1763),
.C(n_1775),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1865),
.A2(n_1760),
.B(n_1785),
.C(n_1775),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1859),
.B(n_1780),
.Y(n_1870)
);

NOR4xp25_ASAP7_75t_L g1871 ( 
.A(n_1861),
.B(n_1785),
.C(n_1775),
.D(n_1784),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1870),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1867),
.A2(n_1862),
.B1(n_1760),
.B2(n_1780),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1866),
.A2(n_1785),
.B1(n_1771),
.B2(n_1769),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1868),
.A2(n_1771),
.B1(n_1769),
.B2(n_1783),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1871),
.B(n_1854),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1869),
.B(n_1373),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1867),
.A2(n_1771),
.B1(n_1783),
.B2(n_1864),
.Y(n_1878)
);

CKINVDCx6p67_ASAP7_75t_R g1879 ( 
.A(n_1876),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1873),
.A2(n_1713),
.B1(n_1668),
.B2(n_1686),
.C(n_1711),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1872),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1878),
.B(n_1694),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1877),
.Y(n_1883)
);

OAI322xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1874),
.A2(n_1713),
.A3(n_1697),
.B1(n_1696),
.B2(n_1650),
.C1(n_1699),
.C2(n_1706),
.Y(n_1884)
);

NOR3x1_ASAP7_75t_L g1885 ( 
.A(n_1882),
.B(n_1879),
.C(n_1881),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1883),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1880),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1886),
.B(n_1875),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1888),
.B(n_1887),
.C(n_1885),
.Y(n_1889)
);

OAI21x1_ASAP7_75t_SL g1890 ( 
.A1(n_1889),
.A2(n_1373),
.B(n_1884),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1889),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1891),
.A2(n_1416),
.B1(n_1458),
.B2(n_1495),
.Y(n_1892)
);

OAI21x1_ASAP7_75t_L g1893 ( 
.A1(n_1890),
.A2(n_1495),
.B(n_1696),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1892),
.B(n_1495),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1893),
.A2(n_1675),
.B(n_1458),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1894),
.B(n_1416),
.Y(n_1896)
);

OAI222xp33_ASAP7_75t_L g1897 ( 
.A1(n_1896),
.A2(n_1895),
.B1(n_1675),
.B2(n_1707),
.C1(n_1706),
.C2(n_1699),
.Y(n_1897)
);

AOI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1707),
.B1(n_1658),
.B2(n_1647),
.C(n_1649),
.Y(n_1898)
);

AOI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1360),
.B(n_1371),
.C(n_1424),
.Y(n_1899)
);


endmodule