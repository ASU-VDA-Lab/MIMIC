module fake_ibex_439_n_3928 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_658, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3928);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_658;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3928;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_3097;
wire n_2906;
wire n_3030;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_772;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3780;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_1969;
wire n_3798;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3634;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_738;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_2880;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2423;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_669;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_724;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_2999;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_705;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2699;
wire n_2160;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_1115;
wire n_1395;
wire n_998;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_2094;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3880;
wire n_721;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_3034;
wire n_2612;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1694;
wire n_1458;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_3773;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_2732;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_768;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2675;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2348;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_2867;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3576;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_3225;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_3124;
wire n_999;
wire n_2634;
wire n_2982;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_3081;
wire n_2492;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_783;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2148;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2302;
wire n_2560;
wire n_2082;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2619;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_3180;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_866;

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_504),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_518),
.Y(n_668)
);

INVx4_ASAP7_75t_R g669 ( 
.A(n_168),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_126),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_324),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_189),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_428),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_594),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_299),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_0),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_192),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_115),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_296),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_93),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_77),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_538),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_459),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_29),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_270),
.Y(n_685)
);

INVxp33_ASAP7_75t_SL g686 ( 
.A(n_447),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_659),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_473),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_558),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_419),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_511),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_336),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_106),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_145),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_311),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_473),
.Y(n_696)
);

CKINVDCx16_ASAP7_75t_R g697 ( 
.A(n_321),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_229),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_62),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_503),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_158),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_218),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_469),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_173),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_406),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_608),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_553),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_605),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_418),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_421),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_602),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_361),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_482),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_500),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_438),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_609),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_630),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_629),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_647),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_453),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_644),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_238),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_115),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_160),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_640),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_456),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_614),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_593),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_385),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_118),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_604),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_458),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_444),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_645),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_11),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_419),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_522),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_348),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_231),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_120),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_478),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_617),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_306),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_302),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_635),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_327),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_60),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_347),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_598),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_491),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_510),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_497),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_378),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_216),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_124),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_512),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_516),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_498),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_540),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_428),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_296),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_590),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_260),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_592),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_356),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_0),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_380),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_453),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_297),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_224),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_619),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_401),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_316),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_661),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_666),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_497),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_663),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_411),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_443),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_649),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_185),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_578),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_621),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_16),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_41),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_361),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_198),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_637),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_401),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_611),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_600),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_175),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_37),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_73),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_106),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_295),
.Y(n_797)
);

BUFx5_ASAP7_75t_L g798 ( 
.A(n_439),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_350),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_17),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_131),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_394),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_19),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_359),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_90),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_19),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_454),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_189),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_606),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_620),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_58),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_76),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_581),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_622),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_197),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_562),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_481),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_35),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_632),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_664),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_631),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_35),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_484),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_174),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_359),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_138),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_398),
.Y(n_827)
);

BUFx2_ASAP7_75t_SL g828 ( 
.A(n_229),
.Y(n_828)
);

CKINVDCx14_ASAP7_75t_R g829 ( 
.A(n_29),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_83),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_439),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_146),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_251),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_613),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_555),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_535),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_476),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_627),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_564),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_662),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_648),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_612),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_179),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_131),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_646),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_546),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_290),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_651),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_340),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_132),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_47),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_579),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_653),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_23),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_658),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_325),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_352),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_108),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_435),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_267),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_62),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_599),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_323),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_328),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_418),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_449),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_109),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_164),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_245),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_650),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_228),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_149),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_251),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_96),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_618),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_652),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_68),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_641),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_329),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_519),
.Y(n_880)
);

CKINVDCx16_ASAP7_75t_R g881 ( 
.A(n_286),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_125),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_438),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_616),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_413),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_493),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_596),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_166),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_407),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_138),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_657),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_642),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_603),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_542),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_496),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_625),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_404),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_520),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_343),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_364),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_6),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_557),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_332),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_633),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_34),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_51),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_654),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_160),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_410),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_420),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_526),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_308),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_159),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_194),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_499),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_218),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_283),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_554),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_566),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_282),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_533),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_125),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_394),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_31),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_576),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_525),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_121),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_634),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_37),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_230),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_3),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_71),
.Y(n_932)
);

CKINVDCx16_ASAP7_75t_R g933 ( 
.A(n_234),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_95),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_583),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_503),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_468),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_315),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_87),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_199),
.Y(n_940)
);

BUFx5_ASAP7_75t_L g941 ( 
.A(n_41),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_201),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_79),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_515),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_20),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_639),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_431),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_595),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_615),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_90),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_517),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_350),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_344),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_430),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_8),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_434),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_610),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_607),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_187),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_436),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_74),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_312),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_338),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_141),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_409),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_290),
.Y(n_966)
);

CKINVDCx16_ASAP7_75t_R g967 ( 
.A(n_159),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_242),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_660),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_32),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_281),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_414),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_626),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_478),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_156),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_100),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_623),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_588),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_74),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_638),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_482),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_113),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_457),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_283),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_500),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_383),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_85),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_366),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_529),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_572),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_83),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_527),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_114),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_204),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_474),
.Y(n_995)
);

BUFx10_ASAP7_75t_L g996 ( 
.A(n_501),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_45),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_539),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_111),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_413),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_591),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_384),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_445),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_330),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_47),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_387),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_247),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_521),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_335),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_423),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_156),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_147),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_449),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_655),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_168),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_560),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_402),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_457),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_577),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_567),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_321),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_446),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_109),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_227),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_246),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_110),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_101),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_569),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_280),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_534),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_216),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_293),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_376),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_113),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_228),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_149),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_58),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_136),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_132),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_34),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_60),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_226),
.Y(n_1042)
);

BUFx10_ASAP7_75t_L g1043 ( 
.A(n_51),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_323),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_66),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_434),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_366),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_523),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_587),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_103),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_411),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_456),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_73),
.Y(n_1053)
);

CKINVDCx14_ASAP7_75t_R g1054 ( 
.A(n_141),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_258),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_88),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_636),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_380),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_643),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_240),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_80),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_133),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_18),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_86),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_112),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_447),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_423),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_597),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_601),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_563),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_342),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_624),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_388),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_92),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_30),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_87),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_165),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_13),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_334),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_589),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_510),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_341),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_369),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_532),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_48),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_310),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_31),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_400),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_907),
.Y(n_1089)
);

AND2x6_ASAP7_75t_L g1090 ( 
.A(n_809),
.B(n_656),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_907),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_937),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_937),
.B(n_1),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_781),
.B(n_1),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_867),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_937),
.B(n_2),
.Y(n_1096)
);

BUFx12f_ASAP7_75t_L g1097 ( 
.A(n_672),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_829),
.B(n_2),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_798),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_829),
.B(n_3),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_768),
.B(n_4),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_750),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_768),
.B(n_4),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_721),
.B(n_5),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_907),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1076),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_721),
.B(n_5),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_861),
.B(n_6),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_861),
.B(n_7),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1054),
.B(n_7),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_1031),
.B(n_8),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_672),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_798),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1031),
.B(n_9),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_672),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1034),
.B(n_9),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_798),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1034),
.B(n_10),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1054),
.B(n_10),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1044),
.B(n_11),
.Y(n_1120)
);

BUFx8_ASAP7_75t_L g1121 ( 
.A(n_673),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_693),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1044),
.B(n_12),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_907),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_750),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1056),
.B(n_12),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_688),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_853),
.B(n_13),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_859),
.B(n_14),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_798),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_853),
.B(n_14),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_750),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_798),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_688),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_938),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_679),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_726),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1056),
.B(n_15),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_891),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_891),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_726),
.B(n_15),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_918),
.B(n_16),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_688),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_679),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_697),
.B(n_17),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_769),
.B(n_18),
.Y(n_1146)
);

BUFx8_ASAP7_75t_SL g1147 ( 
.A(n_756),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_679),
.Y(n_1148)
);

BUFx8_ASAP7_75t_L g1149 ( 
.A(n_798),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_688),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_720),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_891),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_720),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_698),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_782),
.B(n_20),
.Y(n_1155)
);

BUFx12f_ASAP7_75t_L g1156 ( 
.A(n_713),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_753),
.B(n_21),
.Y(n_1157)
);

INVx5_ASAP7_75t_L g1158 ( 
.A(n_918),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_765),
.B(n_21),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_798),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_720),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_720),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_863),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_723),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_682),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_753),
.B(n_22),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_674),
.B(n_22),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_713),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_723),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_881),
.B(n_23),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_723),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_723),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_698),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_809),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_687),
.Y(n_1175)
);

BUFx8_ASAP7_75t_SL g1176 ( 
.A(n_756),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_837),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_713),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_837),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1088),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_933),
.B(n_24),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_760),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_706),
.B(n_24),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1088),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_722),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_837),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_837),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_716),
.B(n_25),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_675),
.B(n_25),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_676),
.B(n_26),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_777),
.Y(n_1191)
);

BUFx8_ASAP7_75t_SL g1192 ( 
.A(n_758),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_777),
.B(n_26),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_879),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_831),
.B(n_27),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_879),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_831),
.B(n_27),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_879),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_677),
.B(n_28),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_690),
.B(n_28),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_863),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_863),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_870),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_936),
.Y(n_1204)
);

AO22x2_ASAP7_75t_L g1205 ( 
.A1(n_1145),
.A2(n_986),
.B1(n_828),
.B2(n_744),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1146),
.A2(n_747),
.B1(n_812),
.B2(n_696),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1122),
.A2(n_1135),
.B1(n_1173),
.B2(n_1154),
.Y(n_1207)
);

OAI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1094),
.A2(n_967),
.B1(n_686),
.B2(n_668),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1093),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_1097),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1180),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1095),
.A2(n_686),
.B1(n_778),
.B2(n_718),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1184),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1106),
.A2(n_778),
.B1(n_846),
.B2(n_718),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1137),
.B(n_722),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1191),
.B(n_722),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1204),
.B(n_779),
.Y(n_1217)
);

AO22x2_ASAP7_75t_L g1218 ( 
.A1(n_1155),
.A2(n_866),
.B1(n_930),
.B2(n_850),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1174),
.Y(n_1219)
);

AOI22x1_ASAP7_75t_L g1220 ( 
.A1(n_1113),
.A2(n_1019),
.B1(n_727),
.B2(n_728),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1165),
.B(n_1081),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1178),
.B(n_1185),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1178),
.B(n_779),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1185),
.B(n_1102),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1125),
.B(n_779),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_1112),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1094),
.A2(n_787),
.B1(n_794),
.B2(n_758),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1170),
.A2(n_1002),
.B1(n_1047),
.B2(n_953),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1125),
.B(n_799),
.Y(n_1229)
);

AO22x2_ASAP7_75t_L g1230 ( 
.A1(n_1181),
.A2(n_1055),
.B1(n_699),
.B2(n_710),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_1109),
.A2(n_1086),
.B1(n_1082),
.B2(n_705),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1125),
.B(n_799),
.Y(n_1232)
);

NAND3x1_ASAP7_75t_L g1233 ( 
.A(n_1159),
.B(n_794),
.C(n_787),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1129),
.A2(n_875),
.B1(n_904),
.B2(n_846),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1132),
.B(n_799),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_904),
.B1(n_925),
.B2(n_875),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1111),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1203),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1111),
.A2(n_948),
.B1(n_925),
.B2(n_956),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1159),
.A2(n_1101),
.B1(n_1108),
.B2(n_1103),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1092),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1101),
.A2(n_670),
.B1(n_671),
.B2(n_667),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1093),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1182),
.A2(n_1189),
.B1(n_1199),
.B2(n_1190),
.Y(n_1244)
);

OAI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1189),
.A2(n_871),
.B1(n_920),
.B2(n_865),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1114),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_1114),
.A2(n_715),
.B1(n_742),
.B2(n_730),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1147),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_R g1249 ( 
.A1(n_1176),
.A2(n_749),
.B1(n_752),
.B2(n_745),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1103),
.A2(n_678),
.B1(n_681),
.B2(n_680),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1132),
.B(n_807),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1116),
.A2(n_948),
.B1(n_683),
.B2(n_685),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1116),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1108),
.A2(n_684),
.B1(n_692),
.B2(n_691),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1190),
.A2(n_871),
.B1(n_920),
.B2(n_865),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1165),
.B(n_1071),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1132),
.B(n_807),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1118),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1092),
.Y(n_1259)
);

AO22x2_ASAP7_75t_L g1260 ( 
.A1(n_1118),
.A2(n_755),
.B1(n_759),
.B2(n_754),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1126),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1144),
.B(n_766),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_695),
.B1(n_700),
.B2(n_694),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1162),
.Y(n_1264)
);

AO22x2_ASAP7_75t_L g1265 ( 
.A1(n_1138),
.A2(n_1157),
.B1(n_1166),
.B2(n_1141),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1162),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1162),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1138),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1172),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1172),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1139),
.B(n_717),
.Y(n_1271)
);

AO22x2_ASAP7_75t_L g1272 ( 
.A1(n_1141),
.A2(n_1166),
.B1(n_1193),
.B2(n_1157),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1139),
.B(n_807),
.Y(n_1273)
);

OAI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1199),
.A2(n_1018),
.B1(n_1037),
.B2(n_931),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1193),
.A2(n_1197),
.B1(n_1195),
.B2(n_1136),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1115),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1195),
.Y(n_1277)
);

AND2x4_ASAP7_75t_SL g1278 ( 
.A(n_1098),
.B(n_1100),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1148),
.A2(n_1018),
.B1(n_1037),
.B2(n_931),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1197),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1172),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1200),
.A2(n_1078),
.B1(n_780),
.B2(n_785),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1200),
.A2(n_1096),
.B1(n_1123),
.B2(n_1120),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1156),
.B(n_987),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1168),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1120),
.A2(n_701),
.B1(n_703),
.B2(n_702),
.Y(n_1286)
);

OA22x2_ASAP7_75t_L g1287 ( 
.A1(n_1123),
.A2(n_734),
.B1(n_764),
.B2(n_714),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_R g1288 ( 
.A1(n_1192),
.A2(n_786),
.B1(n_800),
.B2(n_770),
.Y(n_1288)
);

AO22x2_ASAP7_75t_L g1289 ( 
.A1(n_1110),
.A2(n_826),
.B1(n_854),
.B2(n_802),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1096),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1186),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_R g1292 ( 
.A1(n_1167),
.A2(n_857),
.B1(n_858),
.B2(n_856),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1119),
.A2(n_709),
.B1(n_712),
.B2(n_704),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1139),
.B(n_732),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1140),
.A2(n_1078),
.B1(n_873),
.B2(n_874),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1140),
.B(n_1152),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1099),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1140),
.A2(n_877),
.B1(n_880),
.B2(n_864),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1089),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1099),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1149),
.A2(n_731),
.B1(n_733),
.B2(n_724),
.Y(n_1301)
);

AO22x2_ASAP7_75t_L g1302 ( 
.A1(n_1131),
.A2(n_886),
.B1(n_889),
.B2(n_885),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1152),
.A2(n_736),
.B1(n_738),
.B2(n_737),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1117),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1186),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1186),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1152),
.A2(n_900),
.B1(n_905),
.B2(n_890),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1175),
.B(n_987),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1117),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1158),
.A2(n_914),
.B1(n_923),
.B2(n_908),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1175),
.B(n_987),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1149),
.A2(n_739),
.B1(n_741),
.B2(n_740),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1104),
.A2(n_751),
.B1(n_757),
.B2(n_748),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1107),
.A2(n_762),
.B1(n_767),
.B2(n_761),
.Y(n_1314)
);

AO22x2_ASAP7_75t_L g1315 ( 
.A1(n_1121),
.A2(n_932),
.B1(n_940),
.B2(n_927),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1196),
.Y(n_1316)
);

AO22x2_ASAP7_75t_L g1317 ( 
.A1(n_1121),
.A2(n_954),
.B1(n_959),
.B2(n_951),
.Y(n_1317)
);

AO22x2_ASAP7_75t_L g1318 ( 
.A1(n_1201),
.A2(n_963),
.B1(n_966),
.B2(n_960),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1089),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1158),
.A2(n_972),
.B1(n_974),
.B2(n_970),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1128),
.A2(n_773),
.B1(n_774),
.B2(n_771),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1183),
.B(n_808),
.Y(n_1322)
);

OA22x2_ASAP7_75t_L g1323 ( 
.A1(n_1201),
.A2(n_830),
.B1(n_849),
.B2(n_796),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1196),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1202),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1158),
.B(n_996),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_R g1327 ( 
.A1(n_1188),
.A2(n_985),
.B1(n_995),
.B2(n_984),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1142),
.A2(n_790),
.B1(n_793),
.B2(n_788),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1202),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1196),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1130),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1133),
.B(n_735),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1160),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1163),
.A2(n_797),
.B1(n_801),
.B2(n_795),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1090),
.A2(n_804),
.B1(n_805),
.B2(n_803),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1090),
.A2(n_811),
.B1(n_815),
.B2(n_806),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1124),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1124),
.A2(n_1011),
.B1(n_1015),
.B2(n_1003),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1124),
.A2(n_1024),
.B1(n_1025),
.B2(n_1023),
.Y(n_1339)
);

AOI22x1_ASAP7_75t_SL g1340 ( 
.A1(n_1090),
.A2(n_817),
.B1(n_822),
.B2(n_818),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1090),
.B(n_996),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1127),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1127),
.A2(n_823),
.B1(n_825),
.B2(n_824),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1127),
.A2(n_827),
.B1(n_833),
.B2(n_832),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1134),
.Y(n_1345)
);

AO22x2_ASAP7_75t_L g1346 ( 
.A1(n_1134),
.A2(n_1040),
.B1(n_1045),
.B2(n_1033),
.Y(n_1346)
);

AND2x2_ASAP7_75t_SL g1347 ( 
.A(n_1134),
.B(n_808),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1143),
.B(n_996),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1143),
.A2(n_847),
.B1(n_851),
.B2(n_844),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1143),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1150),
.A2(n_860),
.B1(n_869),
.B2(n_868),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1150),
.A2(n_882),
.B1(n_883),
.B2(n_872),
.Y(n_1352)
);

NAND2xp33_ASAP7_75t_SL g1353 ( 
.A(n_1150),
.B(n_888),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1151),
.B(n_1043),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1151),
.B(n_1046),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1151),
.A2(n_1058),
.B1(n_1060),
.B2(n_1051),
.Y(n_1356)
);

OR2x6_ASAP7_75t_L g1357 ( 
.A(n_1153),
.B(n_1026),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1153),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1153),
.B(n_1074),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1161),
.A2(n_1062),
.B1(n_1063),
.B2(n_1061),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1161),
.A2(n_897),
.B1(n_898),
.B2(n_895),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1161),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1164),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1164),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1164),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1169),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1169),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1169),
.B(n_1043),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1171),
.A2(n_901),
.B1(n_903),
.B2(n_899),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1171),
.Y(n_1370)
);

INVx8_ASAP7_75t_L g1371 ( 
.A(n_1171),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1177),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1177),
.A2(n_1067),
.B1(n_1073),
.B2(n_1066),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1177),
.B(n_1043),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1179),
.A2(n_909),
.B1(n_910),
.B2(n_906),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1179),
.A2(n_913),
.B1(n_915),
.B2(n_912),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1179),
.A2(n_1085),
.B1(n_1087),
.B2(n_1083),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1187),
.A2(n_968),
.B1(n_1010),
.B2(n_843),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1187),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1187),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1194),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1194),
.A2(n_916),
.B1(n_924),
.B2(n_917),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1194),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1198),
.B(n_936),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1198),
.B(n_945),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1198),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1089),
.A2(n_934),
.B1(n_942),
.B2(n_929),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1091),
.B(n_945),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1091),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1091),
.A2(n_968),
.B1(n_1010),
.B2(n_843),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1105),
.A2(n_943),
.B1(n_947),
.B2(n_944),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1105),
.B(n_863),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1105),
.A2(n_950),
.B1(n_955),
.B2(n_952),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1122),
.A2(n_962),
.B1(n_964),
.B2(n_961),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1097),
.B(n_1026),
.Y(n_1395)
);

AO22x2_ASAP7_75t_L g1396 ( 
.A1(n_1145),
.A2(n_746),
.B1(n_792),
.B2(n_784),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1122),
.A2(n_1075),
.B1(n_1077),
.B2(n_1065),
.Y(n_1397)
);

INVxp67_ASAP7_75t_SL g1398 ( 
.A(n_1149),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1093),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1174),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1174),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1165),
.B(n_1079),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1174),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1093),
.Y(n_1404)
);

OA22x2_ASAP7_75t_L g1405 ( 
.A1(n_1095),
.A2(n_994),
.B1(n_1006),
.B2(n_982),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1094),
.A2(n_965),
.B1(n_975),
.B2(n_971),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1093),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1122),
.A2(n_979),
.B1(n_981),
.B2(n_976),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1094),
.A2(n_983),
.B1(n_991),
.B2(n_988),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1093),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1093),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1097),
.B(n_993),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1122),
.A2(n_999),
.B1(n_1000),
.B2(n_997),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1125),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1174),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1122),
.A2(n_1005),
.B1(n_1007),
.B2(n_1004),
.Y(n_1416)
);

XOR2xp5_ASAP7_75t_L g1417 ( 
.A(n_1212),
.B(n_1009),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1290),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1210),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1211),
.Y(n_1420)
);

XOR2xp5_ASAP7_75t_L g1421 ( 
.A(n_1214),
.B(n_1012),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1222),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1213),
.B(n_1013),
.Y(n_1423)
);

XOR2xp5_ASAP7_75t_L g1424 ( 
.A(n_1234),
.B(n_1017),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1388),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1237),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1388),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1246),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1253),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1268),
.Y(n_1430)
);

XOR2xp5_ASAP7_75t_L g1431 ( 
.A(n_1340),
.B(n_1048),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1355),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1283),
.B(n_941),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1241),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1259),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1265),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1265),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1348),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1354),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1395),
.B(n_879),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1368),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1217),
.B(n_1021),
.Y(n_1442)
);

BUFx5_ASAP7_75t_L g1443 ( 
.A(n_1331),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1385),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1279),
.Y(n_1445)
);

XOR2xp5_ASAP7_75t_L g1446 ( 
.A(n_1236),
.B(n_1050),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1357),
.Y(n_1447)
);

CKINVDCx16_ASAP7_75t_R g1448 ( 
.A(n_1284),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1374),
.Y(n_1449)
);

XOR2xp5_ASAP7_75t_L g1450 ( 
.A(n_1248),
.B(n_1239),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1258),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1261),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1272),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1272),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1221),
.B(n_839),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1226),
.B(n_1053),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1209),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1243),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1285),
.Y(n_1459)
);

XOR2xp5_ASAP7_75t_L g1460 ( 
.A(n_1207),
.B(n_1064),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1399),
.Y(n_1461)
);

XOR2xp5_ASAP7_75t_L g1462 ( 
.A(n_1315),
.B(n_1022),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1404),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1407),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1410),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1411),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1385),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1318),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1276),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1335),
.B(n_528),
.Y(n_1470)
);

AOI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1297),
.A2(n_819),
.B(n_814),
.Y(n_1471)
);

AND2x6_ASAP7_75t_L g1472 ( 
.A(n_1341),
.B(n_870),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1318),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1384),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1395),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1215),
.B(n_1027),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1300),
.A2(n_836),
.B(n_835),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1240),
.B(n_689),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1346),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1278),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1216),
.B(n_1029),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1346),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1231),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1231),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1247),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1252),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1247),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1260),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1260),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1277),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1304),
.A2(n_848),
.B(n_838),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1390),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1280),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1359),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1390),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1256),
.B(n_973),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1392),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1402),
.B(n_1028),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1394),
.B(n_1408),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1378),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1413),
.B(n_1032),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1416),
.B(n_1035),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1366),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1378),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1219),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1308),
.B(n_707),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1366),
.Y(n_1507)
);

XNOR2x2_ASAP7_75t_L g1508 ( 
.A(n_1230),
.B(n_1206),
.Y(n_1508)
);

HAxp5_ASAP7_75t_SL g1509 ( 
.A(n_1249),
.B(n_892),
.CON(n_1509),
.SN(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1238),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1400),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1401),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1403),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1397),
.B(n_1244),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1415),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1301),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1398),
.B(n_1038),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1311),
.B(n_1039),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1223),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1264),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1224),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1262),
.Y(n_1522)
);

INVxp67_ASAP7_75t_SL g1523 ( 
.A(n_1309),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1289),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1412),
.B(n_922),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1245),
.B(n_1041),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1289),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1302),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1293),
.B(n_1052),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1302),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1275),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1296),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1325),
.A2(n_902),
.B(n_894),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1323),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1396),
.B(n_863),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1357),
.Y(n_1536)
);

INVxp33_ASAP7_75t_L g1537 ( 
.A(n_1206),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1225),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1229),
.Y(n_1539)
);

XNOR2x2_ASAP7_75t_L g1540 ( 
.A(n_1230),
.B(n_1218),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1232),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1329),
.B(n_863),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_SL g1543 ( 
.A(n_1322),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_R g1544 ( 
.A(n_1322),
.B(n_708),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1332),
.B(n_941),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1235),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1312),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1251),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1326),
.Y(n_1549)
);

XOR2x2_ASAP7_75t_L g1550 ( 
.A(n_1233),
.B(n_30),
.Y(n_1550)
);

XNOR2x1_ASAP7_75t_L g1551 ( 
.A(n_1315),
.B(n_32),
.Y(n_1551)
);

XOR2xp5_ASAP7_75t_L g1552 ( 
.A(n_1317),
.B(n_33),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1257),
.B(n_1030),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1273),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1396),
.B(n_863),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1287),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1414),
.B(n_711),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1356),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1360),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1220),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1205),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1205),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1338),
.Y(n_1563)
);

INVxp33_ASAP7_75t_L g1564 ( 
.A(n_1218),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1263),
.B(n_719),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1313),
.B(n_941),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1339),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1310),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1320),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1344),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1314),
.B(n_725),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1321),
.B(n_729),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1382),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1334),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1317),
.B(n_922),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1303),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1391),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1393),
.Y(n_1578)
);

INVxp33_ASAP7_75t_L g1579 ( 
.A(n_1228),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1349),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1352),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1361),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1375),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1328),
.B(n_941),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1266),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1271),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1294),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1298),
.B(n_743),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1387),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1405),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1343),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1267),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1351),
.Y(n_1593)
);

XOR2xp5_ASAP7_75t_L g1594 ( 
.A(n_1227),
.B(n_33),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1228),
.B(n_1369),
.Y(n_1595)
);

INVx8_ASAP7_75t_L g1596 ( 
.A(n_1371),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1269),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1249),
.B(n_922),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1376),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1307),
.B(n_763),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1347),
.B(n_941),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1336),
.B(n_941),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1242),
.B(n_772),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1333),
.Y(n_1604)
);

AND2x2_ASAP7_75t_SL g1605 ( 
.A(n_1255),
.B(n_1274),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1270),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1282),
.B(n_941),
.Y(n_1607)
);

XOR2xp5_ASAP7_75t_L g1608 ( 
.A(n_1208),
.B(n_36),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1281),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_R g1610 ( 
.A(n_1288),
.B(n_775),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1250),
.A2(n_1286),
.B(n_1254),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1291),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1305),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1306),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1373),
.B(n_911),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1316),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1353),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1324),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1288),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1406),
.B(n_776),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1330),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1337),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1377),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1409),
.B(n_1068),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1292),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1295),
.B(n_1068),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1292),
.B(n_922),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1327),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1371),
.B(n_921),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1327),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1364),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1379),
.B(n_939),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1342),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_SL g1634 ( 
.A(n_1345),
.B(n_783),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1350),
.Y(n_1635)
);

NAND2xp33_ASAP7_75t_SL g1636 ( 
.A(n_1299),
.B(n_939),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1362),
.B(n_939),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1363),
.B(n_957),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1367),
.Y(n_1639)
);

XOR2x2_ASAP7_75t_L g1640 ( 
.A(n_1372),
.B(n_36),
.Y(n_1640)
);

INVx4_ASAP7_75t_SL g1641 ( 
.A(n_1319),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1381),
.A2(n_977),
.B(n_969),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1319),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1386),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1358),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1299),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1365),
.B(n_789),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1370),
.B(n_939),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1380),
.B(n_1008),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1383),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1389),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1319),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1290),
.Y(n_1653)
);

XOR2xp5_ASAP7_75t_L g1654 ( 
.A(n_1212),
.B(n_38),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1290),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1290),
.B(n_978),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1388),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1290),
.B(n_791),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1290),
.Y(n_1659)
);

CKINVDCx16_ASAP7_75t_R g1660 ( 
.A(n_1210),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1388),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1290),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1290),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1290),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_L g1665 ( 
.A(n_1290),
.B(n_541),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1290),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1290),
.B(n_980),
.Y(n_1667)
);

AND2x2_ASAP7_75t_SL g1668 ( 
.A(n_1210),
.B(n_1008),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1390),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1290),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1290),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1290),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1290),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1290),
.Y(n_1674)
);

XNOR2x2_ASAP7_75t_L g1675 ( 
.A(n_1230),
.B(n_669),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1290),
.B(n_810),
.Y(n_1676)
);

XOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1212),
.B(n_38),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1357),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1290),
.B(n_813),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1290),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1290),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1388),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1290),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1290),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1212),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_1212),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1290),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1211),
.Y(n_1688)
);

XOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1212),
.B(n_39),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1283),
.B(n_816),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1290),
.B(n_989),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1290),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1290),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1290),
.Y(n_1694)
);

XOR2x2_ASAP7_75t_L g1695 ( 
.A(n_1279),
.B(n_39),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1290),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1290),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1388),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1290),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1211),
.B(n_1008),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1388),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1388),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1290),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1290),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1388),
.Y(n_1705)
);

INVxp33_ASAP7_75t_L g1706 ( 
.A(n_1212),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1290),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1357),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1290),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1290),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1388),
.Y(n_1711)
);

XOR2x2_ASAP7_75t_L g1712 ( 
.A(n_1279),
.B(n_40),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1290),
.B(n_820),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1388),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1418),
.B(n_821),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1673),
.B(n_1014),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1688),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1420),
.B(n_1008),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1420),
.B(n_1036),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1459),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1443),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1596),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1596),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1653),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1655),
.B(n_1036),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1596),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1659),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1443),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1443),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1662),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1447),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1423),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1663),
.B(n_1036),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1664),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1666),
.B(n_834),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1670),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_1419),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1443),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1665),
.A2(n_1059),
.B(n_1057),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1671),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1443),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1672),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1674),
.B(n_840),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1447),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1665),
.B(n_1069),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1700),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1680),
.B(n_841),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1447),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1681),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1434),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1435),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1678),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1683),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1684),
.B(n_842),
.Y(n_1754)
);

NAND2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1678),
.B(n_1036),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1678),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1522),
.B(n_1042),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1479),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1648),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1433),
.A2(n_1080),
.B(n_1072),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1708),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1456),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1440),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1708),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1687),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1692),
.B(n_1042),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1693),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1574),
.B(n_1084),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1694),
.B(n_1696),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1697),
.B(n_1042),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1699),
.B(n_845),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1469),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1440),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1703),
.B(n_1704),
.Y(n_1774)
);

AND2x2_ASAP7_75t_SL g1775 ( 
.A(n_1525),
.B(n_1042),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1707),
.B(n_1019),
.Y(n_1776)
);

INVx3_ASAP7_75t_SL g1777 ( 
.A(n_1660),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1709),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1574),
.B(n_1710),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1708),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1426),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1497),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1523),
.B(n_40),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1436),
.B(n_42),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1605),
.B(n_42),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1433),
.A2(n_855),
.B(n_852),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1625),
.B(n_43),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1440),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1417),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1637),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1637),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1654),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1677),
.Y(n_1793)
);

INVx6_ASAP7_75t_L g1794 ( 
.A(n_1475),
.Y(n_1794)
);

AND2x2_ASAP7_75t_SL g1795 ( 
.A(n_1482),
.B(n_43),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1523),
.B(n_1656),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1560),
.A2(n_876),
.B(n_862),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1646),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1478),
.B(n_1531),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1656),
.B(n_878),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1689),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1517),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1514),
.B(n_44),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1589),
.B(n_884),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1667),
.B(n_887),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1575),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1428),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1575),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1667),
.B(n_893),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1691),
.B(n_1519),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1691),
.B(n_44),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1451),
.B(n_896),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1575),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1524),
.B(n_45),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1480),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1452),
.B(n_919),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1477),
.A2(n_928),
.B(n_926),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1480),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1425),
.Y(n_1819)
);

AND2x2_ASAP7_75t_SL g1820 ( 
.A(n_1448),
.B(n_46),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1668),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1527),
.B(n_1492),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1646),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1457),
.B(n_935),
.Y(n_1824)
);

NAND2x1p5_ASAP7_75t_L g1825 ( 
.A(n_1437),
.B(n_46),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1492),
.B(n_1495),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1429),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1685),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1649),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1430),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1504),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1591),
.B(n_946),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1422),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1458),
.B(n_949),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1521),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1468),
.B(n_958),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1438),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1504),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1508),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1593),
.B(n_990),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1495),
.B(n_48),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1461),
.B(n_992),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1599),
.B(n_998),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1543),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1669),
.B(n_49),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1669),
.B(n_49),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1540),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1474),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1463),
.B(n_1001),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1471),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1464),
.B(n_1016),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1427),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1686),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1646),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1473),
.B(n_50),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1444),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1535),
.B(n_50),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1465),
.B(n_1020),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1442),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1555),
.B(n_52),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1467),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1657),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1439),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1661),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1682),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1483),
.B(n_52),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1698),
.Y(n_1867)
);

INVx5_ASAP7_75t_L g1868 ( 
.A(n_1472),
.Y(n_1868)
);

AND2x2_ASAP7_75t_SL g1869 ( 
.A(n_1500),
.B(n_53),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1484),
.B(n_53),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1701),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1441),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1449),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1702),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1628),
.B(n_54),
.Y(n_1875)
);

AND2x2_ASAP7_75t_SL g1876 ( 
.A(n_1562),
.B(n_54),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1705),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1630),
.B(n_55),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1477),
.A2(n_1070),
.B(n_1049),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1466),
.B(n_55),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1706),
.B(n_56),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1432),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1472),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1711),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1460),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1526),
.B(n_56),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1714),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1490),
.Y(n_1888)
);

AND2x2_ASAP7_75t_SL g1889 ( 
.A(n_1485),
.B(n_57),
.Y(n_1889)
);

INVx4_ASAP7_75t_L g1890 ( 
.A(n_1472),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1503),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1493),
.B(n_57),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1658),
.B(n_59),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1542),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1487),
.B(n_59),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1488),
.B(n_61),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1491),
.A2(n_530),
.B(n_524),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1542),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1520),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1585),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1518),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1536),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1489),
.B(n_61),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1592),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1538),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1675),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1453),
.B(n_63),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1676),
.B(n_63),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1679),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1454),
.B(n_64),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1597),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1470),
.B(n_531),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1594),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1539),
.B(n_64),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1713),
.B(n_65),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1633),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1541),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1635),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1626),
.Y(n_1919)
);

BUFx4_ASAP7_75t_SL g1920 ( 
.A(n_1598),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1639),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1626),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1598),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1546),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1507),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1476),
.B(n_65),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1568),
.B(n_66),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1481),
.B(n_67),
.Y(n_1928)
);

NAND2x1p5_ASAP7_75t_L g1929 ( 
.A(n_1528),
.B(n_67),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1510),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1548),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1644),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1627),
.B(n_1569),
.Y(n_1933)
);

INVx4_ASAP7_75t_L g1934 ( 
.A(n_1472),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1532),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1566),
.B(n_68),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1606),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1584),
.B(n_69),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1607),
.B(n_69),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1563),
.B(n_70),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1491),
.B(n_70),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1494),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1505),
.Y(n_1943)
);

BUFx2_ASAP7_75t_L g1944 ( 
.A(n_1598),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1421),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1543),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1629),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1424),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1609),
.Y(n_1949)
);

BUFx5_ASAP7_75t_L g1950 ( 
.A(n_1652),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1533),
.B(n_1567),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_R g1952 ( 
.A(n_1544),
.B(n_1486),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1623),
.B(n_1690),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1558),
.B(n_71),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1612),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1446),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1534),
.B(n_72),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1511),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1512),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1513),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1613),
.Y(n_1961)
);

AND2x6_ASAP7_75t_L g1962 ( 
.A(n_1530),
.B(n_1601),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1559),
.B(n_72),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1533),
.B(n_75),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1595),
.B(n_75),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1614),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1602),
.B(n_76),
.Y(n_1967)
);

BUFx12f_ASAP7_75t_SL g1968 ( 
.A(n_1624),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1616),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1618),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1515),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1554),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1537),
.B(n_77),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1621),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1604),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1549),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1550),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1695),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1622),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1586),
.A2(n_537),
.B(n_536),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1712),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1564),
.B(n_78),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1579),
.B(n_78),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1529),
.B(n_79),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1499),
.B(n_80),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1577),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1553),
.B(n_81),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1501),
.B(n_81),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1553),
.B(n_82),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1502),
.B(n_82),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1561),
.B(n_84),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1643),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1643),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1629),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1565),
.B(n_84),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1632),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1455),
.B(n_85),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1624),
.B(n_1556),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1578),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1645),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1496),
.B(n_86),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1580),
.B(n_88),
.Y(n_2002)
);

INVxp67_ASAP7_75t_L g2003 ( 
.A(n_1590),
.Y(n_2003)
);

OAI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1587),
.A2(n_544),
.B(n_543),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1570),
.B(n_89),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1573),
.B(n_89),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1650),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1638),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1581),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1498),
.B(n_91),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1506),
.B(n_91),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1582),
.B(n_92),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1583),
.B(n_1611),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1638),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1462),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1651),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1611),
.B(n_93),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1470),
.B(n_1642),
.Y(n_2018)
);

AND2x6_ASAP7_75t_L g2019 ( 
.A(n_1617),
.B(n_545),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1615),
.Y(n_2020)
);

INVxp67_ASAP7_75t_SL g2021 ( 
.A(n_1450),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1620),
.B(n_94),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1603),
.B(n_94),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1641),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1571),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1615),
.B(n_1572),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1642),
.A2(n_1545),
.B(n_1647),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1588),
.B(n_97),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1641),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1617),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1631),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1600),
.B(n_98),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1545),
.B(n_98),
.Y(n_2033)
);

CKINVDCx20_ASAP7_75t_R g2034 ( 
.A(n_1576),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1557),
.B(n_99),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1608),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1634),
.B(n_99),
.Y(n_2037)
);

NOR2xp67_ASAP7_75t_R g2038 ( 
.A(n_1610),
.B(n_100),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_SL g2039 ( 
.A(n_1516),
.B(n_101),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1551),
.B(n_102),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1634),
.B(n_665),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1552),
.B(n_102),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1547),
.B(n_103),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1640),
.B(n_104),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1431),
.B(n_104),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1445),
.B(n_105),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1619),
.B(n_105),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1636),
.Y(n_2048)
);

NAND2x1p5_ASAP7_75t_L g2049 ( 
.A(n_1509),
.B(n_107),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1443),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1418),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1418),
.B(n_107),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1418),
.B(n_108),
.Y(n_2053)
);

AND2x4_ASAP7_75t_SL g2054 ( 
.A(n_1440),
.B(n_110),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1596),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1726),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1796),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1779),
.B(n_111),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1778),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1779),
.B(n_112),
.Y(n_2060)
);

INVx4_ASAP7_75t_L g2061 ( 
.A(n_1726),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1769),
.B(n_114),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1778),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1769),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_SL g2065 ( 
.A(n_1883),
.B(n_547),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1798),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1774),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1774),
.B(n_116),
.Y(n_2068)
);

CKINVDCx16_ASAP7_75t_R g2069 ( 
.A(n_1737),
.Y(n_2069)
);

OR2x6_ASAP7_75t_L g2070 ( 
.A(n_1726),
.B(n_116),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1951),
.B(n_117),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_1717),
.Y(n_2072)
);

OR2x6_ASAP7_75t_L g2073 ( 
.A(n_1726),
.B(n_117),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_2055),
.B(n_118),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1951),
.B(n_119),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1762),
.B(n_119),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1942),
.B(n_120),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1770),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1947),
.B(n_121),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1798),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1798),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1901),
.B(n_122),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_2055),
.B(n_122),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2026),
.B(n_123),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1720),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1732),
.B(n_123),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1859),
.B(n_124),
.Y(n_2087)
);

BUFx12f_ASAP7_75t_L g2088 ( 
.A(n_1844),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1828),
.B(n_126),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1722),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1994),
.B(n_127),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_1853),
.B(n_127),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1985),
.B(n_128),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1770),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1798),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_1777),
.Y(n_2096)
);

NAND2x1p5_ASAP7_75t_L g2097 ( 
.A(n_1722),
.B(n_128),
.Y(n_2097)
);

OR2x6_ASAP7_75t_L g2098 ( 
.A(n_1723),
.B(n_129),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1724),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_SL g2100 ( 
.A(n_1883),
.B(n_548),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1810),
.B(n_129),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_1788),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1823),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1737),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_2051),
.B(n_130),
.Y(n_2105)
);

INVx3_ASAP7_75t_L g2106 ( 
.A(n_1748),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1727),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1985),
.B(n_130),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_SL g2109 ( 
.A(n_1883),
.B(n_549),
.Y(n_2109)
);

INVx5_ASAP7_75t_L g2110 ( 
.A(n_1723),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1770),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1777),
.B(n_133),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1730),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1734),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1736),
.B(n_134),
.Y(n_2115)
);

NAND2x1p5_ASAP7_75t_L g2116 ( 
.A(n_1788),
.B(n_1731),
.Y(n_2116)
);

BUFx5_ASAP7_75t_L g2117 ( 
.A(n_1744),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_1885),
.B(n_134),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1740),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1742),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2054),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1749),
.B(n_135),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1753),
.Y(n_2123)
);

OR2x6_ASAP7_75t_L g2124 ( 
.A(n_1923),
.B(n_135),
.Y(n_2124)
);

BUFx4_ASAP7_75t_SL g2125 ( 
.A(n_1844),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1748),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2054),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_SL g2128 ( 
.A(n_1890),
.B(n_550),
.Y(n_2128)
);

BUFx12f_ASAP7_75t_L g2129 ( 
.A(n_1794),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1765),
.B(n_136),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1767),
.B(n_137),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1799),
.B(n_137),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1933),
.B(n_139),
.Y(n_2133)
);

AND2x6_ASAP7_75t_L g2134 ( 
.A(n_1784),
.B(n_139),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1888),
.Y(n_2135)
);

BUFx8_ASAP7_75t_SL g2136 ( 
.A(n_1906),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1750),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1933),
.B(n_140),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1799),
.B(n_140),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1750),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1820),
.B(n_1802),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1751),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1986),
.B(n_1999),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1751),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2013),
.B(n_142),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1725),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_1794),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2013),
.B(n_142),
.Y(n_2148)
);

INVx5_ASAP7_75t_L g2149 ( 
.A(n_1731),
.Y(n_2149)
);

BUFx12f_ASAP7_75t_L g2150 ( 
.A(n_1794),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1894),
.Y(n_2151)
);

INVx2_ASAP7_75t_SL g2152 ( 
.A(n_1920),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1725),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1733),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1820),
.B(n_1746),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1894),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1823),
.Y(n_2157)
);

BUFx3_ASAP7_75t_L g2158 ( 
.A(n_1744),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_1731),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1733),
.Y(n_2160)
);

BUFx4f_ASAP7_75t_L g2161 ( 
.A(n_1889),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2020),
.B(n_143),
.Y(n_2162)
);

NAND2x1_ASAP7_75t_SL g2163 ( 
.A(n_1789),
.B(n_143),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1986),
.B(n_144),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1783),
.B(n_144),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_1909),
.B(n_145),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1898),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1766),
.Y(n_2168)
);

BUFx12f_ASAP7_75t_L g2169 ( 
.A(n_2049),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1783),
.B(n_146),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_1913),
.B(n_147),
.Y(n_2171)
);

INVx4_ASAP7_75t_L g2172 ( 
.A(n_1761),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_1999),
.B(n_148),
.Y(n_2173)
);

BUFx2_ASAP7_75t_SL g2174 ( 
.A(n_1761),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_1773),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_1772),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_SL g2177 ( 
.A(n_1890),
.B(n_551),
.Y(n_2177)
);

NAND2x1p5_ASAP7_75t_L g2178 ( 
.A(n_1815),
.B(n_148),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_2009),
.B(n_150),
.Y(n_2179)
);

OR2x6_ASAP7_75t_L g2180 ( 
.A(n_1944),
.B(n_150),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_1988),
.B(n_151),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1823),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1898),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1748),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_2009),
.B(n_151),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_1968),
.B(n_152),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_1988),
.B(n_152),
.Y(n_2187)
);

BUFx12f_ASAP7_75t_L g2188 ( 
.A(n_2049),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1775),
.B(n_153),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_1818),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_1990),
.B(n_153),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1882),
.B(n_154),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_1945),
.B(n_154),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1823),
.Y(n_2194)
);

BUFx8_ASAP7_75t_L g2195 ( 
.A(n_2042),
.Y(n_2195)
);

AO21x2_ASAP7_75t_L g2196 ( 
.A1(n_1739),
.A2(n_556),
.B(n_552),
.Y(n_2196)
);

BUFx12f_ASAP7_75t_L g2197 ( 
.A(n_1957),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1998),
.B(n_155),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1768),
.B(n_155),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2008),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2014),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1916),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_SL g2203 ( 
.A(n_1890),
.B(n_559),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1998),
.B(n_157),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1833),
.B(n_157),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1990),
.B(n_158),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1766),
.Y(n_2207)
);

OR2x6_ASAP7_75t_L g2208 ( 
.A(n_1946),
.B(n_161),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1768),
.B(n_161),
.Y(n_2209)
);

AND2x6_ASAP7_75t_L g2210 ( 
.A(n_1784),
.B(n_2002),
.Y(n_2210)
);

BUFx2_ASAP7_75t_L g2211 ( 
.A(n_2034),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_1902),
.B(n_162),
.Y(n_2212)
);

INVx6_ASAP7_75t_L g2213 ( 
.A(n_1848),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1916),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_1752),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1811),
.B(n_162),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1918),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1918),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1752),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1984),
.B(n_163),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1921),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1811),
.B(n_163),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1921),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1803),
.B(n_164),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1902),
.B(n_165),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1854),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1984),
.B(n_166),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1803),
.B(n_167),
.Y(n_2228)
);

BUFx12f_ASAP7_75t_L g2229 ( 
.A(n_1957),
.Y(n_2229)
);

AND2x2_ASAP7_75t_SL g2230 ( 
.A(n_1775),
.B(n_167),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1759),
.Y(n_2231)
);

NOR2xp67_ASAP7_75t_L g2232 ( 
.A(n_1934),
.B(n_1868),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1932),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_1934),
.B(n_1822),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1759),
.Y(n_2235)
);

AND2x2_ASAP7_75t_SL g2236 ( 
.A(n_1876),
.B(n_1889),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1835),
.B(n_169),
.Y(n_2237)
);

BUFx3_ASAP7_75t_L g2238 ( 
.A(n_1752),
.Y(n_2238)
);

NAND2x1p5_ASAP7_75t_L g2239 ( 
.A(n_1756),
.B(n_169),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1764),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1932),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1905),
.B(n_170),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_1934),
.B(n_170),
.Y(n_2243)
);

NAND2x1p5_ASAP7_75t_L g2244 ( 
.A(n_1756),
.B(n_171),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1917),
.B(n_171),
.Y(n_2245)
);

CKINVDCx6p67_ASAP7_75t_R g2246 ( 
.A(n_1914),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1854),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_1822),
.B(n_172),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1876),
.B(n_172),
.Y(n_2249)
);

BUFx8_ASAP7_75t_SL g2250 ( 
.A(n_2034),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_1848),
.B(n_173),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1924),
.B(n_1931),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_1935),
.B(n_174),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1968),
.B(n_175),
.Y(n_2254)
);

BUFx3_ASAP7_75t_L g2255 ( 
.A(n_1764),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1804),
.B(n_176),
.Y(n_2256)
);

OR2x6_ASAP7_75t_L g2257 ( 
.A(n_1957),
.B(n_176),
.Y(n_2257)
);

OR2x6_ASAP7_75t_L g2258 ( 
.A(n_2002),
.B(n_177),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_1837),
.B(n_177),
.Y(n_2259)
);

AND2x6_ASAP7_75t_L g2260 ( 
.A(n_1784),
.B(n_2002),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1937),
.Y(n_2261)
);

BUFx8_ASAP7_75t_SL g2262 ( 
.A(n_2047),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1804),
.B(n_178),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_1764),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_1832),
.B(n_1840),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1856),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_1863),
.B(n_1872),
.Y(n_2267)
);

BUFx2_ASAP7_75t_SL g2268 ( 
.A(n_1914),
.Y(n_2268)
);

BUFx2_ASAP7_75t_L g2269 ( 
.A(n_1763),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_1919),
.B(n_178),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_1873),
.B(n_179),
.Y(n_2271)
);

NAND2x1p5_ASAP7_75t_L g2272 ( 
.A(n_1780),
.B(n_180),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1854),
.Y(n_2273)
);

NAND2x1p5_ASAP7_75t_L g2274 ( 
.A(n_1780),
.B(n_180),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1922),
.B(n_2040),
.Y(n_2275)
);

CKINVDCx8_ASAP7_75t_R g2276 ( 
.A(n_1914),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2044),
.B(n_181),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_1926),
.B(n_1928),
.Y(n_2278)
);

CKINVDCx16_ASAP7_75t_R g2279 ( 
.A(n_1952),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1886),
.B(n_181),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1856),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1937),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1832),
.B(n_182),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1862),
.Y(n_2284)
);

BUFx4f_ASAP7_75t_L g2285 ( 
.A(n_1795),
.Y(n_2285)
);

INVxp67_ASAP7_75t_L g2286 ( 
.A(n_2039),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_1780),
.B(n_182),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1738),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1862),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1840),
.B(n_183),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_1948),
.B(n_183),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_1831),
.Y(n_2292)
);

INVx4_ASAP7_75t_L g2293 ( 
.A(n_1854),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_1956),
.B(n_1792),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1864),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1864),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_1891),
.B(n_184),
.Y(n_2297)
);

BUFx3_ASAP7_75t_L g2298 ( 
.A(n_1891),
.Y(n_2298)
);

BUFx4f_ASAP7_75t_L g2299 ( 
.A(n_1795),
.Y(n_2299)
);

BUFx12f_ASAP7_75t_L g2300 ( 
.A(n_2047),
.Y(n_2300)
);

NAND2x1p5_ASAP7_75t_L g2301 ( 
.A(n_1821),
.B(n_1868),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_1925),
.B(n_184),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1843),
.B(n_1995),
.Y(n_2303)
);

BUFx4f_ASAP7_75t_L g2304 ( 
.A(n_1869),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_1868),
.B(n_185),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1949),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_1843),
.B(n_186),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1949),
.Y(n_2308)
);

BUFx3_ASAP7_75t_L g2309 ( 
.A(n_1925),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1941),
.B(n_186),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_L g2311 ( 
.A(n_1972),
.B(n_187),
.Y(n_2311)
);

NAND2x1_ASAP7_75t_SL g2312 ( 
.A(n_1941),
.B(n_188),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_1976),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1964),
.B(n_188),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1955),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_1793),
.B(n_190),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_1965),
.B(n_190),
.Y(n_2317)
);

BUFx4f_ASAP7_75t_L g2318 ( 
.A(n_1869),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1964),
.B(n_191),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_1801),
.B(n_191),
.Y(n_2320)
);

INVx4_ASAP7_75t_L g2321 ( 
.A(n_1868),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_SL g2322 ( 
.A(n_1806),
.B(n_561),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1955),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_SL g2324 ( 
.A(n_1808),
.B(n_565),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2043),
.B(n_192),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_1718),
.Y(n_2326)
);

OR2x2_ASAP7_75t_L g2327 ( 
.A(n_2021),
.B(n_193),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_1965),
.B(n_193),
.Y(n_2328)
);

BUFx12f_ASAP7_75t_L g2329 ( 
.A(n_1825),
.Y(n_2329)
);

BUFx3_ASAP7_75t_L g2330 ( 
.A(n_1718),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1969),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1969),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_SL g2333 ( 
.A(n_1813),
.B(n_568),
.Y(n_2333)
);

AND2x4_ASAP7_75t_L g2334 ( 
.A(n_1781),
.B(n_194),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1979),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1871),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_1787),
.B(n_195),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1875),
.B(n_195),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_1878),
.B(n_196),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_1738),
.Y(n_2340)
);

NOR2x1_ASAP7_75t_L g2341 ( 
.A(n_1912),
.B(n_196),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_1939),
.B(n_197),
.Y(n_2342)
);

BUFx12f_ASAP7_75t_L g2343 ( 
.A(n_1825),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1738),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2003),
.B(n_198),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_1979),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1939),
.B(n_1716),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2050),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1716),
.B(n_199),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1881),
.B(n_200),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1871),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1874),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_SL g2353 ( 
.A(n_1868),
.B(n_570),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1874),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2050),
.Y(n_2355)
);

NAND2x1p5_ASAP7_75t_L g2356 ( 
.A(n_1966),
.B(n_200),
.Y(n_2356)
);

INVx4_ASAP7_75t_L g2357 ( 
.A(n_1755),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2022),
.B(n_201),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1899),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_1807),
.B(n_202),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_SL g2361 ( 
.A(n_1826),
.B(n_571),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2022),
.B(n_202),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1899),
.Y(n_2363)
);

AND2x6_ASAP7_75t_L g2364 ( 
.A(n_1826),
.B(n_203),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_1877),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_1838),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1877),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1884),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2023),
.B(n_203),
.Y(n_2369)
);

CKINVDCx20_ASAP7_75t_R g2370 ( 
.A(n_1952),
.Y(n_2370)
);

INVx4_ASAP7_75t_L g2371 ( 
.A(n_1755),
.Y(n_2371)
);

BUFx12f_ASAP7_75t_L g2372 ( 
.A(n_1929),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2023),
.B(n_204),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1900),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_1836),
.B(n_205),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2015),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1884),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_1719),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_1978),
.B(n_1981),
.Y(n_2379)
);

INVx6_ASAP7_75t_L g2380 ( 
.A(n_1719),
.Y(n_2380)
);

NAND2x1p5_ASAP7_75t_L g2381 ( 
.A(n_1966),
.B(n_205),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1900),
.Y(n_2382)
);

NAND2xp33_ASAP7_75t_L g2383 ( 
.A(n_2019),
.B(n_573),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1953),
.B(n_206),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1904),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_1977),
.B(n_1785),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_1839),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_2050),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_1827),
.B(n_206),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_1836),
.B(n_207),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_1927),
.B(n_207),
.Y(n_2391)
);

BUFx2_ASAP7_75t_L g2392 ( 
.A(n_1758),
.Y(n_2392)
);

BUFx3_ASAP7_75t_L g2393 ( 
.A(n_2024),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_SL g2394 ( 
.A(n_2019),
.B(n_574),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2046),
.B(n_208),
.Y(n_2395)
);

OR2x2_ASAP7_75t_L g2396 ( 
.A(n_2036),
.B(n_208),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_1830),
.B(n_209),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2028),
.B(n_209),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_1975),
.B(n_1814),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2032),
.B(n_210),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_SL g2401 ( 
.A(n_2019),
.B(n_575),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1927),
.B(n_210),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2017),
.B(n_211),
.Y(n_2403)
);

BUFx2_ASAP7_75t_L g2404 ( 
.A(n_1841),
.Y(n_2404)
);

BUFx12f_ASAP7_75t_L g2405 ( 
.A(n_1929),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2046),
.B(n_211),
.Y(n_2406)
);

BUFx2_ASAP7_75t_L g2407 ( 
.A(n_1841),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2017),
.B(n_2012),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1904),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_1847),
.B(n_212),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_1782),
.B(n_212),
.Y(n_2411)
);

NAND2x1p5_ASAP7_75t_L g2412 ( 
.A(n_1782),
.B(n_213),
.Y(n_2412)
);

OR2x6_ASAP7_75t_L g2413 ( 
.A(n_1973),
.B(n_213),
.Y(n_2413)
);

NOR2xp67_ASAP7_75t_L g2414 ( 
.A(n_2024),
.B(n_580),
.Y(n_2414)
);

INVxp67_ASAP7_75t_L g2415 ( 
.A(n_1857),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_1782),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_1814),
.B(n_214),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1855),
.Y(n_2418)
);

BUFx4f_ASAP7_75t_L g2419 ( 
.A(n_2019),
.Y(n_2419)
);

AND2x6_ASAP7_75t_L g2420 ( 
.A(n_1845),
.B(n_214),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2012),
.B(n_215),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_1973),
.Y(n_2422)
);

BUFx8_ASAP7_75t_SL g2423 ( 
.A(n_2045),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_1943),
.B(n_1958),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2011),
.B(n_215),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_2029),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1855),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_1866),
.B(n_1870),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_1866),
.B(n_217),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_1845),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2000),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_1870),
.B(n_1895),
.Y(n_2432)
);

OR2x6_ASAP7_75t_L g2433 ( 
.A(n_1982),
.B(n_1983),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1959),
.Y(n_2434)
);

CKINVDCx20_ASAP7_75t_R g2435 ( 
.A(n_2025),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_2029),
.Y(n_2436)
);

NAND2x1p5_ASAP7_75t_L g2437 ( 
.A(n_1961),
.B(n_1852),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2005),
.B(n_217),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2000),
.Y(n_2439)
);

AND2x4_ASAP7_75t_L g2440 ( 
.A(n_1895),
.B(n_219),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1960),
.Y(n_2441)
);

INVx4_ASAP7_75t_L g2442 ( 
.A(n_1970),
.Y(n_2442)
);

INVx5_ASAP7_75t_L g2443 ( 
.A(n_2019),
.Y(n_2443)
);

INVxp67_ASAP7_75t_SL g2444 ( 
.A(n_1846),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2007),
.Y(n_2445)
);

INVx5_ASAP7_75t_L g2446 ( 
.A(n_2019),
.Y(n_2446)
);

CKINVDCx8_ASAP7_75t_R g2447 ( 
.A(n_1962),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_1971),
.B(n_219),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_SL g2449 ( 
.A(n_1846),
.B(n_582),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2006),
.B(n_220),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2011),
.B(n_220),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_1907),
.B(n_221),
.Y(n_2452)
);

NAND2x1_ASAP7_75t_L g2453 ( 
.A(n_1721),
.B(n_584),
.Y(n_2453)
);

NAND2x1p5_ASAP7_75t_L g2454 ( 
.A(n_1961),
.B(n_221),
.Y(n_2454)
);

OR2x6_ASAP7_75t_L g2455 ( 
.A(n_1982),
.B(n_222),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_1896),
.B(n_222),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_1896),
.B(n_223),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_1721),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_1857),
.B(n_1860),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_1983),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_1860),
.B(n_223),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_1907),
.B(n_224),
.Y(n_2462)
);

OR2x6_ASAP7_75t_L g2463 ( 
.A(n_1903),
.B(n_225),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_1903),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_1910),
.B(n_225),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_1757),
.Y(n_2466)
);

AND2x4_ASAP7_75t_L g2467 ( 
.A(n_1910),
.B(n_1991),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_1817),
.B(n_226),
.Y(n_2468)
);

INVx4_ASAP7_75t_L g2469 ( 
.A(n_1970),
.Y(n_2469)
);

OR2x6_ASAP7_75t_L g2470 ( 
.A(n_1987),
.B(n_227),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_1940),
.B(n_1800),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2007),
.Y(n_2472)
);

NAND2x1p5_ASAP7_75t_L g2473 ( 
.A(n_1961),
.B(n_1852),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_1728),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_1805),
.B(n_230),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2016),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_1991),
.B(n_231),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_2038),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2016),
.Y(n_2479)
);

NAND2x1p5_ASAP7_75t_L g2480 ( 
.A(n_1867),
.B(n_232),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_1819),
.Y(n_2481)
);

OR2x6_ASAP7_75t_L g2482 ( 
.A(n_1989),
.B(n_232),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_1954),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_1809),
.B(n_233),
.Y(n_2484)
);

OR2x6_ASAP7_75t_L g2485 ( 
.A(n_2052),
.B(n_233),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_1728),
.Y(n_2486)
);

NOR2x1_ASAP7_75t_L g2487 ( 
.A(n_1912),
.B(n_234),
.Y(n_2487)
);

INVx2_ASAP7_75t_SL g2488 ( 
.A(n_2053),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1963),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_1879),
.B(n_235),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_1760),
.B(n_235),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_1729),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_1867),
.B(n_236),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_2033),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_1911),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_1911),
.Y(n_2496)
);

OR2x2_ASAP7_75t_L g2497 ( 
.A(n_1715),
.B(n_236),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_1911),
.Y(n_2498)
);

BUFx4f_ASAP7_75t_L g2499 ( 
.A(n_1962),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1930),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1930),
.Y(n_2501)
);

INVxp67_ASAP7_75t_SL g2502 ( 
.A(n_1729),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_1741),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1936),
.B(n_237),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_1938),
.Y(n_2505)
);

INVx4_ASAP7_75t_L g2506 ( 
.A(n_1970),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2033),
.B(n_237),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_1970),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_1887),
.B(n_238),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_1962),
.Y(n_2510)
);

NAND2x1_ASAP7_75t_SL g2511 ( 
.A(n_2030),
.B(n_239),
.Y(n_2511)
);

BUFx2_ASAP7_75t_L g2512 ( 
.A(n_1962),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_1887),
.B(n_1967),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_1974),
.Y(n_2514)
);

INVx4_ASAP7_75t_L g2515 ( 
.A(n_1974),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_1735),
.B(n_239),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_1819),
.B(n_240),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_1819),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_1974),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_1743),
.B(n_241),
.Y(n_2520)
);

HB1xp67_ASAP7_75t_L g2521 ( 
.A(n_2151),
.Y(n_2521)
);

CKINVDCx16_ASAP7_75t_R g2522 ( 
.A(n_2069),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2252),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2129),
.Y(n_2524)
);

BUFx2_ASAP7_75t_L g2525 ( 
.A(n_2197),
.Y(n_2525)
);

INVx8_ASAP7_75t_L g2526 ( 
.A(n_2150),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2066),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2057),
.B(n_1962),
.Y(n_2528)
);

BUFx8_ASAP7_75t_L g2529 ( 
.A(n_2169),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_2125),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_2110),
.Y(n_2531)
);

BUFx2_ASAP7_75t_R g2532 ( 
.A(n_2250),
.Y(n_2532)
);

INVx1_ASAP7_75t_SL g2533 ( 
.A(n_2268),
.Y(n_2533)
);

INVx6_ASAP7_75t_SL g2534 ( 
.A(n_2070),
.Y(n_2534)
);

BUFx5_ASAP7_75t_L g2535 ( 
.A(n_2151),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2156),
.Y(n_2536)
);

BUFx6f_ASAP7_75t_L g2537 ( 
.A(n_2066),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2057),
.B(n_1962),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2229),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2424),
.Y(n_2540)
);

CKINVDCx14_ASAP7_75t_R g2541 ( 
.A(n_2104),
.Y(n_2541)
);

BUFx4_ASAP7_75t_SL g2542 ( 
.A(n_2070),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2176),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2088),
.Y(n_2544)
);

BUFx12f_ASAP7_75t_L g2545 ( 
.A(n_2188),
.Y(n_2545)
);

BUFx12f_ASAP7_75t_L g2546 ( 
.A(n_2152),
.Y(n_2546)
);

BUFx10_ASAP7_75t_L g2547 ( 
.A(n_2074),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2236),
.B(n_1861),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2110),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2386),
.B(n_1861),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2200),
.B(n_1880),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2156),
.Y(n_2552)
);

INVx3_ASAP7_75t_SL g2553 ( 
.A(n_2069),
.Y(n_2553)
);

INVx3_ASAP7_75t_SL g2554 ( 
.A(n_2096),
.Y(n_2554)
);

BUFx8_ASAP7_75t_SL g2555 ( 
.A(n_2211),
.Y(n_2555)
);

BUFx2_ASAP7_75t_L g2556 ( 
.A(n_2246),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2085),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2167),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2200),
.B(n_1892),
.Y(n_2559)
);

BUFx2_ASAP7_75t_SL g2560 ( 
.A(n_2074),
.Y(n_2560)
);

INVx5_ASAP7_75t_L g2561 ( 
.A(n_2073),
.Y(n_2561)
);

BUFx2_ASAP7_75t_SL g2562 ( 
.A(n_2083),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2298),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2099),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2067),
.B(n_1861),
.Y(n_2565)
);

BUFx12f_ASAP7_75t_L g2566 ( 
.A(n_2208),
.Y(n_2566)
);

CKINVDCx11_ASAP7_75t_R g2567 ( 
.A(n_2370),
.Y(n_2567)
);

BUFx2_ASAP7_75t_L g2568 ( 
.A(n_2210),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2167),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2183),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2447),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2210),
.Y(n_2572)
);

INVx4_ASAP7_75t_L g2573 ( 
.A(n_2210),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2066),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2099),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2061),
.Y(n_2576)
);

INVxp67_ASAP7_75t_SL g2577 ( 
.A(n_2444),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_2080),
.Y(n_2578)
);

BUFx6f_ASAP7_75t_L g2579 ( 
.A(n_2080),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2183),
.Y(n_2580)
);

INVx5_ASAP7_75t_L g2581 ( 
.A(n_2210),
.Y(n_2581)
);

CKINVDCx11_ASAP7_75t_R g2582 ( 
.A(n_2279),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2107),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2309),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2110),
.Y(n_2585)
);

BUFx3_ASAP7_75t_L g2586 ( 
.A(n_2190),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2201),
.Y(n_2587)
);

BUFx4_ASAP7_75t_SL g2588 ( 
.A(n_2073),
.Y(n_2588)
);

CKINVDCx14_ASAP7_75t_R g2589 ( 
.A(n_2208),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2061),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2107),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2149),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2201),
.B(n_2027),
.Y(n_2593)
);

INVx3_ASAP7_75t_SL g2594 ( 
.A(n_2279),
.Y(n_2594)
);

BUFx2_ASAP7_75t_SL g2595 ( 
.A(n_2083),
.Y(n_2595)
);

INVx3_ASAP7_75t_L g2596 ( 
.A(n_2149),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2059),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2260),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2277),
.B(n_1865),
.Y(n_2599)
);

INVx1_ASAP7_75t_SL g2600 ( 
.A(n_2260),
.Y(n_2600)
);

INVx2_ASAP7_75t_SL g2601 ( 
.A(n_2329),
.Y(n_2601)
);

BUFx3_ASAP7_75t_L g2602 ( 
.A(n_2213),
.Y(n_2602)
);

BUFx8_ASAP7_75t_L g2603 ( 
.A(n_2343),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_2260),
.Y(n_2604)
);

INVx3_ASAP7_75t_SL g2605 ( 
.A(n_2376),
.Y(n_2605)
);

INVx6_ASAP7_75t_L g2606 ( 
.A(n_2149),
.Y(n_2606)
);

BUFx4f_ASAP7_75t_L g2607 ( 
.A(n_2260),
.Y(n_2607)
);

BUFx2_ASAP7_75t_L g2608 ( 
.A(n_2372),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2113),
.Y(n_2609)
);

BUFx4f_ASAP7_75t_L g2610 ( 
.A(n_2257),
.Y(n_2610)
);

INVx2_ASAP7_75t_SL g2611 ( 
.A(n_2405),
.Y(n_2611)
);

NAND2x1p5_ASAP7_75t_L g2612 ( 
.A(n_2499),
.B(n_1741),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2113),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_2213),
.Y(n_2614)
);

INVx4_ASAP7_75t_L g2615 ( 
.A(n_2257),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2147),
.Y(n_2616)
);

INVx5_ASAP7_75t_L g2617 ( 
.A(n_2134),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_2121),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2064),
.B(n_2018),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2392),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2059),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2063),
.Y(n_2622)
);

BUFx12f_ASAP7_75t_L g2623 ( 
.A(n_2112),
.Y(n_2623)
);

INVx5_ASAP7_75t_SL g2624 ( 
.A(n_2098),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2499),
.Y(n_2625)
);

BUFx2_ASAP7_75t_R g2626 ( 
.A(n_2262),
.Y(n_2626)
);

INVx1_ASAP7_75t_SL g2627 ( 
.A(n_2297),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2123),
.Y(n_2628)
);

INVx4_ASAP7_75t_L g2629 ( 
.A(n_2258),
.Y(n_2629)
);

BUFx12f_ASAP7_75t_L g2630 ( 
.A(n_2195),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2072),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2064),
.B(n_2018),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_L g2633 ( 
.A(n_2080),
.Y(n_2633)
);

BUFx6f_ASAP7_75t_SL g2634 ( 
.A(n_2124),
.Y(n_2634)
);

INVxp67_ASAP7_75t_SL g2635 ( 
.A(n_2297),
.Y(n_2635)
);

INVx4_ASAP7_75t_L g2636 ( 
.A(n_2258),
.Y(n_2636)
);

BUFx4_ASAP7_75t_SL g2637 ( 
.A(n_2098),
.Y(n_2637)
);

INVx4_ASAP7_75t_L g2638 ( 
.A(n_2134),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2408),
.B(n_1865),
.Y(n_2639)
);

BUFx3_ASAP7_75t_L g2640 ( 
.A(n_2056),
.Y(n_2640)
);

BUFx2_ASAP7_75t_L g2641 ( 
.A(n_2134),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2123),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2159),
.Y(n_2643)
);

BUFx3_ASAP7_75t_L g2644 ( 
.A(n_2056),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2135),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2275),
.B(n_2161),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2159),
.Y(n_2647)
);

INVx3_ASAP7_75t_L g2648 ( 
.A(n_2357),
.Y(n_2648)
);

NAND2x1p5_ASAP7_75t_L g2649 ( 
.A(n_2302),
.B(n_1974),
.Y(n_2649)
);

NAND2x1p5_ASAP7_75t_L g2650 ( 
.A(n_2302),
.B(n_1930),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2135),
.Y(n_2651)
);

INVx3_ASAP7_75t_SL g2652 ( 
.A(n_2124),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2161),
.A2(n_2001),
.B1(n_2010),
.B2(n_1997),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2285),
.A2(n_1908),
.B1(n_1915),
.B2(n_1893),
.Y(n_2654)
);

BUFx3_ASAP7_75t_L g2655 ( 
.A(n_2195),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2114),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_2357),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2285),
.B(n_1865),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2063),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2202),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2119),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2202),
.Y(n_2662)
);

INVx8_ASAP7_75t_L g2663 ( 
.A(n_2134),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2120),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2267),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2180),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2267),
.Y(n_2667)
);

INVx2_ASAP7_75t_SL g2668 ( 
.A(n_2127),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2299),
.B(n_1747),
.Y(n_2669)
);

INVx2_ASAP7_75t_SL g2670 ( 
.A(n_2251),
.Y(n_2670)
);

NAND2x1p5_ASAP7_75t_L g2671 ( 
.A(n_2243),
.B(n_2031),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2434),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2434),
.Y(n_2673)
);

BUFx5_ASAP7_75t_L g2674 ( 
.A(n_2214),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2214),
.Y(n_2675)
);

INVx5_ASAP7_75t_L g2676 ( 
.A(n_2364),
.Y(n_2676)
);

NAND2x1p5_ASAP7_75t_L g2677 ( 
.A(n_2243),
.B(n_2251),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2418),
.B(n_1776),
.Y(n_2678)
);

BUFx12f_ASAP7_75t_L g2679 ( 
.A(n_2180),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2299),
.A2(n_1776),
.B1(n_2035),
.B2(n_2037),
.Y(n_2680)
);

INVx4_ASAP7_75t_L g2681 ( 
.A(n_2364),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_2136),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2304),
.A2(n_2030),
.B1(n_1850),
.B2(n_1996),
.Y(n_2683)
);

BUFx6f_ASAP7_75t_L g2684 ( 
.A(n_2081),
.Y(n_2684)
);

CKINVDCx16_ASAP7_75t_R g2685 ( 
.A(n_2300),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2217),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2418),
.B(n_1996),
.Y(n_2687)
);

BUFx5_ASAP7_75t_L g2688 ( 
.A(n_2217),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2304),
.B(n_1754),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_2313),
.Y(n_2690)
);

BUFx3_ASAP7_75t_L g2691 ( 
.A(n_2116),
.Y(n_2691)
);

BUFx2_ASAP7_75t_SL g2692 ( 
.A(n_2276),
.Y(n_2692)
);

BUFx3_ASAP7_75t_L g2693 ( 
.A(n_2158),
.Y(n_2693)
);

BUFx3_ASAP7_75t_L g2694 ( 
.A(n_2292),
.Y(n_2694)
);

INVx1_ASAP7_75t_SL g2695 ( 
.A(n_2493),
.Y(n_2695)
);

CKINVDCx20_ASAP7_75t_R g2696 ( 
.A(n_2423),
.Y(n_2696)
);

INVx1_ASAP7_75t_SL g2697 ( 
.A(n_2493),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2097),
.Y(n_2698)
);

BUFx12f_ASAP7_75t_L g2699 ( 
.A(n_2316),
.Y(n_2699)
);

INVx1_ASAP7_75t_SL g2700 ( 
.A(n_2175),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2441),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_L g2702 ( 
.A1(n_2318),
.A2(n_2030),
.B1(n_1850),
.B2(n_1897),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2441),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_2318),
.A2(n_1786),
.B1(n_1829),
.B2(n_1745),
.Y(n_2704)
);

BUFx3_ASAP7_75t_L g2705 ( 
.A(n_2287),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2448),
.Y(n_2706)
);

BUFx6f_ASAP7_75t_L g2707 ( 
.A(n_2081),
.Y(n_2707)
);

CKINVDCx11_ASAP7_75t_R g2708 ( 
.A(n_2413),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2212),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2218),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2427),
.B(n_1829),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2427),
.B(n_1771),
.Y(n_2712)
);

BUFx2_ASAP7_75t_SL g2713 ( 
.A(n_2115),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2212),
.Y(n_2714)
);

NAND2x1p5_ASAP7_75t_L g2715 ( 
.A(n_2172),
.B(n_2510),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2225),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2218),
.Y(n_2717)
);

CKINVDCx16_ASAP7_75t_R g2718 ( 
.A(n_2463),
.Y(n_2718)
);

INVx5_ASAP7_75t_L g2719 ( 
.A(n_2364),
.Y(n_2719)
);

INVxp67_ASAP7_75t_SL g2720 ( 
.A(n_2419),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2459),
.B(n_1812),
.Y(n_2721)
);

INVx5_ASAP7_75t_SL g2722 ( 
.A(n_2230),
.Y(n_2722)
);

BUFx3_ASAP7_75t_L g2723 ( 
.A(n_2287),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_SL g2724 ( 
.A(n_2115),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2221),
.Y(n_2725)
);

BUFx2_ASAP7_75t_L g2726 ( 
.A(n_2364),
.Y(n_2726)
);

INVx1_ASAP7_75t_SL g2727 ( 
.A(n_2175),
.Y(n_2727)
);

BUFx24_ASAP7_75t_L g2728 ( 
.A(n_2205),
.Y(n_2728)
);

INVx4_ASAP7_75t_L g2729 ( 
.A(n_2172),
.Y(n_2729)
);

OR2x6_ASAP7_75t_L g2730 ( 
.A(n_2463),
.B(n_2031),
.Y(n_2730)
);

INVx1_ASAP7_75t_SL g2731 ( 
.A(n_2380),
.Y(n_2731)
);

INVx5_ASAP7_75t_L g2732 ( 
.A(n_2081),
.Y(n_2732)
);

INVx5_ASAP7_75t_L g2733 ( 
.A(n_2095),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_L g2734 ( 
.A(n_2265),
.B(n_1816),
.Y(n_2734)
);

NAND2x1p5_ASAP7_75t_L g2735 ( 
.A(n_2512),
.B(n_2031),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2269),
.Y(n_2736)
);

CKINVDCx20_ASAP7_75t_R g2737 ( 
.A(n_2286),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2225),
.Y(n_2738)
);

INVxp67_ASAP7_75t_SL g2739 ( 
.A(n_2419),
.Y(n_2739)
);

NAND2x1p5_ASAP7_75t_L g2740 ( 
.A(n_2164),
.B(n_2031),
.Y(n_2740)
);

CKINVDCx20_ASAP7_75t_R g2741 ( 
.A(n_2366),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2221),
.B(n_1824),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2248),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2248),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2387),
.Y(n_2745)
);

INVx5_ASAP7_75t_L g2746 ( 
.A(n_2095),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2223),
.B(n_1834),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2223),
.B(n_1842),
.Y(n_2748)
);

BUFx12f_ASAP7_75t_L g2749 ( 
.A(n_2320),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2105),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2089),
.Y(n_2751)
);

BUFx3_ASAP7_75t_L g2752 ( 
.A(n_2105),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2143),
.B(n_1790),
.Y(n_2753)
);

BUFx12f_ASAP7_75t_L g2754 ( 
.A(n_2294),
.Y(n_2754)
);

CKINVDCx20_ASAP7_75t_R g2755 ( 
.A(n_2092),
.Y(n_2755)
);

INVx2_ASAP7_75t_SL g2756 ( 
.A(n_2205),
.Y(n_2756)
);

NAND2x1p5_ASAP7_75t_L g2757 ( 
.A(n_2164),
.B(n_1790),
.Y(n_2757)
);

NAND2x1p5_ASAP7_75t_L g2758 ( 
.A(n_2173),
.B(n_1790),
.Y(n_2758)
);

BUFx12f_ASAP7_75t_L g2759 ( 
.A(n_2118),
.Y(n_2759)
);

BUFx3_ASAP7_75t_L g2760 ( 
.A(n_2090),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2379),
.Y(n_2761)
);

NAND2x1p5_ASAP7_75t_L g2762 ( 
.A(n_2173),
.B(n_1791),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2233),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2460),
.B(n_1849),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2233),
.Y(n_2765)
);

BUFx12f_ASAP7_75t_L g2766 ( 
.A(n_2193),
.Y(n_2766)
);

NAND2x1p5_ASAP7_75t_L g2767 ( 
.A(n_2179),
.B(n_1791),
.Y(n_2767)
);

OR2x6_ASAP7_75t_L g2768 ( 
.A(n_2179),
.B(n_2185),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2241),
.B(n_2483),
.Y(n_2769)
);

INVx3_ASAP7_75t_SL g2770 ( 
.A(n_2171),
.Y(n_2770)
);

BUFx4f_ASAP7_75t_SL g2771 ( 
.A(n_2143),
.Y(n_2771)
);

BUFx3_ASAP7_75t_L g2772 ( 
.A(n_2356),
.Y(n_2772)
);

INVx1_ASAP7_75t_SL g2773 ( 
.A(n_2380),
.Y(n_2773)
);

INVx4_ASAP7_75t_L g2774 ( 
.A(n_2420),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_2241),
.Y(n_2775)
);

BUFx3_ASAP7_75t_L g2776 ( 
.A(n_2381),
.Y(n_2776)
);

BUFx2_ASAP7_75t_SL g2777 ( 
.A(n_2253),
.Y(n_2777)
);

INVx5_ASAP7_75t_L g2778 ( 
.A(n_2095),
.Y(n_2778)
);

BUFx12f_ASAP7_75t_L g2779 ( 
.A(n_2291),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2192),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2483),
.B(n_1851),
.Y(n_2781)
);

BUFx12f_ASAP7_75t_L g2782 ( 
.A(n_2327),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2103),
.Y(n_2783)
);

INVx1_ASAP7_75t_SL g2784 ( 
.A(n_2517),
.Y(n_2784)
);

BUFx2_ASAP7_75t_SL g2785 ( 
.A(n_2253),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2399),
.B(n_1791),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_2371),
.Y(n_2787)
);

INVx5_ASAP7_75t_L g2788 ( 
.A(n_2293),
.Y(n_2788)
);

INVx2_ASAP7_75t_SL g2789 ( 
.A(n_2259),
.Y(n_2789)
);

BUFx3_ASAP7_75t_L g2790 ( 
.A(n_2259),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2155),
.B(n_1797),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2141),
.B(n_1858),
.Y(n_2792)
);

BUFx2_ASAP7_75t_L g2793 ( 
.A(n_2185),
.Y(n_2793)
);

CKINVDCx5p33_ASAP7_75t_R g2794 ( 
.A(n_2464),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2371),
.Y(n_2795)
);

NAND2x1p5_ASAP7_75t_L g2796 ( 
.A(n_2442),
.B(n_1992),
.Y(n_2796)
);

INVx3_ASAP7_75t_L g2797 ( 
.A(n_2442),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2271),
.Y(n_2798)
);

INVx2_ASAP7_75t_SL g2799 ( 
.A(n_2271),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2103),
.Y(n_2800)
);

BUFx2_ASAP7_75t_L g2801 ( 
.A(n_2420),
.Y(n_2801)
);

INVx6_ASAP7_75t_L g2802 ( 
.A(n_2413),
.Y(n_2802)
);

BUFx2_ASAP7_75t_SL g2803 ( 
.A(n_2334),
.Y(n_2803)
);

BUFx3_ASAP7_75t_L g2804 ( 
.A(n_2137),
.Y(n_2804)
);

CKINVDCx8_ASAP7_75t_R g2805 ( 
.A(n_2420),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2137),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2142),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2334),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2142),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2489),
.B(n_1745),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2360),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2360),
.Y(n_2812)
);

INVx6_ASAP7_75t_SL g2813 ( 
.A(n_2389),
.Y(n_2813)
);

BUFx3_ASAP7_75t_L g2814 ( 
.A(n_2261),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2389),
.Y(n_2815)
);

BUFx2_ASAP7_75t_L g2816 ( 
.A(n_2420),
.Y(n_2816)
);

NAND2x1_ASAP7_75t_L g2817 ( 
.A(n_2469),
.B(n_1992),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2261),
.Y(n_2818)
);

CKINVDCx5p33_ASAP7_75t_R g2819 ( 
.A(n_2455),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2062),
.Y(n_2820)
);

INVx3_ASAP7_75t_L g2821 ( 
.A(n_2469),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2103),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2404),
.B(n_241),
.Y(n_2823)
);

INVx8_ASAP7_75t_L g2824 ( 
.A(n_2455),
.Y(n_2824)
);

CKINVDCx6p67_ASAP7_75t_R g2825 ( 
.A(n_2470),
.Y(n_2825)
);

INVx4_ASAP7_75t_L g2826 ( 
.A(n_2506),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2435),
.A2(n_1980),
.B1(n_2004),
.B2(n_2041),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2282),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_2282),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2399),
.B(n_2048),
.Y(n_2830)
);

BUFx10_ASAP7_75t_L g2831 ( 
.A(n_2198),
.Y(n_2831)
);

BUFx3_ASAP7_75t_L g2832 ( 
.A(n_2306),
.Y(n_2832)
);

INVx1_ASAP7_75t_SL g2833 ( 
.A(n_2517),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_2470),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2306),
.Y(n_2835)
);

BUFx4_ASAP7_75t_SL g2836 ( 
.A(n_2482),
.Y(n_2836)
);

INVxp67_ASAP7_75t_SL g2837 ( 
.A(n_2361),
.Y(n_2837)
);

BUFx3_ASAP7_75t_L g2838 ( 
.A(n_2308),
.Y(n_2838)
);

INVx1_ASAP7_75t_SL g2839 ( 
.A(n_2308),
.Y(n_2839)
);

BUFx8_ASAP7_75t_L g2840 ( 
.A(n_2249),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2068),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2315),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2237),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2315),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2242),
.Y(n_2845)
);

BUFx4f_ASAP7_75t_SL g2846 ( 
.A(n_2506),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2323),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2489),
.B(n_1950),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2157),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2407),
.B(n_242),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_2102),
.Y(n_2851)
);

BUFx10_ASAP7_75t_L g2852 ( 
.A(n_2198),
.Y(n_2852)
);

NAND2x1p5_ASAP7_75t_L g2853 ( 
.A(n_2515),
.B(n_1993),
.Y(n_2853)
);

BUFx6f_ASAP7_75t_SL g2854 ( 
.A(n_2204),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2428),
.B(n_1950),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2323),
.Y(n_2856)
);

BUFx12f_ASAP7_75t_L g2857 ( 
.A(n_2480),
.Y(n_2857)
);

BUFx4_ASAP7_75t_SL g2858 ( 
.A(n_2482),
.Y(n_2858)
);

INVx3_ASAP7_75t_L g2859 ( 
.A(n_2515),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_2331),
.Y(n_2860)
);

BUFx12f_ASAP7_75t_L g2861 ( 
.A(n_2178),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2245),
.Y(n_2862)
);

BUFx4f_ASAP7_75t_SL g2863 ( 
.A(n_2117),
.Y(n_2863)
);

OR2x6_ASAP7_75t_L g2864 ( 
.A(n_2454),
.B(n_2048),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_2331),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2204),
.Y(n_2866)
);

INVxp33_ASAP7_75t_SL g2867 ( 
.A(n_2505),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_2332),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2303),
.B(n_1993),
.Y(n_2869)
);

INVx1_ASAP7_75t_SL g2870 ( 
.A(n_2332),
.Y(n_2870)
);

AND2x4_ASAP7_75t_L g2871 ( 
.A(n_2234),
.B(n_2041),
.Y(n_2871)
);

AOI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_2347),
.A2(n_1950),
.B1(n_245),
.B2(n_243),
.Y(n_2872)
);

BUFx12f_ASAP7_75t_L g2873 ( 
.A(n_2396),
.Y(n_2873)
);

CKINVDCx5p33_ASAP7_75t_R g2874 ( 
.A(n_2485),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2335),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2077),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2122),
.Y(n_2877)
);

BUFx6f_ASAP7_75t_L g2878 ( 
.A(n_2157),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2335),
.Y(n_2879)
);

OAI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2494),
.A2(n_2430),
.B1(n_2415),
.B2(n_2429),
.Y(n_2880)
);

CKINVDCx5p33_ASAP7_75t_R g2881 ( 
.A(n_2485),
.Y(n_2881)
);

BUFx6f_ASAP7_75t_L g2882 ( 
.A(n_2157),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2130),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2346),
.Y(n_2884)
);

INVx8_ASAP7_75t_L g2885 ( 
.A(n_2417),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_SL g2886 ( 
.A(n_2417),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2346),
.Y(n_2887)
);

INVx2_ASAP7_75t_SL g2888 ( 
.A(n_2079),
.Y(n_2888)
);

INVxp67_ASAP7_75t_SL g2889 ( 
.A(n_2361),
.Y(n_2889)
);

INVx2_ASAP7_75t_SL g2890 ( 
.A(n_2429),
.Y(n_2890)
);

INVxp67_ASAP7_75t_SL g2891 ( 
.A(n_2472),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2472),
.Y(n_2892)
);

OR2x6_ASAP7_75t_L g2893 ( 
.A(n_2305),
.B(n_1950),
.Y(n_2893)
);

INVx1_ASAP7_75t_SL g2894 ( 
.A(n_2476),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2428),
.B(n_1950),
.Y(n_2895)
);

BUFx12f_ASAP7_75t_L g2896 ( 
.A(n_2239),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2131),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2231),
.Y(n_2898)
);

BUFx6f_ASAP7_75t_L g2899 ( 
.A(n_2182),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2620),
.B(n_2076),
.Y(n_2900)
);

INVx4_ASAP7_75t_L g2901 ( 
.A(n_2526),
.Y(n_2901)
);

CKINVDCx6p67_ASAP7_75t_R g2902 ( 
.A(n_2545),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_SL g2903 ( 
.A1(n_2718),
.A2(n_2186),
.B1(n_2254),
.B2(n_2478),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2891),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2722),
.A2(n_2256),
.B1(n_2307),
.B2(n_2278),
.Y(n_2905)
);

CKINVDCx6p67_ASAP7_75t_R g2906 ( 
.A(n_2630),
.Y(n_2906)
);

AOI22xp33_ASAP7_75t_L g2907 ( 
.A1(n_2722),
.A2(n_2278),
.B1(n_2433),
.B2(n_2406),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2891),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2839),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_L g2910 ( 
.A1(n_2722),
.A2(n_2433),
.B1(n_2395),
.B2(n_2432),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_SL g2911 ( 
.A1(n_2589),
.A2(n_2629),
.B1(n_2636),
.B2(n_2615),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2775),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2775),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2610),
.A2(n_2432),
.B1(n_2467),
.B2(n_2166),
.Y(n_2914)
);

CKINVDCx20_ASAP7_75t_R g2915 ( 
.A(n_2603),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2523),
.B(n_2467),
.Y(n_2916)
);

BUFx2_ASAP7_75t_L g2917 ( 
.A(n_2768),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2540),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2768),
.Y(n_2919)
);

OAI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2734),
.A2(n_2471),
.B(n_2283),
.Y(n_2920)
);

BUFx6f_ASAP7_75t_L g2921 ( 
.A(n_2606),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2734),
.B(n_2317),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2656),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2661),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2664),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2839),
.Y(n_2926)
);

AOI22xp33_ASAP7_75t_SL g2927 ( 
.A1(n_2560),
.A2(n_2449),
.B1(n_2401),
.B2(n_2394),
.Y(n_2927)
);

INVx2_ASAP7_75t_SL g2928 ( 
.A(n_2603),
.Y(n_2928)
);

AOI22xp33_ASAP7_75t_L g2929 ( 
.A1(n_2610),
.A2(n_2456),
.B1(n_2457),
.B2(n_2440),
.Y(n_2929)
);

AOI22xp33_ASAP7_75t_SL g2930 ( 
.A1(n_2562),
.A2(n_2595),
.B1(n_2624),
.B2(n_2824),
.Y(n_2930)
);

AOI22xp33_ASAP7_75t_SL g2931 ( 
.A1(n_2624),
.A2(n_2449),
.B1(n_2401),
.B2(n_2394),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2768),
.B(n_2082),
.Y(n_2932)
);

CKINVDCx11_ASAP7_75t_R g2933 ( 
.A(n_2526),
.Y(n_2933)
);

OAI22xp33_ASAP7_75t_L g2934 ( 
.A1(n_2885),
.A2(n_2412),
.B1(n_2410),
.B2(n_2324),
.Y(n_2934)
);

INVx5_ASAP7_75t_L g2935 ( 
.A(n_2526),
.Y(n_2935)
);

BUFx12f_ASAP7_75t_L g2936 ( 
.A(n_2529),
.Y(n_2936)
);

INVx4_ASAP7_75t_L g2937 ( 
.A(n_2663),
.Y(n_2937)
);

CKINVDCx20_ASAP7_75t_R g2938 ( 
.A(n_2529),
.Y(n_2938)
);

AOI22xp33_ASAP7_75t_L g2939 ( 
.A1(n_2634),
.A2(n_2456),
.B1(n_2457),
.B2(n_2440),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2805),
.A2(n_2465),
.B1(n_2477),
.B2(n_2461),
.Y(n_2940)
);

OAI21xp5_ASAP7_75t_SL g2941 ( 
.A1(n_2677),
.A2(n_2244),
.B(n_2465),
.Y(n_2941)
);

INVx4_ASAP7_75t_L g2942 ( 
.A(n_2663),
.Y(n_2942)
);

AOI22xp33_ASAP7_75t_L g2943 ( 
.A1(n_2634),
.A2(n_2477),
.B1(n_2375),
.B2(n_2390),
.Y(n_2943)
);

CKINVDCx20_ASAP7_75t_R g2944 ( 
.A(n_2696),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2708),
.A2(n_2325),
.B1(n_2400),
.B2(n_2398),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2870),
.Y(n_2946)
);

BUFx2_ASAP7_75t_R g2947 ( 
.A(n_2544),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2870),
.Y(n_2948)
);

BUFx6f_ASAP7_75t_L g2949 ( 
.A(n_2606),
.Y(n_2949)
);

INVx4_ASAP7_75t_L g2950 ( 
.A(n_2663),
.Y(n_2950)
);

INVx1_ASAP7_75t_SL g2951 ( 
.A(n_2608),
.Y(n_2951)
);

BUFx2_ASAP7_75t_L g2952 ( 
.A(n_2534),
.Y(n_2952)
);

NAND2x1p5_ASAP7_75t_L g2953 ( 
.A(n_2524),
.B(n_2293),
.Y(n_2953)
);

AOI22xp33_ASAP7_75t_SL g2954 ( 
.A1(n_2624),
.A2(n_2324),
.B1(n_2333),
.B2(n_2322),
.Y(n_2954)
);

HB1xp67_ASAP7_75t_L g2955 ( 
.A(n_2631),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2564),
.Y(n_2956)
);

OAI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2677),
.A2(n_2328),
.B1(n_2093),
.B2(n_2342),
.Y(n_2957)
);

OAI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2885),
.A2(n_2333),
.B1(n_2322),
.B2(n_2100),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2894),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_SL g2960 ( 
.A1(n_2824),
.A2(n_2100),
.B1(n_2109),
.B2(n_2065),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2828),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2828),
.Y(n_2962)
);

CKINVDCx20_ASAP7_75t_R g2963 ( 
.A(n_2554),
.Y(n_2963)
);

BUFx10_ASAP7_75t_L g2964 ( 
.A(n_2530),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2527),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_SL g2966 ( 
.A1(n_2824),
.A2(n_2109),
.B1(n_2128),
.B2(n_2065),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_SL g2967 ( 
.A1(n_2713),
.A2(n_2177),
.B1(n_2203),
.B2(n_2128),
.Y(n_2967)
);

BUFx12f_ASAP7_75t_L g2968 ( 
.A(n_2582),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2575),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2583),
.Y(n_2970)
);

INVx8_ASAP7_75t_L g2971 ( 
.A(n_2546),
.Y(n_2971)
);

AOI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2886),
.A2(n_2422),
.B1(n_2087),
.B2(n_2187),
.Y(n_2972)
);

BUFx8_ASAP7_75t_L g2973 ( 
.A(n_2566),
.Y(n_2973)
);

OAI21xp33_ASAP7_75t_L g2974 ( 
.A1(n_2654),
.A2(n_2312),
.B(n_2290),
.Y(n_2974)
);

AOI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2837),
.A2(n_2889),
.B(n_2383),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_SL g2976 ( 
.A1(n_2777),
.A2(n_2203),
.B1(n_2177),
.B2(n_2468),
.Y(n_2976)
);

CKINVDCx20_ASAP7_75t_R g2977 ( 
.A(n_2541),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2792),
.B(n_2181),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2591),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2527),
.Y(n_2980)
);

CKINVDCx6p67_ASAP7_75t_R g2981 ( 
.A(n_2728),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2894),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2609),
.Y(n_2983)
);

OAI21xp5_ASAP7_75t_SL g2984 ( 
.A1(n_2801),
.A2(n_2490),
.B(n_2274),
.Y(n_2984)
);

AOI22xp5_ASAP7_75t_L g2985 ( 
.A1(n_2886),
.A2(n_2206),
.B1(n_2220),
.B2(n_2191),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2601),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2536),
.Y(n_2987)
);

OAI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2885),
.A2(n_2272),
.B1(n_2263),
.B2(n_2310),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2552),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2587),
.B(n_2227),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2558),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2521),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_2741),
.Y(n_2993)
);

INVx11_ASAP7_75t_L g2994 ( 
.A(n_2857),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2615),
.A2(n_2138),
.B1(n_2133),
.B2(n_2280),
.Y(n_2995)
);

AOI22xp33_ASAP7_75t_L g2996 ( 
.A1(n_2629),
.A2(n_2209),
.B1(n_2199),
.B2(n_2520),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_2836),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2613),
.Y(n_2998)
);

BUFx12f_ASAP7_75t_L g2999 ( 
.A(n_2567),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2569),
.Y(n_3000)
);

AOI22xp33_ASAP7_75t_L g3001 ( 
.A1(n_2636),
.A2(n_2349),
.B1(n_2337),
.B2(n_2339),
.Y(n_3001)
);

INVx6_ASAP7_75t_L g3002 ( 
.A(n_2685),
.Y(n_3002)
);

INVx6_ASAP7_75t_L g3003 ( 
.A(n_2896),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2635),
.A2(n_2108),
.B1(n_2319),
.B2(n_2314),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2854),
.A2(n_2338),
.B1(n_2311),
.B2(n_2345),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2854),
.A2(n_2397),
.B1(n_2402),
.B2(n_2391),
.Y(n_3006)
);

INVx1_ASAP7_75t_SL g3007 ( 
.A(n_2836),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2550),
.B(n_2646),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2690),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2823),
.B(n_2086),
.Y(n_3010)
);

INVx6_ASAP7_75t_L g3011 ( 
.A(n_2547),
.Y(n_3011)
);

AOI22xp33_ASAP7_75t_L g3012 ( 
.A1(n_2802),
.A2(n_2326),
.B1(n_2378),
.B2(n_2330),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2867),
.A2(n_2450),
.B1(n_2438),
.B2(n_2224),
.Y(n_3013)
);

CKINVDCx11_ASAP7_75t_R g3014 ( 
.A(n_2605),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2521),
.Y(n_3015)
);

AOI22xp33_ASAP7_75t_L g3016 ( 
.A1(n_2802),
.A2(n_2679),
.B1(n_2724),
.B2(n_2681),
.Y(n_3016)
);

INVx1_ASAP7_75t_SL g3017 ( 
.A(n_2858),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2597),
.Y(n_3018)
);

BUFx6f_ASAP7_75t_L g3019 ( 
.A(n_2527),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2621),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2570),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2724),
.A2(n_2084),
.B1(n_2234),
.B2(n_2058),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2622),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_2681),
.A2(n_2060),
.B1(n_2228),
.B2(n_2139),
.Y(n_3024)
);

BUFx6f_ASAP7_75t_L g3025 ( 
.A(n_2537),
.Y(n_3025)
);

CKINVDCx11_ASAP7_75t_R g3026 ( 
.A(n_2553),
.Y(n_3026)
);

BUFx2_ASAP7_75t_SL g3027 ( 
.A(n_2611),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_SL g3028 ( 
.A1(n_2785),
.A2(n_2353),
.B1(n_2446),
.B2(n_2443),
.Y(n_3028)
);

INVx1_ASAP7_75t_SL g3029 ( 
.A(n_2858),
.Y(n_3029)
);

BUFx2_ASAP7_75t_L g3030 ( 
.A(n_2534),
.Y(n_3030)
);

BUFx10_ASAP7_75t_L g3031 ( 
.A(n_2730),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2850),
.B(n_2270),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2580),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2774),
.A2(n_2132),
.B1(n_2484),
.B2(n_2475),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2628),
.Y(n_3035)
);

INVx5_ASAP7_75t_L g3036 ( 
.A(n_2730),
.Y(n_3036)
);

BUFx10_ASAP7_75t_L g3037 ( 
.A(n_2730),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2642),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2543),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2659),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2645),
.Y(n_3041)
);

INVx6_ASAP7_75t_L g3042 ( 
.A(n_2547),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_L g3043 ( 
.A1(n_2774),
.A2(n_2466),
.B1(n_2189),
.B2(n_2362),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2706),
.B(n_2403),
.Y(n_3044)
);

BUFx4f_ASAP7_75t_SL g3045 ( 
.A(n_2655),
.Y(n_3045)
);

HB1xp67_ASAP7_75t_L g3046 ( 
.A(n_2637),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2651),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2672),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2803),
.B(n_2235),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2563),
.Y(n_3050)
);

NAND2x1p5_ASAP7_75t_L g3051 ( 
.A(n_2561),
.B(n_2443),
.Y(n_3051)
);

CKINVDCx5p33_ASAP7_75t_R g3052 ( 
.A(n_2532),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2673),
.Y(n_3053)
);

CKINVDCx20_ASAP7_75t_R g3054 ( 
.A(n_2555),
.Y(n_3054)
);

OAI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2825),
.A2(n_2491),
.B1(n_2353),
.B2(n_2497),
.Y(n_3055)
);

OAI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_2652),
.A2(n_2446),
.B1(n_2443),
.B2(n_2101),
.Y(n_3056)
);

OAI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_2635),
.A2(n_2369),
.B1(n_2373),
.B2(n_2358),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2701),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2703),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2769),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2769),
.Y(n_3061)
);

BUFx6f_ASAP7_75t_L g3062 ( 
.A(n_2537),
.Y(n_3062)
);

INVx3_ASAP7_75t_L g3063 ( 
.A(n_2863),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2660),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_SL g3065 ( 
.A1(n_2638),
.A2(n_2446),
.B1(n_2196),
.B2(n_2488),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2662),
.Y(n_3066)
);

BUFx12f_ASAP7_75t_L g3067 ( 
.A(n_2682),
.Y(n_3067)
);

OAI22xp5_ASAP7_75t_SL g3068 ( 
.A1(n_2819),
.A2(n_2163),
.B1(n_2421),
.B2(n_2301),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2880),
.A2(n_2638),
.B1(n_2666),
.B2(n_2754),
.Y(n_3069)
);

BUFx2_ASAP7_75t_L g3070 ( 
.A(n_2813),
.Y(n_3070)
);

INVxp67_ASAP7_75t_SL g3071 ( 
.A(n_2757),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2880),
.A2(n_2782),
.B1(n_2791),
.B2(n_2561),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2675),
.Y(n_3073)
);

OAI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2607),
.A2(n_2451),
.B1(n_2425),
.B2(n_2507),
.Y(n_3074)
);

CKINVDCx11_ASAP7_75t_R g3075 ( 
.A(n_2594),
.Y(n_3075)
);

INVx1_ASAP7_75t_SL g3076 ( 
.A(n_2586),
.Y(n_3076)
);

INVx3_ASAP7_75t_L g3077 ( 
.A(n_2863),
.Y(n_3077)
);

INVx3_ASAP7_75t_L g3078 ( 
.A(n_2573),
.Y(n_3078)
);

CKINVDCx6p67_ASAP7_75t_R g3079 ( 
.A(n_2561),
.Y(n_3079)
);

OAI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2607),
.A2(n_2170),
.B1(n_2165),
.B2(n_2216),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2686),
.Y(n_3081)
);

INVxp67_ASAP7_75t_SL g3082 ( 
.A(n_2757),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2898),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2710),
.Y(n_3084)
);

OAI21xp5_ASAP7_75t_SL g3085 ( 
.A1(n_2816),
.A2(n_2487),
.B(n_2341),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_SL g3086 ( 
.A1(n_2793),
.A2(n_2196),
.B1(n_2174),
.B2(n_2476),
.Y(n_3086)
);

BUFx8_ASAP7_75t_L g3087 ( 
.A(n_2525),
.Y(n_3087)
);

BUFx6f_ASAP7_75t_L g3088 ( 
.A(n_2537),
.Y(n_3088)
);

OAI22xp33_ASAP7_75t_L g3089 ( 
.A1(n_2834),
.A2(n_2091),
.B1(n_2222),
.B2(n_2411),
.Y(n_3089)
);

NAND2x1p5_ASAP7_75t_L g3090 ( 
.A(n_2581),
.B(n_2232),
.Y(n_3090)
);

INVx6_ASAP7_75t_L g3091 ( 
.A(n_2729),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_2873),
.A2(n_2350),
.B1(n_2516),
.B2(n_2504),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2868),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2717),
.Y(n_3094)
);

CKINVDCx8_ASAP7_75t_R g3095 ( 
.A(n_2692),
.Y(n_3095)
);

OAI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_2874),
.A2(n_2881),
.B1(n_2813),
.B2(n_2762),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2755),
.A2(n_2071),
.B1(n_2075),
.B2(n_2162),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2725),
.Y(n_3098)
);

AOI22xp33_ASAP7_75t_L g3099 ( 
.A1(n_2726),
.A2(n_2462),
.B1(n_2452),
.B2(n_2148),
.Y(n_3099)
);

OAI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2758),
.A2(n_2513),
.B1(n_2479),
.B2(n_2509),
.Y(n_3100)
);

BUFx3_ASAP7_75t_L g3101 ( 
.A(n_2584),
.Y(n_3101)
);

BUFx10_ASAP7_75t_L g3102 ( 
.A(n_2794),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2763),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2758),
.A2(n_2479),
.B1(n_2359),
.B2(n_2374),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2765),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2806),
.Y(n_3106)
);

BUFx4f_ASAP7_75t_SL g3107 ( 
.A(n_2861),
.Y(n_3107)
);

INVx3_ASAP7_75t_L g3108 ( 
.A(n_2573),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2699),
.A2(n_2145),
.B1(n_2153),
.B2(n_2146),
.Y(n_3109)
);

CKINVDCx11_ASAP7_75t_R g3110 ( 
.A(n_2522),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_2749),
.A2(n_2160),
.B1(n_2168),
.B2(n_2154),
.Y(n_3111)
);

INVx6_ASAP7_75t_L g3112 ( 
.A(n_2729),
.Y(n_3112)
);

CKINVDCx6p67_ASAP7_75t_R g3113 ( 
.A(n_2557),
.Y(n_3113)
);

CKINVDCx11_ASAP7_75t_R g3114 ( 
.A(n_2539),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2809),
.Y(n_3115)
);

AOI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_2764),
.A2(n_2384),
.B1(n_2207),
.B2(n_2363),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_2846),
.Y(n_3117)
);

AOI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2764),
.A2(n_2359),
.B1(n_2374),
.B2(n_2363),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2818),
.Y(n_3119)
);

AOI22xp33_ASAP7_75t_L g3120 ( 
.A1(n_2759),
.A2(n_2487),
.B1(n_2341),
.B2(n_2416),
.Y(n_3120)
);

OAI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2762),
.A2(n_2385),
.B1(n_2409),
.B2(n_2382),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2767),
.A2(n_2385),
.B1(n_2409),
.B2(n_2382),
.Y(n_3122)
);

BUFx6f_ASAP7_75t_L g3123 ( 
.A(n_2574),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_SL g3124 ( 
.A1(n_2719),
.A2(n_2321),
.B1(n_2473),
.B2(n_2437),
.Y(n_3124)
);

BUFx8_ASAP7_75t_L g3125 ( 
.A(n_2556),
.Y(n_3125)
);

BUFx12f_ASAP7_75t_L g3126 ( 
.A(n_2745),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2835),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_SL g3128 ( 
.A1(n_2719),
.A2(n_2321),
.B1(n_2117),
.B2(n_2288),
.Y(n_3128)
);

OAI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2767),
.A2(n_2144),
.B1(n_2431),
.B2(n_2140),
.Y(n_3129)
);

AOI22xp33_ASAP7_75t_L g3130 ( 
.A1(n_2766),
.A2(n_2078),
.B1(n_2111),
.B2(n_2094),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2842),
.Y(n_3131)
);

INVx4_ASAP7_75t_L g3132 ( 
.A(n_2846),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_L g3133 ( 
.A1(n_2779),
.A2(n_2496),
.B1(n_2498),
.B2(n_2495),
.Y(n_3133)
);

CKINVDCx6p67_ASAP7_75t_R g3134 ( 
.A(n_2694),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_2744),
.A2(n_2653),
.B1(n_2890),
.B2(n_2798),
.Y(n_3135)
);

AND2x4_ASAP7_75t_L g3136 ( 
.A(n_2581),
.B(n_2439),
.Y(n_3136)
);

BUFx2_ASAP7_75t_L g3137 ( 
.A(n_2771),
.Y(n_3137)
);

BUFx12f_ASAP7_75t_L g3138 ( 
.A(n_2532),
.Y(n_3138)
);

BUFx3_ASAP7_75t_L g3139 ( 
.A(n_2693),
.Y(n_3139)
);

BUFx2_ASAP7_75t_L g3140 ( 
.A(n_2771),
.Y(n_3140)
);

INVxp67_ASAP7_75t_SL g3141 ( 
.A(n_2650),
.Y(n_3141)
);

BUFx3_ASAP7_75t_L g3142 ( 
.A(n_2602),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2875),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2844),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2887),
.Y(n_3145)
);

INVx6_ASAP7_75t_L g3146 ( 
.A(n_2840),
.Y(n_3146)
);

INVxp67_ASAP7_75t_L g3147 ( 
.A(n_2736),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2577),
.Y(n_3148)
);

INVx1_ASAP7_75t_SL g3149 ( 
.A(n_2637),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_2653),
.A2(n_2495),
.B1(n_2498),
.B2(n_2496),
.Y(n_3150)
);

CKINVDCx16_ASAP7_75t_R g3151 ( 
.A(n_2751),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_2790),
.A2(n_2500),
.B1(n_2501),
.B2(n_2445),
.Y(n_3152)
);

BUFx10_ASAP7_75t_L g3153 ( 
.A(n_2531),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2847),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2856),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2577),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_2654),
.A2(n_2501),
.B1(n_2500),
.B2(n_2436),
.Y(n_3157)
);

BUFx2_ASAP7_75t_L g3158 ( 
.A(n_2691),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_SL g3159 ( 
.A1(n_2837),
.A2(n_2194),
.B(n_2182),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_SL g3160 ( 
.A1(n_2719),
.A2(n_2676),
.B1(n_2641),
.B2(n_2617),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2669),
.A2(n_2393),
.B1(n_2518),
.B2(n_2481),
.Y(n_3161)
);

OAI22xp5_ASAP7_75t_L g3162 ( 
.A1(n_2650),
.A2(n_2502),
.B1(n_2266),
.B2(n_2284),
.Y(n_3162)
);

CKINVDCx11_ASAP7_75t_R g3163 ( 
.A(n_2623),
.Y(n_3163)
);

BUFx8_ASAP7_75t_SL g3164 ( 
.A(n_2737),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2879),
.Y(n_3165)
);

BUFx12f_ASAP7_75t_L g3166 ( 
.A(n_2761),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2884),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_2574),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2804),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2807),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2814),
.Y(n_3171)
);

BUFx3_ASAP7_75t_L g3172 ( 
.A(n_2614),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2829),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_2750),
.B(n_2281),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2832),
.Y(n_3175)
);

AOI22xp33_ASAP7_75t_L g3176 ( 
.A1(n_2689),
.A2(n_2426),
.B1(n_2295),
.B2(n_2296),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2838),
.Y(n_3177)
);

NAND2x1p5_ASAP7_75t_L g3178 ( 
.A(n_2581),
.B(n_2232),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2619),
.Y(n_3179)
);

HB1xp67_ASAP7_75t_L g3180 ( 
.A(n_2860),
.Y(n_3180)
);

HB1xp67_ASAP7_75t_L g3181 ( 
.A(n_2865),
.Y(n_3181)
);

OAI22xp33_ASAP7_75t_L g3182 ( 
.A1(n_2676),
.A2(n_2289),
.B1(n_2351),
.B2(n_2336),
.Y(n_3182)
);

OAI22x1_ASAP7_75t_SL g3183 ( 
.A1(n_2626),
.A2(n_246),
.B1(n_243),
.B2(n_244),
.Y(n_3183)
);

OAI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_2676),
.A2(n_2352),
.B1(n_2365),
.B2(n_2354),
.Y(n_3184)
);

AOI22xp33_ASAP7_75t_SL g3185 ( 
.A1(n_2676),
.A2(n_2117),
.B1(n_2288),
.B2(n_2508),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2721),
.B(n_2367),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_SL g3187 ( 
.A(n_2617),
.B(n_2674),
.Y(n_3187)
);

INVx1_ASAP7_75t_SL g3188 ( 
.A(n_2542),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_2626),
.Y(n_3189)
);

CKINVDCx20_ASAP7_75t_R g3190 ( 
.A(n_2840),
.Y(n_3190)
);

OAI22xp33_ASAP7_75t_L g3191 ( 
.A1(n_2627),
.A2(n_2377),
.B1(n_2368),
.B2(n_2414),
.Y(n_3191)
);

AOI22xp33_ASAP7_75t_L g3192 ( 
.A1(n_2940),
.A2(n_2866),
.B1(n_2756),
.B2(n_2799),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2918),
.Y(n_3193)
);

OAI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_2929),
.A2(n_2695),
.B1(n_2697),
.B2(n_2627),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3060),
.B(n_2700),
.Y(n_3195)
);

INVx1_ASAP7_75t_SL g3196 ( 
.A(n_3180),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_3008),
.B(n_2892),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_L g3198 ( 
.A1(n_3080),
.A2(n_2789),
.B1(n_2811),
.B2(n_2548),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_3074),
.A2(n_2770),
.B1(n_2888),
.B2(n_2752),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_3032),
.B(n_2700),
.Y(n_3200)
);

AOI22xp5_ASAP7_75t_L g3201 ( 
.A1(n_3013),
.A2(n_2957),
.B1(n_2981),
.B2(n_2941),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_2936),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2923),
.Y(n_3203)
);

AOI22xp33_ASAP7_75t_SL g3204 ( 
.A1(n_2917),
.A2(n_2617),
.B1(n_2889),
.B2(n_2723),
.Y(n_3204)
);

OAI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_2954),
.A2(n_2617),
.B1(n_2697),
.B2(n_2695),
.Y(n_3205)
);

NOR2x1_ASAP7_75t_SL g3206 ( 
.A(n_2935),
.B(n_2581),
.Y(n_3206)
);

OAI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_2931),
.A2(n_2833),
.B1(n_2784),
.B2(n_2740),
.Y(n_3207)
);

AOI22xp33_ASAP7_75t_L g3208 ( 
.A1(n_2920),
.A2(n_2772),
.B1(n_2776),
.B2(n_2670),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_2963),
.Y(n_3209)
);

OAI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_2960),
.A2(n_2966),
.B1(n_2939),
.B2(n_2927),
.Y(n_3210)
);

AOI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_2974),
.A2(n_2780),
.B1(n_2845),
.B2(n_2843),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2924),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2925),
.Y(n_3213)
);

OAI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_2967),
.A2(n_2784),
.B1(n_2833),
.B2(n_2740),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2956),
.Y(n_3215)
);

OAI21xp33_ASAP7_75t_L g3216 ( 
.A1(n_3097),
.A2(n_2511),
.B(n_2872),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3181),
.B(n_2727),
.Y(n_3217)
);

AOI22xp33_ASAP7_75t_SL g3218 ( 
.A1(n_2919),
.A2(n_2705),
.B1(n_2568),
.B2(n_2572),
.Y(n_3218)
);

AOI22xp33_ASAP7_75t_L g3219 ( 
.A1(n_3004),
.A2(n_3089),
.B1(n_3055),
.B2(n_2996),
.Y(n_3219)
);

AOI22xp33_ASAP7_75t_L g3220 ( 
.A1(n_3057),
.A2(n_2876),
.B1(n_2877),
.B2(n_2862),
.Y(n_3220)
);

OAI22xp5_ASAP7_75t_L g3221 ( 
.A1(n_2976),
.A2(n_2649),
.B1(n_2872),
.B2(n_2827),
.Y(n_3221)
);

AOI22xp33_ASAP7_75t_L g3222 ( 
.A1(n_2905),
.A2(n_2897),
.B1(n_2883),
.B2(n_2743),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_L g3223 ( 
.A1(n_2922),
.A2(n_2841),
.B1(n_2820),
.B2(n_2827),
.Y(n_3223)
);

OAI21xp5_ASAP7_75t_SL g3224 ( 
.A1(n_2984),
.A2(n_2600),
.B(n_2598),
.Y(n_3224)
);

AOI22xp33_ASAP7_75t_L g3225 ( 
.A1(n_3135),
.A2(n_2808),
.B1(n_2815),
.B2(n_2812),
.Y(n_3225)
);

BUFx4f_ASAP7_75t_SL g3226 ( 
.A(n_2915),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_3010),
.B(n_2727),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_SL g3228 ( 
.A1(n_3091),
.A2(n_3112),
.B1(n_2937),
.B2(n_2950),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2987),
.Y(n_3229)
);

AOI22xp33_ASAP7_75t_L g3230 ( 
.A1(n_2934),
.A2(n_2864),
.B1(n_2721),
.B2(n_2830),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2989),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_SL g3232 ( 
.A(n_2958),
.B(n_2674),
.Y(n_3232)
);

OAI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_3118),
.A2(n_2649),
.B1(n_2864),
.B2(n_2893),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2969),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_L g3235 ( 
.A1(n_2943),
.A2(n_2864),
.B1(n_2830),
.B2(n_2852),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_2937),
.Y(n_3236)
);

AOI22xp33_ASAP7_75t_L g3237 ( 
.A1(n_3001),
.A2(n_2852),
.B1(n_2831),
.B2(n_2869),
.Y(n_3237)
);

OAI21xp5_ASAP7_75t_SL g3238 ( 
.A1(n_2930),
.A2(n_2600),
.B(n_2598),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2970),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2979),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_2991),
.Y(n_3241)
);

AOI22xp33_ASAP7_75t_SL g3242 ( 
.A1(n_3091),
.A2(n_2831),
.B1(n_2604),
.B2(n_2533),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3072),
.A2(n_2869),
.B1(n_2709),
.B2(n_2716),
.Y(n_3243)
);

AOI22xp33_ASAP7_75t_SL g3244 ( 
.A1(n_3112),
.A2(n_2604),
.B1(n_2533),
.B2(n_2588),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_L g3245 ( 
.A1(n_3006),
.A2(n_2714),
.B1(n_2738),
.B2(n_2704),
.Y(n_3245)
);

AOI222xp33_ASAP7_75t_L g3246 ( 
.A1(n_3183),
.A2(n_2781),
.B1(n_2712),
.B2(n_2559),
.C1(n_2551),
.C2(n_2665),
.Y(n_3246)
);

CKINVDCx20_ASAP7_75t_R g3247 ( 
.A(n_2938),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_L g3248 ( 
.A(n_2993),
.B(n_2618),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3000),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2983),
.Y(n_3250)
);

INVx3_ASAP7_75t_L g3251 ( 
.A(n_2942),
.Y(n_3251)
);

AOI22xp33_ASAP7_75t_L g3252 ( 
.A1(n_2995),
.A2(n_2704),
.B1(n_2528),
.B2(n_2538),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3021),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3061),
.B(n_2667),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2998),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_3099),
.A2(n_2528),
.B1(n_2538),
.B2(n_2698),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_2903),
.A2(n_2781),
.B1(n_2680),
.B2(n_2855),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2900),
.B(n_2851),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3035),
.B(n_2619),
.Y(n_3259)
);

INVx2_ASAP7_75t_SL g3260 ( 
.A(n_2935),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3033),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2955),
.B(n_2549),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3038),
.B(n_2632),
.Y(n_3263)
);

OAI21xp5_ASAP7_75t_SL g3264 ( 
.A1(n_3069),
.A2(n_2588),
.B(n_2542),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3041),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3047),
.B(n_2632),
.Y(n_3266)
);

CKINVDCx20_ASAP7_75t_R g3267 ( 
.A(n_2933),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_L g3268 ( 
.A1(n_2985),
.A2(n_3116),
.B1(n_2910),
.B2(n_2907),
.Y(n_3268)
);

AOI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_3024),
.A2(n_2786),
.B1(n_2871),
.B2(n_2599),
.Y(n_3269)
);

INVx3_ASAP7_75t_L g3270 ( 
.A(n_2942),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3048),
.B(n_2687),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3170),
.B(n_2585),
.Y(n_3272)
);

AOI22xp33_ASAP7_75t_L g3273 ( 
.A1(n_2945),
.A2(n_2786),
.B1(n_2871),
.B2(n_2855),
.Y(n_3273)
);

INVx4_ASAP7_75t_L g3274 ( 
.A(n_2935),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_2902),
.Y(n_3275)
);

INVx4_ASAP7_75t_L g3276 ( 
.A(n_2901),
.Y(n_3276)
);

OAI222xp33_ASAP7_75t_L g3277 ( 
.A1(n_3149),
.A2(n_2893),
.B1(n_2671),
.B2(n_2895),
.C1(n_2680),
.C2(n_2683),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3053),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3058),
.Y(n_3279)
);

OAI222xp33_ASAP7_75t_L g3280 ( 
.A1(n_2997),
.A2(n_2893),
.B1(n_2671),
.B2(n_2895),
.C1(n_2683),
.C2(n_2702),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_3046),
.A2(n_2658),
.B1(n_2712),
.B2(n_2571),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3059),
.Y(n_3282)
);

CKINVDCx20_ASAP7_75t_R g3283 ( 
.A(n_2944),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3083),
.Y(n_3284)
);

BUFx12f_ASAP7_75t_L g3285 ( 
.A(n_3014),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_2914),
.A2(n_2571),
.B1(n_2559),
.B2(n_2551),
.Y(n_3286)
);

HB1xp67_ASAP7_75t_L g3287 ( 
.A(n_3148),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3186),
.B(n_2687),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3156),
.Y(n_3289)
);

AOI22xp33_ASAP7_75t_L g3290 ( 
.A1(n_3068),
.A2(n_2668),
.B1(n_2702),
.B2(n_2742),
.Y(n_3290)
);

INVx4_ASAP7_75t_L g3291 ( 
.A(n_2901),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3018),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_2950),
.Y(n_3293)
);

CKINVDCx6p67_ASAP7_75t_R g3294 ( 
.A(n_2971),
.Y(n_3294)
);

AOI22xp33_ASAP7_75t_L g3295 ( 
.A1(n_3034),
.A2(n_2747),
.B1(n_2748),
.B2(n_2742),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_3092),
.A2(n_2748),
.B1(n_2747),
.B2(n_2753),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3018),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3020),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3020),
.Y(n_3299)
);

AOI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_2972),
.A2(n_3005),
.B1(n_2978),
.B2(n_3109),
.Y(n_3300)
);

HB1xp67_ASAP7_75t_L g3301 ( 
.A(n_3169),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3040),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_3150),
.A2(n_2753),
.B1(n_2535),
.B2(n_2848),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3044),
.B(n_2711),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3049),
.B(n_2592),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3023),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3064),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_2988),
.A2(n_2535),
.B1(n_2848),
.B2(n_2639),
.Y(n_3308)
);

OAI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_3022),
.A2(n_2643),
.B1(n_2647),
.B2(n_2648),
.Y(n_3309)
);

NOR3xp33_ASAP7_75t_L g3310 ( 
.A(n_3096),
.B(n_2773),
.C(n_2731),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3066),
.Y(n_3311)
);

BUFx2_ASAP7_75t_L g3312 ( 
.A(n_3117),
.Y(n_3312)
);

AOI22xp33_ASAP7_75t_L g3313 ( 
.A1(n_2932),
.A2(n_2535),
.B1(n_2639),
.B2(n_2593),
.Y(n_3313)
);

AOI22xp33_ASAP7_75t_SL g3314 ( 
.A1(n_2911),
.A2(n_2688),
.B1(n_2674),
.B2(n_2657),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_3171),
.Y(n_3315)
);

AOI22xp33_ASAP7_75t_SL g3316 ( 
.A1(n_3146),
.A2(n_3036),
.B1(n_3140),
.B2(n_3137),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3176),
.A2(n_2647),
.B1(n_2643),
.B2(n_2648),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3081),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_SL g3319 ( 
.A1(n_3146),
.A2(n_2674),
.B1(n_2688),
.B2(n_2657),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_SL g3320 ( 
.A1(n_3036),
.A2(n_2688),
.B1(n_2674),
.B2(n_2787),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3093),
.A2(n_2535),
.B1(n_2593),
.B2(n_2731),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_3143),
.A2(n_2535),
.B1(n_2773),
.B2(n_2810),
.Y(n_3322)
);

AOI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_3145),
.A2(n_2810),
.B1(n_2760),
.B2(n_2688),
.Y(n_3323)
);

AOI22xp33_ASAP7_75t_L g3324 ( 
.A1(n_3157),
.A2(n_2688),
.B1(n_2616),
.B2(n_2565),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_3023),
.B(n_2592),
.Y(n_3325)
);

OAI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3007),
.A2(n_2787),
.B1(n_2795),
.B2(n_2596),
.Y(n_3326)
);

OAI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_2904),
.A2(n_2720),
.B1(n_2739),
.B2(n_2711),
.Y(n_3327)
);

INVx2_ASAP7_75t_SL g3328 ( 
.A(n_2994),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_2951),
.B(n_2795),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3151),
.B(n_2596),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_2916),
.A2(n_2678),
.B1(n_2576),
.B2(n_2590),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3073),
.Y(n_3332)
);

OAI22xp33_ASAP7_75t_L g3333 ( 
.A1(n_3017),
.A2(n_3029),
.B1(n_3188),
.B2(n_3132),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3084),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3173),
.A2(n_2678),
.B1(n_2576),
.B2(n_2590),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_3175),
.A2(n_2826),
.B1(n_2625),
.B2(n_2821),
.Y(n_3336)
);

INVxp67_ASAP7_75t_L g3337 ( 
.A(n_3027),
.Y(n_3337)
);

OAI22xp33_ASAP7_75t_SL g3338 ( 
.A1(n_3147),
.A2(n_2715),
.B1(n_2826),
.B2(n_2821),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3073),
.Y(n_3339)
);

INVx4_ASAP7_75t_L g3340 ( 
.A(n_3132),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_SL g3341 ( 
.A1(n_3036),
.A2(n_2720),
.B1(n_2739),
.B2(n_2715),
.Y(n_3341)
);

AOI22xp33_ASAP7_75t_L g3342 ( 
.A1(n_3177),
.A2(n_2625),
.B1(n_2859),
.B2(n_2797),
.Y(n_3342)
);

BUFx5_ASAP7_75t_L g3343 ( 
.A(n_3136),
.Y(n_3343)
);

BUFx3_ASAP7_75t_L g3344 ( 
.A(n_3003),
.Y(n_3344)
);

BUFx4f_ASAP7_75t_SL g3345 ( 
.A(n_2906),
.Y(n_3345)
);

CKINVDCx11_ASAP7_75t_R g3346 ( 
.A(n_2999),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_SL g3347 ( 
.A1(n_3078),
.A2(n_2797),
.B1(n_2859),
.B2(n_2788),
.Y(n_3347)
);

OAI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_2904),
.A2(n_2908),
.B1(n_2913),
.B2(n_2912),
.Y(n_3348)
);

BUFx2_ASAP7_75t_L g3349 ( 
.A(n_3039),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3094),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3110),
.A2(n_2640),
.B1(n_2644),
.B2(n_2426),
.Y(n_3351)
);

INVx1_ASAP7_75t_SL g3352 ( 
.A(n_2909),
.Y(n_3352)
);

OAI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_2908),
.A2(n_2612),
.B1(n_2788),
.B2(n_2735),
.Y(n_3353)
);

OAI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3016),
.A2(n_2788),
.B1(n_2612),
.B2(n_2735),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_L g3355 ( 
.A1(n_2912),
.A2(n_2238),
.B1(n_2255),
.B2(n_2117),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3098),
.Y(n_3356)
);

NOR2x1_ASAP7_75t_L g3357 ( 
.A(n_3190),
.B(n_2817),
.Y(n_3357)
);

INVx3_ASAP7_75t_SL g3358 ( 
.A(n_3003),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_2913),
.A2(n_2961),
.B1(n_2992),
.B2(n_2962),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_SL g3360 ( 
.A1(n_3078),
.A2(n_2733),
.B1(n_2746),
.B2(n_2732),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3094),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_2961),
.A2(n_2117),
.B1(n_2126),
.B2(n_2106),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_SL g3363 ( 
.A1(n_3108),
.A2(n_2733),
.B1(n_2746),
.B2(n_2732),
.Y(n_3363)
);

OAI21xp33_ASAP7_75t_L g3364 ( 
.A1(n_3120),
.A2(n_2853),
.B(n_2796),
.Y(n_3364)
);

OAI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_3085),
.A2(n_2414),
.B(n_2453),
.Y(n_3365)
);

NOR2xp33_ASAP7_75t_L g3366 ( 
.A(n_2986),
.B(n_244),
.Y(n_3366)
);

BUFx3_ASAP7_75t_L g3367 ( 
.A(n_3087),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_2962),
.A2(n_2106),
.B1(n_2184),
.B2(n_2126),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3165),
.B(n_2732),
.Y(n_3369)
);

OAI21xp33_ASAP7_75t_L g3370 ( 
.A1(n_3086),
.A2(n_3111),
.B(n_2990),
.Y(n_3370)
);

OAI21xp5_ASAP7_75t_SL g3371 ( 
.A1(n_3160),
.A2(n_2853),
.B(n_2796),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3103),
.Y(n_3372)
);

AOI22xp33_ASAP7_75t_L g3373 ( 
.A1(n_2992),
.A2(n_2215),
.B1(n_2219),
.B2(n_2184),
.Y(n_3373)
);

CKINVDCx5p33_ASAP7_75t_R g3374 ( 
.A(n_3164),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3015),
.A2(n_2219),
.B1(n_2240),
.B2(n_2215),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3015),
.A2(n_2264),
.B1(n_2240),
.B2(n_2508),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_3100),
.A2(n_2264),
.B1(n_2519),
.B2(n_2514),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3105),
.Y(n_3378)
);

OAI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3113),
.A2(n_2733),
.B1(n_2746),
.B2(n_2732),
.Y(n_3379)
);

AOI222xp33_ASAP7_75t_L g3380 ( 
.A1(n_3138),
.A2(n_249),
.B1(n_252),
.B2(n_247),
.C1(n_248),
.C2(n_250),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_3063),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_L g3382 ( 
.A1(n_3043),
.A2(n_2519),
.B1(n_2514),
.B2(n_2344),
.Y(n_3382)
);

BUFx5_ASAP7_75t_L g3383 ( 
.A(n_3136),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3167),
.B(n_2733),
.Y(n_3384)
);

CKINVDCx11_ASAP7_75t_R g3385 ( 
.A(n_3054),
.Y(n_3385)
);

OAI21xp33_ASAP7_75t_L g3386 ( 
.A1(n_3076),
.A2(n_2474),
.B(n_2458),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_3079),
.A2(n_2344),
.B1(n_2348),
.B2(n_2340),
.Y(n_3387)
);

HB1xp67_ASAP7_75t_L g3388 ( 
.A(n_3103),
.Y(n_3388)
);

INVx5_ASAP7_75t_SL g3389 ( 
.A(n_3134),
.Y(n_3389)
);

BUFx3_ASAP7_75t_L g3390 ( 
.A(n_3087),
.Y(n_3390)
);

OAI21xp5_ASAP7_75t_SL g3391 ( 
.A1(n_3028),
.A2(n_2344),
.B(n_2340),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_3179),
.A2(n_2348),
.B1(n_2355),
.B2(n_2340),
.Y(n_3392)
);

INVx4_ASAP7_75t_R g3393 ( 
.A(n_2928),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3115),
.B(n_2746),
.Y(n_3394)
);

BUFx12f_ASAP7_75t_L g3395 ( 
.A(n_2973),
.Y(n_3395)
);

AOI222xp33_ASAP7_75t_L g3396 ( 
.A1(n_2973),
.A2(n_3026),
.B1(n_2968),
.B2(n_3052),
.C1(n_3189),
.C2(n_3107),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_SL g3397 ( 
.A1(n_3108),
.A2(n_3071),
.B1(n_3082),
.B2(n_3077),
.Y(n_3397)
);

OAI222xp33_ASAP7_75t_L g3398 ( 
.A1(n_3104),
.A2(n_2778),
.B1(n_250),
.B2(n_253),
.C1(n_248),
.C2(n_249),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3174),
.B(n_252),
.Y(n_3399)
);

INVx2_ASAP7_75t_SL g3400 ( 
.A(n_2971),
.Y(n_3400)
);

BUFx12f_ASAP7_75t_L g3401 ( 
.A(n_3075),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3115),
.B(n_2778),
.Y(n_3402)
);

AOI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3179),
.A2(n_2355),
.B1(n_2388),
.B2(n_2348),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_SL g3404 ( 
.A1(n_3063),
.A2(n_2778),
.B1(n_2899),
.B2(n_2578),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3153),
.B(n_253),
.Y(n_3405)
);

OAI22xp5_ASAP7_75t_L g3406 ( 
.A1(n_3121),
.A2(n_2778),
.B1(n_2388),
.B2(n_2355),
.Y(n_3406)
);

INVxp67_ASAP7_75t_SL g3407 ( 
.A(n_2926),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_SL g3408 ( 
.A1(n_3077),
.A2(n_2574),
.B1(n_2579),
.B2(n_2578),
.Y(n_3408)
);

CKINVDCx11_ASAP7_75t_R g3409 ( 
.A(n_3067),
.Y(n_3409)
);

AOI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_3122),
.A2(n_2388),
.B1(n_2474),
.B2(n_2458),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3106),
.Y(n_3411)
);

AOI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_3161),
.A2(n_2458),
.B1(n_2486),
.B2(n_2474),
.Y(n_3412)
);

AOI222xp33_ASAP7_75t_L g3413 ( 
.A1(n_3002),
.A2(n_256),
.B1(n_258),
.B2(n_254),
.C1(n_255),
.C2(n_257),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_3090),
.Y(n_3414)
);

INVxp67_ASAP7_75t_L g3415 ( 
.A(n_3158),
.Y(n_3415)
);

AOI22xp33_ASAP7_75t_L g3416 ( 
.A1(n_3002),
.A2(n_2492),
.B1(n_2503),
.B2(n_2486),
.Y(n_3416)
);

BUFx2_ASAP7_75t_L g3417 ( 
.A(n_3009),
.Y(n_3417)
);

OAI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3141),
.A2(n_2492),
.B1(n_2503),
.B2(n_2486),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3119),
.B(n_2492),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3127),
.B(n_2503),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3131),
.B(n_2578),
.Y(n_3421)
);

CKINVDCx5p33_ASAP7_75t_R g3422 ( 
.A(n_3114),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3070),
.A2(n_3030),
.B1(n_2952),
.B2(n_3125),
.Y(n_3423)
);

OAI221xp5_ASAP7_75t_L g3424 ( 
.A1(n_3219),
.A2(n_3133),
.B1(n_3130),
.B2(n_3012),
.C(n_3095),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3246),
.A2(n_3216),
.B1(n_3210),
.B2(n_3268),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_3246),
.A2(n_3042),
.B1(n_3011),
.B2(n_3166),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3380),
.A2(n_3042),
.B1(n_3011),
.B2(n_3152),
.Y(n_3427)
);

OAI221xp5_ASAP7_75t_L g3428 ( 
.A1(n_3201),
.A2(n_2953),
.B1(n_3065),
.B2(n_3172),
.C(n_3142),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3380),
.A2(n_3125),
.B1(n_3037),
.B2(n_3031),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3229),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3215),
.Y(n_3431)
);

OAI22xp5_ASAP7_75t_L g3432 ( 
.A1(n_3230),
.A2(n_3264),
.B1(n_3290),
.B2(n_3198),
.Y(n_3432)
);

OAI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3398),
.A2(n_3129),
.B(n_3162),
.Y(n_3433)
);

AOI22xp33_ASAP7_75t_L g3434 ( 
.A1(n_3223),
.A2(n_3037),
.B1(n_3031),
.B2(n_3144),
.Y(n_3434)
);

OAI222xp33_ASAP7_75t_L g3435 ( 
.A1(n_3207),
.A2(n_3314),
.B1(n_3397),
.B2(n_3196),
.C1(n_3205),
.C2(n_3291),
.Y(n_3435)
);

AOI22xp33_ASAP7_75t_SL g3436 ( 
.A1(n_3207),
.A2(n_3045),
.B1(n_2977),
.B2(n_3153),
.Y(n_3436)
);

AOI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3300),
.A2(n_2964),
.B1(n_3056),
.B2(n_3163),
.Y(n_3437)
);

AOI22xp33_ASAP7_75t_L g3438 ( 
.A1(n_3220),
.A2(n_3155),
.B1(n_3154),
.B2(n_2946),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_3226),
.B(n_3050),
.Y(n_3439)
);

NOR3xp33_ASAP7_75t_SL g3440 ( 
.A(n_3264),
.B(n_2947),
.C(n_3187),
.Y(n_3440)
);

AOI222xp33_ASAP7_75t_L g3441 ( 
.A1(n_3370),
.A2(n_3296),
.B1(n_3276),
.B2(n_3291),
.C1(n_3199),
.C2(n_3222),
.Y(n_3441)
);

OAI211xp5_ASAP7_75t_SL g3442 ( 
.A1(n_3396),
.A2(n_3124),
.B(n_3128),
.C(n_2975),
.Y(n_3442)
);

OAI21xp33_ASAP7_75t_L g3443 ( 
.A1(n_3211),
.A2(n_3139),
.B(n_3101),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_L g3444 ( 
.A1(n_3221),
.A2(n_2949),
.B1(n_2921),
.B2(n_2948),
.Y(n_3444)
);

AOI22xp33_ASAP7_75t_L g3445 ( 
.A1(n_3413),
.A2(n_2949),
.B1(n_2921),
.B2(n_2959),
.Y(n_3445)
);

OA21x2_ASAP7_75t_L g3446 ( 
.A1(n_3365),
.A2(n_2982),
.B(n_3184),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3413),
.A2(n_2949),
.B1(n_2921),
.B2(n_3051),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3200),
.A2(n_3182),
.B1(n_3191),
.B2(n_3185),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3234),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3227),
.B(n_2965),
.Y(n_3450)
);

AOI22xp33_ASAP7_75t_L g3451 ( 
.A1(n_3273),
.A2(n_2964),
.B1(n_3178),
.B2(n_2980),
.Y(n_3451)
);

AOI222xp33_ASAP7_75t_L g3452 ( 
.A1(n_3276),
.A2(n_3126),
.B1(n_3102),
.B2(n_256),
.C1(n_259),
.C2(n_254),
.Y(n_3452)
);

OAI221xp5_ASAP7_75t_L g3453 ( 
.A1(n_3192),
.A2(n_3159),
.B1(n_3168),
.B2(n_3019),
.C(n_3025),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3269),
.A2(n_2980),
.B1(n_3019),
.B2(n_2965),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_3258),
.A2(n_2980),
.B1(n_3019),
.B2(n_2965),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3197),
.B(n_3025),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3252),
.A2(n_3310),
.B1(n_3243),
.B2(n_3281),
.Y(n_3457)
);

AOI22xp33_ASAP7_75t_L g3458 ( 
.A1(n_3205),
.A2(n_3062),
.B1(n_3088),
.B2(n_3025),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_3308),
.A2(n_3088),
.B1(n_3123),
.B2(n_3062),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3286),
.A2(n_3102),
.B1(n_3088),
.B2(n_3062),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3295),
.A2(n_3168),
.B1(n_3123),
.B2(n_2633),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3193),
.B(n_3196),
.Y(n_3462)
);

OAI22xp5_ASAP7_75t_SL g3463 ( 
.A1(n_3267),
.A2(n_3168),
.B1(n_3123),
.B2(n_2633),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3313),
.A2(n_2633),
.B1(n_2684),
.B2(n_2579),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3217),
.B(n_255),
.Y(n_3465)
);

AOI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3214),
.A2(n_2684),
.B1(n_2707),
.B2(n_2579),
.Y(n_3466)
);

NAND3xp33_ASAP7_75t_L g3467 ( 
.A(n_3366),
.B(n_2707),
.C(n_2684),
.Y(n_3467)
);

AOI22xp33_ASAP7_75t_L g3468 ( 
.A1(n_3237),
.A2(n_2783),
.B1(n_2800),
.B2(n_2707),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3233),
.A2(n_2800),
.B1(n_2822),
.B2(n_2783),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3203),
.B(n_257),
.Y(n_3470)
);

INVx4_ASAP7_75t_L g3471 ( 
.A(n_3274),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3327),
.A2(n_2800),
.B1(n_2822),
.B2(n_2783),
.Y(n_3472)
);

OAI222xp33_ASAP7_75t_L g3473 ( 
.A1(n_3349),
.A2(n_261),
.B1(n_263),
.B2(n_259),
.C1(n_260),
.C2(n_262),
.Y(n_3473)
);

AOI22xp5_ASAP7_75t_L g3474 ( 
.A1(n_3257),
.A2(n_2822),
.B1(n_2878),
.B2(n_2849),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3327),
.A2(n_2878),
.B1(n_2882),
.B2(n_2849),
.Y(n_3475)
);

OAI221xp5_ASAP7_75t_SL g3476 ( 
.A1(n_3224),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.C(n_264),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3212),
.B(n_264),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3231),
.Y(n_3478)
);

OAI222xp33_ASAP7_75t_L g3479 ( 
.A1(n_3340),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.C1(n_268),
.C2(n_269),
.Y(n_3479)
);

OAI221xp5_ASAP7_75t_SL g3480 ( 
.A1(n_3224),
.A2(n_268),
.B1(n_265),
.B2(n_266),
.C(n_269),
.Y(n_3480)
);

OAI22xp5_ASAP7_75t_L g3481 ( 
.A1(n_3244),
.A2(n_2878),
.B1(n_2882),
.B2(n_2849),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3256),
.A2(n_2899),
.B1(n_2882),
.B2(n_2182),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3245),
.A2(n_2899),
.B1(n_2194),
.B2(n_2247),
.Y(n_3483)
);

OAI22xp5_ASAP7_75t_SL g3484 ( 
.A1(n_3345),
.A2(n_2226),
.B1(n_2247),
.B2(n_2194),
.Y(n_3484)
);

OAI221xp5_ASAP7_75t_L g3485 ( 
.A1(n_3208),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.C(n_273),
.Y(n_3485)
);

AOI222xp33_ASAP7_75t_SL g3486 ( 
.A1(n_3337),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.C1(n_274),
.C2(n_275),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3305),
.B(n_274),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3213),
.B(n_275),
.Y(n_3488)
);

AOI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3225),
.A2(n_2226),
.B1(n_2273),
.B2(n_2247),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_L g3490 ( 
.A1(n_3301),
.A2(n_3315),
.B1(n_3399),
.B2(n_3340),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3194),
.A2(n_2226),
.B1(n_2273),
.B2(n_1950),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3241),
.Y(n_3492)
);

NAND2xp33_ASAP7_75t_SL g3493 ( 
.A(n_3274),
.B(n_2273),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_L g3494 ( 
.A1(n_3304),
.A2(n_3312),
.B1(n_3235),
.B2(n_3367),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_SL g3495 ( 
.A(n_3294),
.B(n_3390),
.Y(n_3495)
);

AOI22xp33_ASAP7_75t_L g3496 ( 
.A1(n_3303),
.A2(n_1950),
.B1(n_278),
.B2(n_276),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3284),
.B(n_276),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_SL g3498 ( 
.A1(n_3338),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3239),
.B(n_277),
.Y(n_3499)
);

INVxp67_ASAP7_75t_L g3500 ( 
.A(n_3417),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3240),
.B(n_279),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3272),
.B(n_280),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3249),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3324),
.A2(n_284),
.B1(n_281),
.B2(n_282),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_SL g3505 ( 
.A1(n_3236),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3262),
.B(n_285),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3388),
.B(n_287),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_SL g3508 ( 
.A1(n_3236),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3331),
.A2(n_3330),
.B1(n_3287),
.B2(n_3248),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_3333),
.A2(n_291),
.B1(n_288),
.B2(n_289),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_L g3511 ( 
.A1(n_3405),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3250),
.B(n_292),
.Y(n_3512)
);

AOI22xp33_ASAP7_75t_L g3513 ( 
.A1(n_3323),
.A2(n_297),
.B1(n_294),
.B2(n_295),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3255),
.B(n_294),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3265),
.B(n_298),
.Y(n_3515)
);

OA21x2_ASAP7_75t_L g3516 ( 
.A1(n_3365),
.A2(n_586),
.B(n_585),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3335),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3278),
.B(n_300),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3279),
.B(n_3282),
.Y(n_3519)
);

AOI22xp33_ASAP7_75t_L g3520 ( 
.A1(n_3232),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_L g3521 ( 
.A1(n_3322),
.A2(n_304),
.B1(n_301),
.B2(n_303),
.Y(n_3521)
);

AOI22xp33_ASAP7_75t_L g3522 ( 
.A1(n_3289),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3411),
.B(n_305),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_SL g3524 ( 
.A1(n_3251),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3321),
.A2(n_3369),
.B1(n_3384),
.B2(n_3309),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3329),
.A2(n_310),
.B1(n_307),
.B2(n_309),
.Y(n_3526)
);

AOI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3394),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_3527)
);

OAI22xp33_ASAP7_75t_L g3528 ( 
.A1(n_3371),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3325),
.B(n_314),
.Y(n_3529)
);

AOI22xp33_ASAP7_75t_SL g3530 ( 
.A1(n_3251),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_3530)
);

NOR3xp33_ASAP7_75t_L g3531 ( 
.A(n_3415),
.B(n_317),
.C(n_318),
.Y(n_3531)
);

AOI22xp33_ASAP7_75t_L g3532 ( 
.A1(n_3402),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3228),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.Y(n_3533)
);

AOI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_3317),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_3534)
);

AOI22xp33_ASAP7_75t_L g3535 ( 
.A1(n_3396),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_3535)
);

AOI22xp33_ASAP7_75t_L g3536 ( 
.A1(n_3288),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3395),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3253),
.B(n_333),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3292),
.Y(n_3539)
);

AOI22xp33_ASAP7_75t_L g3540 ( 
.A1(n_3254),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3297),
.B(n_337),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3261),
.B(n_3302),
.Y(n_3542)
);

NAND3xp33_ASAP7_75t_L g3543 ( 
.A(n_3316),
.B(n_337),
.C(n_338),
.Y(n_3543)
);

OAI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3371),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3298),
.B(n_3299),
.Y(n_3545)
);

OAI222xp33_ASAP7_75t_L g3546 ( 
.A1(n_3319),
.A2(n_339),
.B1(n_342),
.B2(n_343),
.C1(n_344),
.C2(n_345),
.Y(n_3546)
);

AOI22xp33_ASAP7_75t_SL g3547 ( 
.A1(n_3270),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3307),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3348),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_3549)
);

AOI22xp33_ASAP7_75t_L g3550 ( 
.A1(n_3271),
.A2(n_352),
.B1(n_349),
.B2(n_351),
.Y(n_3550)
);

AOI22xp5_ASAP7_75t_L g3551 ( 
.A1(n_3270),
.A2(n_3293),
.B1(n_3238),
.B2(n_3260),
.Y(n_3551)
);

AO22x1_ASAP7_75t_L g3552 ( 
.A1(n_3358),
.A2(n_354),
.B1(n_351),
.B2(n_353),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3348),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3553)
);

OAI22xp5_ASAP7_75t_L g3554 ( 
.A1(n_3293),
.A2(n_3218),
.B1(n_3389),
.B2(n_3242),
.Y(n_3554)
);

AOI22xp33_ASAP7_75t_L g3555 ( 
.A1(n_3364),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_3555)
);

OAI22xp5_ASAP7_75t_L g3556 ( 
.A1(n_3389),
.A2(n_360),
.B1(n_357),
.B2(n_358),
.Y(n_3556)
);

OAI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_3389),
.A2(n_3341),
.B1(n_3320),
.B2(n_3377),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3381),
.A2(n_362),
.B1(n_358),
.B2(n_360),
.Y(n_3558)
);

OAI221xp5_ASAP7_75t_SL g3559 ( 
.A1(n_3238),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.C(n_365),
.Y(n_3559)
);

AOI22xp5_ASAP7_75t_SL g3560 ( 
.A1(n_3247),
.A2(n_367),
.B1(n_363),
.B2(n_365),
.Y(n_3560)
);

AOI222xp33_ASAP7_75t_L g3561 ( 
.A1(n_3401),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.C1(n_370),
.C2(n_371),
.Y(n_3561)
);

AOI22xp33_ASAP7_75t_L g3562 ( 
.A1(n_3381),
.A2(n_371),
.B1(n_368),
.B2(n_370),
.Y(n_3562)
);

AOI22xp33_ASAP7_75t_L g3563 ( 
.A1(n_3359),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_3563)
);

OAI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3391),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_3564)
);

OAI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3391),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_3565)
);

AOI22xp33_ASAP7_75t_SL g3566 ( 
.A1(n_3206),
.A2(n_378),
.B1(n_375),
.B2(n_377),
.Y(n_3566)
);

AOI221xp5_ASAP7_75t_L g3567 ( 
.A1(n_3195),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.C(n_383),
.Y(n_3567)
);

OAI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3347),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3306),
.Y(n_3569)
);

AOI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3332),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3339),
.Y(n_3571)
);

AOI22xp33_ASAP7_75t_L g3572 ( 
.A1(n_3350),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3361),
.B(n_389),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3283),
.B(n_389),
.Y(n_3574)
);

OAI221xp5_ASAP7_75t_L g3575 ( 
.A1(n_3423),
.A2(n_3351),
.B1(n_3342),
.B2(n_3336),
.C(n_3357),
.Y(n_3575)
);

OAI22xp5_ASAP7_75t_L g3576 ( 
.A1(n_3360),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_3576)
);

OAI21xp5_ASAP7_75t_SL g3577 ( 
.A1(n_3436),
.A2(n_3277),
.B(n_3280),
.Y(n_3577)
);

NAND4xp25_ASAP7_75t_L g3578 ( 
.A(n_3425),
.B(n_3209),
.C(n_3382),
.D(n_3373),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_3554),
.B(n_3326),
.Y(n_3579)
);

AND2x2_ASAP7_75t_SL g3580 ( 
.A(n_3471),
.B(n_3393),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_3471),
.B(n_3408),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3519),
.B(n_3372),
.Y(n_3582)
);

OAI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_3429),
.A2(n_3204),
.B1(n_3363),
.B2(n_3414),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3456),
.B(n_3407),
.Y(n_3584)
);

AOI221xp5_ASAP7_75t_L g3585 ( 
.A1(n_3426),
.A2(n_3259),
.B1(n_3263),
.B2(n_3266),
.C(n_3352),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3542),
.B(n_3311),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3431),
.B(n_3318),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3449),
.B(n_3334),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3462),
.B(n_3352),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3539),
.B(n_3356),
.Y(n_3590)
);

OAI21xp5_ASAP7_75t_SL g3591 ( 
.A1(n_3452),
.A2(n_3379),
.B(n_3400),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3450),
.B(n_3378),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3500),
.B(n_3343),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_3509),
.B(n_3430),
.Y(n_3594)
);

NAND3xp33_ASAP7_75t_L g3595 ( 
.A(n_3426),
.B(n_3353),
.C(n_3404),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3569),
.B(n_3343),
.Y(n_3596)
);

OAI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3429),
.A2(n_3414),
.B1(n_3353),
.B2(n_3416),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3571),
.B(n_3343),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3545),
.B(n_3343),
.Y(n_3599)
);

NAND3xp33_ASAP7_75t_L g3600 ( 
.A(n_3441),
.B(n_3375),
.C(n_3368),
.Y(n_3600)
);

OAI221xp5_ASAP7_75t_L g3601 ( 
.A1(n_3535),
.A2(n_3344),
.B1(n_3422),
.B2(n_3328),
.C(n_3374),
.Y(n_3601)
);

AOI221xp5_ASAP7_75t_L g3602 ( 
.A1(n_3432),
.A2(n_3535),
.B1(n_3544),
.B2(n_3528),
.C(n_3473),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3478),
.B(n_3343),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3492),
.B(n_3383),
.Y(n_3604)
);

OA21x2_ASAP7_75t_L g3605 ( 
.A1(n_3435),
.A2(n_3386),
.B(n_3421),
.Y(n_3605)
);

OAI21xp5_ASAP7_75t_SL g3606 ( 
.A1(n_3561),
.A2(n_3354),
.B(n_3406),
.Y(n_3606)
);

NAND4xp25_ASAP7_75t_SL g3607 ( 
.A(n_3437),
.B(n_3285),
.C(n_3385),
.D(n_3346),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3503),
.B(n_3383),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3548),
.B(n_3383),
.Y(n_3609)
);

OAI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3528),
.A2(n_3420),
.B(n_3419),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3490),
.B(n_3383),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3507),
.Y(n_3612)
);

OAI221xp5_ASAP7_75t_L g3613 ( 
.A1(n_3494),
.A2(n_3376),
.B1(n_3275),
.B2(n_3202),
.C(n_3355),
.Y(n_3613)
);

OAI221xp5_ASAP7_75t_L g3614 ( 
.A1(n_3494),
.A2(n_3427),
.B1(n_3447),
.B2(n_3537),
.C(n_3457),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3490),
.B(n_3383),
.Y(n_3615)
);

OAI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3445),
.A2(n_3387),
.B1(n_3410),
.B2(n_3412),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3438),
.B(n_3392),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3465),
.B(n_3403),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3438),
.B(n_3362),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3487),
.B(n_3506),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3525),
.B(n_390),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3512),
.B(n_391),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3502),
.B(n_3529),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3518),
.B(n_392),
.Y(n_3624)
);

OAI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3544),
.A2(n_3418),
.B1(n_3409),
.B2(n_396),
.Y(n_3625)
);

NAND3xp33_ASAP7_75t_L g3626 ( 
.A(n_3486),
.B(n_393),
.C(n_395),
.Y(n_3626)
);

NAND3xp33_ASAP7_75t_L g3627 ( 
.A(n_3560),
.B(n_393),
.C(n_395),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3444),
.B(n_396),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3434),
.B(n_397),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3551),
.Y(n_3630)
);

OAI21xp33_ASAP7_75t_L g3631 ( 
.A1(n_3537),
.A2(n_3574),
.B(n_3495),
.Y(n_3631)
);

AOI221xp5_ASAP7_75t_L g3632 ( 
.A1(n_3556),
.A2(n_3479),
.B1(n_3531),
.B2(n_3557),
.C(n_3559),
.Y(n_3632)
);

NAND2xp33_ASAP7_75t_L g3633 ( 
.A(n_3440),
.B(n_397),
.Y(n_3633)
);

OAI21xp5_ASAP7_75t_SL g3634 ( 
.A1(n_3498),
.A2(n_3566),
.B(n_3427),
.Y(n_3634)
);

NAND3xp33_ASAP7_75t_L g3635 ( 
.A(n_3476),
.B(n_398),
.C(n_399),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3434),
.B(n_399),
.Y(n_3636)
);

OA21x2_ASAP7_75t_L g3637 ( 
.A1(n_3458),
.A2(n_400),
.B(n_402),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3538),
.B(n_403),
.Y(n_3638)
);

NAND3xp33_ASAP7_75t_L g3639 ( 
.A(n_3543),
.B(n_403),
.C(n_404),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3455),
.B(n_3472),
.Y(n_3640)
);

NAND3xp33_ASAP7_75t_L g3641 ( 
.A(n_3480),
.B(n_405),
.C(n_406),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3475),
.B(n_405),
.Y(n_3642)
);

OAI221xp5_ASAP7_75t_L g3643 ( 
.A1(n_3428),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.C(n_410),
.Y(n_3643)
);

AOI221xp5_ASAP7_75t_L g3644 ( 
.A1(n_3565),
.A2(n_408),
.B1(n_412),
.B2(n_414),
.C(n_415),
.Y(n_3644)
);

NOR3xp33_ASAP7_75t_L g3645 ( 
.A(n_3552),
.B(n_412),
.C(n_415),
.Y(n_3645)
);

AND2x2_ASAP7_75t_SL g3646 ( 
.A(n_3460),
.B(n_3466),
.Y(n_3646)
);

NAND3xp33_ASAP7_75t_L g3647 ( 
.A(n_3565),
.B(n_416),
.C(n_417),
.Y(n_3647)
);

NAND3xp33_ASAP7_75t_L g3648 ( 
.A(n_3505),
.B(n_416),
.C(n_417),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3470),
.B(n_420),
.Y(n_3649)
);

OAI221xp5_ASAP7_75t_L g3650 ( 
.A1(n_3575),
.A2(n_421),
.B1(n_422),
.B2(n_424),
.C(n_425),
.Y(n_3650)
);

AND2x4_ASAP7_75t_L g3651 ( 
.A(n_3467),
.B(n_422),
.Y(n_3651)
);

HB1xp67_ASAP7_75t_L g3652 ( 
.A(n_3589),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3634),
.A2(n_3442),
.B1(n_3564),
.B2(n_3443),
.Y(n_3653)
);

NAND3xp33_ASAP7_75t_L g3654 ( 
.A(n_3577),
.B(n_3555),
.C(n_3460),
.Y(n_3654)
);

AOI22xp33_ASAP7_75t_L g3655 ( 
.A1(n_3602),
.A2(n_3433),
.B1(n_3424),
.B2(n_3485),
.Y(n_3655)
);

BUFx2_ASAP7_75t_L g3656 ( 
.A(n_3580),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3594),
.B(n_3446),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_L g3658 ( 
.A1(n_3614),
.A2(n_3533),
.B1(n_3568),
.B2(n_3576),
.Y(n_3658)
);

AO221x1_ASAP7_75t_L g3659 ( 
.A1(n_3583),
.A2(n_3463),
.B1(n_3481),
.B2(n_3461),
.C(n_3546),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3630),
.B(n_3477),
.Y(n_3660)
);

NOR3xp33_ASAP7_75t_L g3661 ( 
.A(n_3591),
.B(n_3524),
.C(n_3508),
.Y(n_3661)
);

OR2x2_ASAP7_75t_L g3662 ( 
.A(n_3586),
.B(n_3446),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3584),
.B(n_3469),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3587),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3588),
.B(n_3446),
.Y(n_3665)
);

OR2x2_ASAP7_75t_L g3666 ( 
.A(n_3582),
.B(n_3541),
.Y(n_3666)
);

NOR3xp33_ASAP7_75t_L g3667 ( 
.A(n_3631),
.B(n_3627),
.C(n_3650),
.Y(n_3667)
);

NAND3xp33_ASAP7_75t_L g3668 ( 
.A(n_3579),
.B(n_3550),
.C(n_3536),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3593),
.B(n_3474),
.Y(n_3669)
);

OAI22xp5_ASAP7_75t_L g3670 ( 
.A1(n_3627),
.A2(n_3451),
.B1(n_3448),
.B2(n_3540),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3590),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3592),
.Y(n_3672)
);

AOI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3632),
.A2(n_3530),
.B1(n_3547),
.B2(n_3454),
.Y(n_3673)
);

AOI22xp33_ASAP7_75t_L g3674 ( 
.A1(n_3600),
.A2(n_3510),
.B1(n_3567),
.B2(n_3536),
.Y(n_3674)
);

INVx1_ASAP7_75t_SL g3675 ( 
.A(n_3581),
.Y(n_3675)
);

OR2x2_ASAP7_75t_L g3676 ( 
.A(n_3599),
.B(n_3573),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3596),
.B(n_3488),
.Y(n_3677)
);

NAND3xp33_ASAP7_75t_L g3678 ( 
.A(n_3605),
.B(n_3550),
.C(n_3572),
.Y(n_3678)
);

AOI22xp33_ASAP7_75t_SL g3679 ( 
.A1(n_3595),
.A2(n_3453),
.B1(n_3516),
.B2(n_3484),
.Y(n_3679)
);

NAND2xp33_ASAP7_75t_R g3680 ( 
.A(n_3605),
.B(n_3516),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_SL g3681 ( 
.A(n_3646),
.B(n_3595),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3598),
.Y(n_3682)
);

OAI221xp5_ASAP7_75t_L g3683 ( 
.A1(n_3606),
.A2(n_3511),
.B1(n_3540),
.B2(n_3526),
.C(n_3534),
.Y(n_3683)
);

NAND3xp33_ASAP7_75t_L g3684 ( 
.A(n_3585),
.B(n_3572),
.C(n_3553),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3623),
.B(n_3459),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3620),
.B(n_3464),
.Y(n_3686)
);

OAI211xp5_ASAP7_75t_SL g3687 ( 
.A1(n_3601),
.A2(n_3514),
.B(n_3501),
.C(n_3497),
.Y(n_3687)
);

NOR3xp33_ASAP7_75t_L g3688 ( 
.A(n_3643),
.B(n_3515),
.C(n_3499),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3612),
.B(n_3611),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3615),
.B(n_3523),
.Y(n_3690)
);

OR2x2_ASAP7_75t_L g3691 ( 
.A(n_3608),
.B(n_3482),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3640),
.B(n_3483),
.Y(n_3692)
);

AO21x2_ASAP7_75t_L g3693 ( 
.A1(n_3621),
.A2(n_3439),
.B(n_3516),
.Y(n_3693)
);

NAND3xp33_ASAP7_75t_L g3694 ( 
.A(n_3645),
.B(n_3549),
.C(n_3520),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3617),
.B(n_3468),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_SL g3696 ( 
.A(n_3651),
.B(n_3493),
.Y(n_3696)
);

AND2x2_ASAP7_75t_L g3697 ( 
.A(n_3603),
.B(n_3489),
.Y(n_3697)
);

OR2x2_ASAP7_75t_L g3698 ( 
.A(n_3604),
.B(n_3489),
.Y(n_3698)
);

NAND4xp75_ASAP7_75t_L g3699 ( 
.A(n_3637),
.B(n_3504),
.C(n_3496),
.D(n_3513),
.Y(n_3699)
);

AND2x2_ASAP7_75t_SL g3700 ( 
.A(n_3633),
.B(n_3491),
.Y(n_3700)
);

OAI211xp5_ASAP7_75t_L g3701 ( 
.A1(n_3578),
.A2(n_3532),
.B(n_3527),
.C(n_3562),
.Y(n_3701)
);

NOR3xp33_ASAP7_75t_L g3702 ( 
.A(n_3647),
.B(n_3517),
.C(n_3558),
.Y(n_3702)
);

OR2x2_ASAP7_75t_L g3703 ( 
.A(n_3609),
.B(n_424),
.Y(n_3703)
);

XOR2x2_ASAP7_75t_L g3704 ( 
.A(n_3607),
.B(n_425),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3618),
.B(n_3521),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3651),
.B(n_3563),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3619),
.B(n_3522),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3610),
.B(n_3570),
.Y(n_3708)
);

NAND4xp75_ASAP7_75t_L g3709 ( 
.A(n_3637),
.B(n_426),
.C(n_427),
.D(n_429),
.Y(n_3709)
);

INVx2_ASAP7_75t_SL g3710 ( 
.A(n_3656),
.Y(n_3710)
);

NAND4xp75_ASAP7_75t_L g3711 ( 
.A(n_3681),
.B(n_3642),
.C(n_3644),
.D(n_3629),
.Y(n_3711)
);

INVx2_ASAP7_75t_SL g3712 ( 
.A(n_3652),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3662),
.Y(n_3713)
);

INVxp67_ASAP7_75t_L g3714 ( 
.A(n_3685),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_SL g3715 ( 
.A(n_3675),
.B(n_3625),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3682),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3686),
.B(n_3597),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3653),
.A2(n_3647),
.B1(n_3635),
.B2(n_3641),
.Y(n_3718)
);

XNOR2xp5_ASAP7_75t_L g3719 ( 
.A(n_3704),
.B(n_3613),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3689),
.B(n_3616),
.Y(n_3720)
);

NAND4xp75_ASAP7_75t_SL g3721 ( 
.A(n_3659),
.B(n_3706),
.C(n_3680),
.D(n_3679),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3689),
.B(n_3636),
.Y(n_3722)
);

INVx5_ASAP7_75t_L g3723 ( 
.A(n_3709),
.Y(n_3723)
);

OAI22xp5_ASAP7_75t_L g3724 ( 
.A1(n_3675),
.A2(n_3635),
.B1(n_3641),
.B2(n_3648),
.Y(n_3724)
);

INVx2_ASAP7_75t_SL g3725 ( 
.A(n_3672),
.Y(n_3725)
);

INVx2_ASAP7_75t_SL g3726 ( 
.A(n_3664),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3669),
.B(n_3663),
.Y(n_3727)
);

INVxp67_ASAP7_75t_SL g3728 ( 
.A(n_3665),
.Y(n_3728)
);

NAND4xp75_ASAP7_75t_L g3729 ( 
.A(n_3700),
.B(n_3622),
.C(n_3624),
.D(n_3628),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3671),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3666),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3661),
.A2(n_3648),
.B1(n_3639),
.B2(n_3649),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3677),
.Y(n_3733)
);

INVx2_ASAP7_75t_SL g3734 ( 
.A(n_3703),
.Y(n_3734)
);

INVx1_ASAP7_75t_SL g3735 ( 
.A(n_3676),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3665),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3697),
.B(n_3638),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3691),
.Y(n_3738)
);

OR2x2_ASAP7_75t_L g3739 ( 
.A(n_3657),
.B(n_3626),
.Y(n_3739)
);

NAND3xp33_ASAP7_75t_L g3740 ( 
.A(n_3667),
.B(n_426),
.C(n_427),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3698),
.B(n_429),
.Y(n_3741)
);

AOI22xp5_ASAP7_75t_L g3742 ( 
.A1(n_3654),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_3742)
);

AND2x4_ASAP7_75t_L g3743 ( 
.A(n_3693),
.B(n_3692),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3695),
.B(n_432),
.Y(n_3744)
);

OR2x2_ASAP7_75t_L g3745 ( 
.A(n_3657),
.B(n_433),
.Y(n_3745)
);

XNOR2x2_ASAP7_75t_L g3746 ( 
.A(n_3678),
.B(n_433),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3677),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3690),
.Y(n_3748)
);

XNOR2xp5_ASAP7_75t_L g3749 ( 
.A(n_3655),
.B(n_435),
.Y(n_3749)
);

INVx4_ASAP7_75t_L g3750 ( 
.A(n_3693),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3660),
.Y(n_3751)
);

NAND4xp75_ASAP7_75t_L g3752 ( 
.A(n_3696),
.B(n_436),
.C(n_437),
.D(n_440),
.Y(n_3752)
);

AOI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_3670),
.A2(n_437),
.B1(n_440),
.B2(n_441),
.Y(n_3753)
);

XNOR2xp5_ASAP7_75t_L g3754 ( 
.A(n_3707),
.B(n_441),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3690),
.B(n_442),
.Y(n_3755)
);

NAND4xp75_ASAP7_75t_L g3756 ( 
.A(n_3708),
.B(n_442),
.C(n_443),
.D(n_444),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3705),
.B(n_445),
.Y(n_3757)
);

AND2x4_ASAP7_75t_L g3758 ( 
.A(n_3708),
.B(n_446),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3668),
.B(n_448),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3670),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3684),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3738),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3760),
.A2(n_3715),
.B1(n_3718),
.B2(n_3761),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3712),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3760),
.B(n_3674),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3733),
.Y(n_3766)
);

INVxp67_ASAP7_75t_L g3767 ( 
.A(n_3759),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3719),
.B(n_3687),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3747),
.Y(n_3769)
);

XOR2x2_ASAP7_75t_L g3770 ( 
.A(n_3721),
.B(n_3699),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3726),
.Y(n_3771)
);

INVxp67_ASAP7_75t_L g3772 ( 
.A(n_3739),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3730),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3725),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3713),
.Y(n_3775)
);

INVx2_ASAP7_75t_SL g3776 ( 
.A(n_3710),
.Y(n_3776)
);

XOR2x2_ASAP7_75t_L g3777 ( 
.A(n_3754),
.B(n_3673),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3748),
.B(n_3688),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3716),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3713),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3736),
.Y(n_3781)
);

XNOR2x1_ASAP7_75t_L g3782 ( 
.A(n_3749),
.B(n_3694),
.Y(n_3782)
);

CKINVDCx8_ASAP7_75t_R g3783 ( 
.A(n_3723),
.Y(n_3783)
);

XNOR2x2_ASAP7_75t_L g3784 ( 
.A(n_3746),
.B(n_3683),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3736),
.Y(n_3785)
);

OA22x2_ASAP7_75t_L g3786 ( 
.A1(n_3743),
.A2(n_3701),
.B1(n_3658),
.B2(n_3702),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3731),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3748),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3751),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3728),
.B(n_448),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3727),
.B(n_450),
.Y(n_3791)
);

AOI22x1_ASAP7_75t_L g3792 ( 
.A1(n_3784),
.A2(n_3758),
.B1(n_3750),
.B2(n_3745),
.Y(n_3792)
);

INVx2_ASAP7_75t_SL g3793 ( 
.A(n_3774),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3789),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3762),
.Y(n_3795)
);

AOI22x1_ASAP7_75t_L g3796 ( 
.A1(n_3786),
.A2(n_3758),
.B1(n_3750),
.B2(n_3741),
.Y(n_3796)
);

OA22x2_ASAP7_75t_L g3797 ( 
.A1(n_3763),
.A2(n_3743),
.B1(n_3732),
.B2(n_3717),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3773),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3766),
.Y(n_3799)
);

OA22x2_ASAP7_75t_L g3800 ( 
.A1(n_3765),
.A2(n_3714),
.B1(n_3720),
.B2(n_3753),
.Y(n_3800)
);

INVx1_ASAP7_75t_SL g3801 ( 
.A(n_3791),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3779),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3769),
.Y(n_3803)
);

AOI22x1_ASAP7_75t_L g3804 ( 
.A1(n_3786),
.A2(n_3755),
.B1(n_3734),
.B2(n_3735),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3787),
.Y(n_3805)
);

OA22x2_ASAP7_75t_L g3806 ( 
.A1(n_3765),
.A2(n_3724),
.B1(n_3742),
.B2(n_3737),
.Y(n_3806)
);

OA22x2_ASAP7_75t_L g3807 ( 
.A1(n_3772),
.A2(n_3757),
.B1(n_3744),
.B2(n_3722),
.Y(n_3807)
);

INVx1_ASAP7_75t_SL g3808 ( 
.A(n_3776),
.Y(n_3808)
);

HB1xp67_ASAP7_75t_L g3809 ( 
.A(n_3772),
.Y(n_3809)
);

XOR2x2_ASAP7_75t_L g3810 ( 
.A(n_3770),
.B(n_3729),
.Y(n_3810)
);

INVx1_ASAP7_75t_SL g3811 ( 
.A(n_3790),
.Y(n_3811)
);

NAND2xp33_ASAP7_75t_L g3812 ( 
.A(n_3771),
.B(n_3723),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3785),
.Y(n_3813)
);

INVxp67_ASAP7_75t_L g3814 ( 
.A(n_3790),
.Y(n_3814)
);

XOR2x2_ASAP7_75t_L g3815 ( 
.A(n_3777),
.B(n_3782),
.Y(n_3815)
);

OAI22x1_ASAP7_75t_L g3816 ( 
.A1(n_3768),
.A2(n_3723),
.B1(n_3740),
.B2(n_3711),
.Y(n_3816)
);

XOR2x2_ASAP7_75t_L g3817 ( 
.A(n_3768),
.B(n_3752),
.Y(n_3817)
);

INVx1_ASAP7_75t_SL g3818 ( 
.A(n_3764),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3767),
.B(n_3756),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3788),
.Y(n_3820)
);

AOI22x1_ASAP7_75t_L g3821 ( 
.A1(n_3783),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.Y(n_3821)
);

OA22x2_ASAP7_75t_L g3822 ( 
.A1(n_3767),
.A2(n_451),
.B1(n_452),
.B2(n_454),
.Y(n_3822)
);

OA22x2_ASAP7_75t_L g3823 ( 
.A1(n_3778),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3778),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3809),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3794),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3799),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3803),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3798),
.Y(n_3829)
);

NOR2x1_ASAP7_75t_L g3830 ( 
.A(n_3812),
.B(n_3785),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3805),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3818),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3820),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3795),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3795),
.Y(n_3835)
);

INVxp67_ASAP7_75t_SL g3836 ( 
.A(n_3823),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3802),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3808),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3824),
.Y(n_3839)
);

INVx1_ASAP7_75t_SL g3840 ( 
.A(n_3822),
.Y(n_3840)
);

BUFx3_ASAP7_75t_L g3841 ( 
.A(n_3793),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3814),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3811),
.Y(n_3843)
);

INVx1_ASAP7_75t_SL g3844 ( 
.A(n_3817),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3813),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3792),
.Y(n_3846)
);

OAI322xp33_ASAP7_75t_L g3847 ( 
.A1(n_3797),
.A2(n_3780),
.A3(n_3775),
.B1(n_3781),
.B2(n_462),
.C1(n_463),
.C2(n_464),
.Y(n_3847)
);

INVxp67_ASAP7_75t_L g3848 ( 
.A(n_3816),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3792),
.Y(n_3849)
);

AOI221xp5_ASAP7_75t_L g3850 ( 
.A1(n_3847),
.A2(n_3819),
.B1(n_3801),
.B2(n_3815),
.C(n_3806),
.Y(n_3850)
);

NAND4xp75_ASAP7_75t_L g3851 ( 
.A(n_3846),
.B(n_3804),
.C(n_3796),
.D(n_3810),
.Y(n_3851)
);

AOI22xp5_ASAP7_75t_L g3852 ( 
.A1(n_3848),
.A2(n_3800),
.B1(n_3807),
.B2(n_3796),
.Y(n_3852)
);

NAND4xp75_ASAP7_75t_L g3853 ( 
.A(n_3849),
.B(n_3804),
.C(n_3821),
.D(n_461),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3832),
.Y(n_3854)
);

INVxp67_ASAP7_75t_L g3855 ( 
.A(n_3841),
.Y(n_3855)
);

NAND4xp75_ASAP7_75t_L g3856 ( 
.A(n_3838),
.B(n_3821),
.C(n_460),
.D(n_461),
.Y(n_3856)
);

INVxp67_ASAP7_75t_L g3857 ( 
.A(n_3836),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3848),
.A2(n_455),
.B1(n_460),
.B2(n_462),
.Y(n_3858)
);

INVx3_ASAP7_75t_L g3859 ( 
.A(n_3837),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3825),
.Y(n_3860)
);

NAND4xp75_ASAP7_75t_L g3861 ( 
.A(n_3843),
.B(n_463),
.C(n_464),
.D(n_465),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3842),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3845),
.Y(n_3863)
);

AOI22xp5_ASAP7_75t_L g3864 ( 
.A1(n_3840),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_3864)
);

AOI221xp5_ASAP7_75t_L g3865 ( 
.A1(n_3844),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.C(n_469),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3839),
.Y(n_3866)
);

OAI22xp5_ASAP7_75t_L g3867 ( 
.A1(n_3840),
.A2(n_3844),
.B1(n_3830),
.B2(n_3829),
.Y(n_3867)
);

AOI22x1_ASAP7_75t_L g3868 ( 
.A1(n_3826),
.A2(n_470),
.B1(n_471),
.B2(n_472),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3854),
.Y(n_3869)
);

OAI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_3851),
.A2(n_3831),
.B1(n_3828),
.B2(n_3827),
.Y(n_3870)
);

HB1xp67_ASAP7_75t_L g3871 ( 
.A(n_3857),
.Y(n_3871)
);

BUFx2_ASAP7_75t_L g3872 ( 
.A(n_3855),
.Y(n_3872)
);

AO22x2_ASAP7_75t_L g3873 ( 
.A1(n_3867),
.A2(n_3833),
.B1(n_3835),
.B2(n_3834),
.Y(n_3873)
);

O2A1O1Ixp33_ASAP7_75t_SL g3874 ( 
.A1(n_3850),
.A2(n_470),
.B(n_471),
.C(n_472),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3860),
.Y(n_3875)
);

AOI22xp5_ASAP7_75t_L g3876 ( 
.A1(n_3852),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.Y(n_3876)
);

AOI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_3853),
.A2(n_475),
.B1(n_477),
.B2(n_479),
.Y(n_3877)
);

NOR4xp25_ASAP7_75t_L g3878 ( 
.A(n_3862),
.B(n_477),
.C(n_479),
.D(n_480),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3863),
.Y(n_3879)
);

AOI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3864),
.A2(n_480),
.B1(n_481),
.B2(n_483),
.Y(n_3880)
);

AOI22xp5_ASAP7_75t_L g3881 ( 
.A1(n_3856),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_3859),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3859),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_3883)
);

OAI22xp5_ASAP7_75t_L g3884 ( 
.A1(n_3866),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_3884)
);

AOI22xp33_ASAP7_75t_SL g3885 ( 
.A1(n_3868),
.A2(n_488),
.B1(n_489),
.B2(n_490),
.Y(n_3885)
);

AO22x2_ASAP7_75t_L g3886 ( 
.A1(n_3870),
.A2(n_3861),
.B1(n_3865),
.B2(n_3858),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3872),
.Y(n_3887)
);

AO22x1_ASAP7_75t_L g3888 ( 
.A1(n_3871),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_3888)
);

AOI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3874),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3877),
.A2(n_492),
.B1(n_494),
.B2(n_495),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3879),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3883),
.Y(n_3892)
);

NOR3xp33_ASAP7_75t_L g3893 ( 
.A(n_3884),
.B(n_495),
.C(n_496),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3882),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3869),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3875),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3876),
.A2(n_498),
.B1(n_499),
.B2(n_501),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3887),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3894),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3891),
.Y(n_3900)
);

AOI22xp33_ASAP7_75t_L g3901 ( 
.A1(n_3892),
.A2(n_3873),
.B1(n_3885),
.B2(n_3881),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3888),
.Y(n_3902)
);

AOI22xp33_ASAP7_75t_L g3903 ( 
.A1(n_3886),
.A2(n_3873),
.B1(n_3880),
.B2(n_3878),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3895),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3896),
.Y(n_3905)
);

OR2x2_ASAP7_75t_L g3906 ( 
.A(n_3889),
.B(n_502),
.Y(n_3906)
);

AOI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3902),
.A2(n_3901),
.B1(n_3898),
.B2(n_3903),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3899),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3906),
.Y(n_3909)
);

NOR3xp33_ASAP7_75t_L g3910 ( 
.A(n_3900),
.B(n_3897),
.C(n_3893),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3905),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3907),
.A2(n_3901),
.B1(n_3890),
.B2(n_3904),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3908),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3911),
.Y(n_3914)
);

BUFx2_ASAP7_75t_L g3915 ( 
.A(n_3909),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3910),
.Y(n_3916)
);

AO22x2_ASAP7_75t_L g3917 ( 
.A1(n_3913),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.Y(n_3917)
);

OAI22xp5_ASAP7_75t_L g3918 ( 
.A1(n_3912),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_3918)
);

CKINVDCx20_ASAP7_75t_R g3919 ( 
.A(n_3915),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3914),
.A2(n_506),
.B1(n_507),
.B2(n_508),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3917),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3919),
.Y(n_3922)
);

O2A1O1Ixp33_ASAP7_75t_L g3923 ( 
.A1(n_3922),
.A2(n_3918),
.B(n_3916),
.C(n_3920),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3923),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3924),
.A2(n_3921),
.B1(n_509),
.B2(n_511),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3925),
.Y(n_3926)
);

AOI221xp5_ASAP7_75t_L g3927 ( 
.A1(n_3926),
.A2(n_508),
.B1(n_509),
.B2(n_512),
.C(n_513),
.Y(n_3927)
);

AOI211xp5_ASAP7_75t_L g3928 ( 
.A1(n_3927),
.A2(n_513),
.B(n_514),
.C(n_515),
.Y(n_3928)
);


endmodule