module fake_netlist_1_7981_n_1281 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_191, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1281);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_191;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1281;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_158), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_217), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_26), .B(n_186), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_162), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_137), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_174), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_108), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_244), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_212), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_192), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_301), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_185), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_156), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_305), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_254), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_98), .Y(n_323) );
CKINVDCx16_ASAP7_75t_R g324 ( .A(n_278), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_290), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_255), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_165), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_148), .Y(n_328) );
INVxp33_ASAP7_75t_L g329 ( .A(n_222), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_257), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_184), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_90), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_24), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_102), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_51), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_250), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_198), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_50), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_256), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_161), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_123), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_200), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_34), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_145), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_297), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_269), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_41), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_202), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_159), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_204), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_218), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_47), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_271), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_211), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_136), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_169), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_49), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_120), .Y(n_362) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_231), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_173), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_232), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_201), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_191), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_229), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_273), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_170), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_118), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_168), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_79), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_134), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_50), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_249), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_240), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_69), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_251), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_138), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_209), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_166), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_282), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_112), .Y(n_385) );
BUFx2_ASAP7_75t_R g386 ( .A(n_261), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_90), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_41), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_141), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_40), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_7), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_114), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_139), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_16), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_233), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_296), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_106), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_235), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_276), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_289), .Y(n_400) );
INVxp33_ASAP7_75t_SL g401 ( .A(n_243), .Y(n_401) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_277), .B(n_28), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_179), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_221), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_143), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_283), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_152), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_81), .Y(n_408) );
BUFx10_ASAP7_75t_L g409 ( .A(n_160), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_10), .Y(n_410) );
XNOR2xp5_ASAP7_75t_L g411 ( .A(n_225), .B(n_44), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_121), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_144), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_194), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_268), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_171), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_27), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_247), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_85), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_196), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_195), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_87), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_219), .Y(n_423) );
INVxp33_ASAP7_75t_SL g424 ( .A(n_103), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_234), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_31), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_11), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_53), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_180), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_286), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_26), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_61), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_31), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_270), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_127), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_285), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_199), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_288), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_237), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_150), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_2), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_172), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_187), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_77), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_154), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_163), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_15), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_164), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_298), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_197), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_293), .Y(n_451) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_284), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_20), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_14), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_213), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_181), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_259), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_280), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_167), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_294), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_86), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_14), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_149), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_274), .Y(n_464) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_116), .B(n_275), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_279), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_104), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_258), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_123), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_287), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_193), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_97), .B(n_239), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_108), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_265), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_42), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_224), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_248), .Y(n_477) );
BUFx5_ASAP7_75t_L g478 ( .A(n_292), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_245), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_188), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_135), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_48), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_132), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_133), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_359), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_387), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_359), .B(n_0), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_387), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_409), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_359), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_478), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_410), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_478), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_478), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_315), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_410), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_329), .B(n_0), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_326), .B(n_1), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_478), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_409), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_462), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_478), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_462), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_398), .B(n_1), .Y(n_504) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_312), .A2(n_140), .B(n_131), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_468), .B(n_2), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_324), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_308), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_315), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_313), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_432), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_310), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_405), .B(n_3), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_338), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_478), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_334), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_478), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_379), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_424), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_314), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_363), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_457), .B(n_6), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_316), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_318), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_330), .B(n_7), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_424), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_409), .Y(n_527) );
NAND2xp33_ASAP7_75t_SL g528 ( .A(n_329), .B(n_8), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_519), .A2(n_397), .B1(n_441), .B2(n_386), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_491), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_508), .B(n_455), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_489), .B(n_479), .Y(n_532) );
INVx4_ASAP7_75t_L g533 ( .A(n_487), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_508), .B(n_312), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_516), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_489), .B(n_418), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_514), .B(n_425), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_491), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_487), .Y(n_539) );
OR2x6_ASAP7_75t_L g540 ( .A(n_497), .B(n_309), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_512), .B(n_319), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_489), .B(n_333), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_510), .Y(n_544) );
BUFx8_ASAP7_75t_SL g545 ( .A(n_507), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_491), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_516), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_510), .B(n_427), .Y(n_548) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_522), .A2(n_321), .B(n_320), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_518), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_489), .B(n_452), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_512), .A2(n_339), .B1(n_347), .B2(n_345), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_493), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_516), .Y(n_556) );
BUFx10_ASAP7_75t_L g557 ( .A(n_525), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_494), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_494), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_516), .Y(n_560) );
NOR2xp33_ASAP7_75t_SL g561 ( .A(n_497), .B(n_332), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_494), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_516), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_499), .Y(n_565) );
BUFx4f_ASAP7_75t_L g566 ( .A(n_525), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_485), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_531), .B(n_514), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_531), .B(n_500), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_550), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_561), .A2(n_526), .B1(n_519), .B2(n_518), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_550), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_566), .B(n_525), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_532), .B(n_500), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_542), .B(n_500), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_533), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_542), .B(n_527), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_542), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_550), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_542), .B(n_527), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_566), .A2(n_505), .B(n_527), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_536), .B(n_527), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_564), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_567), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_544), .B(n_521), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_552), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_567), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_529), .B(n_506), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_537), .B(n_506), .Y(n_591) );
AOI221x1_ASAP7_75t_L g592 ( .A1(n_543), .A2(n_522), .B1(n_524), .B2(n_523), .C(n_520), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_553), .B(n_520), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_533), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_567), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_537), .B(n_498), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_552), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_548), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_540), .A2(n_528), .B1(n_524), .B2(n_523), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_540), .B(n_498), .Y(n_602) );
BUFx3_ASAP7_75t_L g603 ( .A(n_557), .Y(n_603) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_529), .B(n_504), .Y(n_604) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_543), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_540), .A2(n_504), .B1(n_509), .B2(n_495), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_540), .A2(n_495), .B1(n_509), .B2(n_513), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_540), .B(n_495), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_543), .Y(n_609) );
O2A1O1Ixp5_ASAP7_75t_L g610 ( .A1(n_534), .A2(n_490), .B(n_503), .C(n_501), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_539), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_561), .A2(n_526), .B1(n_511), .B2(n_441), .Y(n_612) );
BUFx12f_ASAP7_75t_L g613 ( .A(n_548), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_549), .B(n_501), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_549), .B(n_503), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_549), .A2(n_505), .B(n_517), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_534), .B(n_401), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_541), .B(n_307), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_545), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_530), .B(n_502), .Y(n_620) );
NOR2x1p5_ASAP7_75t_L g621 ( .A(n_541), .B(n_376), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_530), .B(n_511), .C(n_388), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_538), .B(n_502), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_546), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_554), .B(n_401), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_554), .B(n_486), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_551), .Y(n_627) );
HB1xp67_ASAP7_75t_SL g628 ( .A(n_551), .Y(n_628) );
INVx4_ASAP7_75t_L g629 ( .A(n_555), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_555), .B(n_335), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_558), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_559), .B(n_486), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_559), .A2(n_397), .B1(n_352), .B2(n_353), .Y(n_633) );
INVx4_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_565), .B(n_502), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_535), .A2(n_505), .B(n_515), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_535), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_603), .B(n_327), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_603), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_600), .B(n_341), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_628), .A2(n_358), .B1(n_378), .B2(n_353), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_631), .A2(n_378), .B1(n_383), .B2(n_358), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_598), .B(n_328), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_582), .A2(n_505), .B(n_515), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_571), .A2(n_361), .B(n_362), .C(n_351), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_621), .B(n_383), .Y(n_646) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_629), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_588), .B(n_389), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_594), .A2(n_490), .B(n_517), .C(n_374), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_573), .A2(n_505), .B(n_517), .Y(n_650) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_597), .B(n_389), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_594), .A2(n_385), .B(n_390), .C(n_372), .Y(n_652) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_629), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_616), .A2(n_395), .B(n_322), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_629), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_577), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_631), .A2(n_439), .B1(n_481), .B2(n_471), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_568), .A2(n_392), .B(n_391), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_602), .A2(n_471), .B1(n_481), .B2(n_439), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_617), .A2(n_412), .B(n_417), .C(n_394), .Y(n_660) );
INVx3_ASAP7_75t_SL g661 ( .A(n_587), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_617), .B(n_336), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_580), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_569), .B(n_342), .Y(n_664) );
INVx11_ASAP7_75t_L g665 ( .A(n_613), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_591), .B(n_356), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_627), .A2(n_411), .B1(n_463), .B2(n_393), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_612), .A2(n_433), .B(n_447), .C(n_428), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_633), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_590), .B(n_408), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_625), .A2(n_422), .B1(n_426), .B2(n_419), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_604), .B(n_435), .Y(n_673) );
INVx3_ASAP7_75t_L g674 ( .A(n_634), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_630), .B(n_461), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_618), .B(n_444), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_622), .A2(n_475), .B(n_467), .C(n_488), .Y(n_677) );
AOI21x1_ASAP7_75t_L g678 ( .A1(n_636), .A2(n_563), .B(n_547), .Y(n_678) );
INVx4_ASAP7_75t_L g679 ( .A(n_634), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_634), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_601), .A2(n_454), .B1(n_469), .B2(n_453), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_606), .A2(n_483), .B1(n_466), .B2(n_482), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_626), .A2(n_323), .B1(n_431), .B2(n_473), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_632), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_599), .Y(n_685) );
BUFx12f_ASAP7_75t_L g686 ( .A(n_619), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_610), .A2(n_465), .B(n_402), .C(n_492), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_614), .A2(n_496), .B(n_337), .C(n_343), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_632), .B(n_496), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_583), .B(n_483), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_611), .A2(n_344), .B(n_331), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_615), .A2(n_348), .B(n_346), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_575), .B(n_323), .Y(n_693) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_607), .A2(n_472), .B1(n_431), .B2(n_323), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_583), .B(n_317), .Y(n_695) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_575), .Y(n_696) );
AO21x1_ASAP7_75t_L g697 ( .A1(n_574), .A2(n_357), .B(n_350), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_608), .B(n_323), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_599), .Y(n_699) );
AOI22x1_ASAP7_75t_L g700 ( .A1(n_609), .A2(n_325), .B1(n_377), .B2(n_319), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_609), .A2(n_366), .B(n_365), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_624), .A2(n_367), .B(n_369), .C(n_368), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_605), .A2(n_371), .B(n_370), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_576), .B(n_380), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_620), .A2(n_382), .B(n_381), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_593), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_623), .A2(n_399), .B(n_396), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_595), .B(n_404), .Y(n_708) );
AOI21x1_ASAP7_75t_L g709 ( .A1(n_623), .A2(n_415), .B(n_413), .Y(n_709) );
CKINVDCx11_ASAP7_75t_R g710 ( .A(n_570), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_635), .A2(n_420), .B(n_416), .Y(n_711) );
AO32x1_ASAP7_75t_L g712 ( .A1(n_592), .A2(n_438), .A3(n_440), .B1(n_437), .B2(n_434), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_635), .A2(n_445), .B(n_443), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g714 ( .A1(n_581), .A2(n_451), .B(n_450), .Y(n_714) );
NOR2xp33_ASAP7_75t_R g715 ( .A(n_595), .B(n_311), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_584), .Y(n_716) );
NOR2xp67_ASAP7_75t_R g717 ( .A(n_585), .B(n_430), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_586), .A2(n_579), .B(n_572), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_572), .A2(n_470), .B(n_459), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_579), .A2(n_477), .B(n_484), .C(n_474), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_589), .Y(n_721) );
BUFx4f_ASAP7_75t_L g722 ( .A(n_596), .Y(n_722) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_637), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_582), .A2(n_460), .B(n_458), .Y(n_724) );
NOR2xp67_ASAP7_75t_L g725 ( .A(n_619), .B(n_9), .Y(n_725) );
CKINVDCx10_ASAP7_75t_R g726 ( .A(n_619), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_568), .B(n_349), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_578), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_603), .B(n_354), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_629), .Y(n_730) );
AO21x1_ASAP7_75t_L g731 ( .A1(n_582), .A2(n_442), .B(n_334), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_629), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_568), .B(n_355), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_621), .B(n_431), .Y(n_734) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_571), .A2(n_421), .B(n_464), .C(n_340), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_SL g736 ( .A1(n_614), .A2(n_146), .B(n_147), .C(n_142), .Y(n_736) );
AOI33xp33_ASAP7_75t_L g737 ( .A1(n_571), .A2(n_431), .A3(n_12), .B1(n_13), .B2(n_15), .B3(n_16), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_568), .B(n_360), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_SL g739 ( .A1(n_617), .A2(n_364), .B(n_375), .C(n_373), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g740 ( .A1(n_594), .A2(n_442), .B(n_334), .C(n_384), .Y(n_740) );
OAI21x1_ASAP7_75t_L g741 ( .A1(n_636), .A2(n_560), .B(n_556), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_603), .B(n_400), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g743 ( .A(n_613), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_628), .A2(n_403), .B1(n_407), .B2(n_406), .Y(n_744) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_639), .Y(n_745) );
NOR4xp25_ASAP7_75t_L g746 ( .A(n_737), .B(n_13), .C(n_11), .D(n_12), .Y(n_746) );
O2A1O1Ixp33_ASAP7_75t_L g747 ( .A1(n_660), .A2(n_19), .B(n_17), .C(n_18), .Y(n_747) );
AOI221x1_ASAP7_75t_L g748 ( .A1(n_644), .A2(n_442), .B1(n_334), .B2(n_560), .C(n_556), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_648), .B(n_414), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_650), .A2(n_429), .B(n_423), .Y(n_750) );
AOI21x1_ASAP7_75t_L g751 ( .A1(n_678), .A2(n_442), .B(n_556), .Y(n_751) );
OAI21x1_ASAP7_75t_L g752 ( .A1(n_741), .A2(n_560), .B(n_556), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_654), .A2(n_446), .B(n_436), .Y(n_753) );
INVx3_ASAP7_75t_SL g754 ( .A(n_743), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_688), .A2(n_19), .B(n_17), .C(n_18), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_693), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g757 ( .A1(n_735), .A2(n_449), .B(n_456), .C(n_448), .Y(n_757) );
BUFx10_ASAP7_75t_L g758 ( .A(n_640), .Y(n_758) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_642), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_718), .A2(n_480), .B(n_476), .Y(n_760) );
AOI21x1_ASAP7_75t_L g761 ( .A1(n_731), .A2(n_560), .B(n_556), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_689), .A2(n_672), .B1(n_679), .B2(n_657), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_684), .B(n_21), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g764 ( .A1(n_692), .A2(n_153), .B(n_151), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_645), .B(n_22), .Y(n_765) );
AO32x2_ASAP7_75t_L g766 ( .A1(n_694), .A2(n_23), .A3(n_25), .B1(n_27), .B2(n_28), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_661), .B(n_29), .Y(n_767) );
O2A1O1Ixp33_ASAP7_75t_L g768 ( .A1(n_652), .A2(n_32), .B(n_29), .C(n_30), .Y(n_768) );
O2A1O1Ixp33_ASAP7_75t_L g769 ( .A1(n_668), .A2(n_33), .B(n_30), .C(n_32), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_647), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_724), .A2(n_157), .B(n_155), .Y(n_771) );
AO31x2_ASAP7_75t_L g772 ( .A1(n_687), .A2(n_35), .A3(n_33), .B(n_34), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_659), .A2(n_37), .B1(n_35), .B2(n_36), .Y(n_773) );
INVx4_ASAP7_75t_L g774 ( .A(n_665), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_647), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_641), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_677), .A2(n_40), .B(n_38), .C(n_39), .Y(n_777) );
OAI21x1_ASAP7_75t_L g778 ( .A1(n_709), .A2(n_176), .B(n_175), .Y(n_778) );
INVx5_ASAP7_75t_L g779 ( .A(n_653), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_734), .B(n_43), .Y(n_780) );
AO32x2_ASAP7_75t_L g781 ( .A1(n_694), .A2(n_44), .A3(n_45), .B1(n_46), .B2(n_47), .Y(n_781) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_649), .A2(n_178), .B(n_177), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_658), .B(n_46), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_646), .B(n_48), .Y(n_784) );
OAI21x1_ASAP7_75t_L g785 ( .A1(n_700), .A2(n_183), .B(n_182), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_683), .B(n_49), .C(n_51), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_740), .A2(n_190), .B(n_189), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_658), .B(n_52), .Y(n_788) );
BUFx3_ASAP7_75t_L g789 ( .A(n_710), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_653), .B(n_54), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_728), .Y(n_791) );
AO31x2_ASAP7_75t_L g792 ( .A1(n_697), .A2(n_712), .A3(n_719), .B(n_701), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_646), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_696), .B(n_55), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_656), .B(n_55), .Y(n_795) );
AND2x2_ASAP7_75t_SL g796 ( .A(n_722), .B(n_56), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_651), .B(n_57), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_675), .B(n_671), .Y(n_798) );
AO21x2_ASAP7_75t_L g799 ( .A1(n_736), .A2(n_205), .B(n_203), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_663), .B(n_58), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_674), .B(n_58), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_685), .Y(n_802) );
INVx1_ASAP7_75t_SL g803 ( .A(n_715), .Y(n_803) );
AOI21x1_ASAP7_75t_L g804 ( .A1(n_698), .A2(n_207), .B(n_206), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_667), .B(n_59), .Y(n_805) );
AO31x2_ASAP7_75t_L g806 ( .A1(n_712), .A2(n_59), .A3(n_60), .B(n_61), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_716), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_666), .B(n_62), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_703), .A2(n_210), .B(n_208), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_699), .Y(n_810) );
AO21x1_ASAP7_75t_L g811 ( .A1(n_720), .A2(n_215), .B(n_214), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_L g812 ( .A1(n_702), .A2(n_62), .B(n_63), .C(n_64), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_673), .B(n_65), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_691), .A2(n_220), .B(n_216), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_722), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_815) );
INVx3_ASAP7_75t_L g816 ( .A(n_674), .Y(n_816) );
AND2x2_ASAP7_75t_SL g817 ( .A(n_680), .B(n_67), .Y(n_817) );
INVx1_ASAP7_75t_SL g818 ( .A(n_726), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_670), .B(n_68), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_664), .Y(n_820) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_662), .A2(n_69), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_744), .Y(n_822) );
NAND3xp33_ASAP7_75t_SL g823 ( .A(n_681), .B(n_72), .C(n_73), .Y(n_823) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_655), .Y(n_824) );
AO22x2_ASAP7_75t_L g825 ( .A1(n_682), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_643), .Y(n_826) );
O2A1O1Ixp33_ASAP7_75t_L g827 ( .A1(n_676), .A2(n_74), .B(n_75), .C(n_76), .Y(n_827) );
AO31x2_ASAP7_75t_L g828 ( .A1(n_712), .A2(n_76), .A3(n_77), .B(n_78), .Y(n_828) );
AO31x2_ASAP7_75t_L g829 ( .A1(n_705), .A2(n_78), .A3(n_79), .B(n_80), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_727), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_714), .A2(n_82), .B(n_83), .C(n_84), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_733), .B(n_738), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_SL g833 ( .A1(n_739), .A2(n_236), .B(n_303), .C(n_302), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_706), .Y(n_834) );
INVx1_ASAP7_75t_SL g835 ( .A(n_638), .Y(n_835) );
INVxp67_ASAP7_75t_SL g836 ( .A(n_723), .Y(n_836) );
AND2x4_ASAP7_75t_L g837 ( .A(n_730), .B(n_83), .Y(n_837) );
BUFx3_ASAP7_75t_L g838 ( .A(n_732), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_725), .B(n_88), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_729), .Y(n_840) );
AO21x1_ASAP7_75t_L g841 ( .A1(n_721), .A2(n_238), .B(n_295), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_695), .B(n_89), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_690), .A2(n_89), .B1(n_91), .B2(n_92), .Y(n_843) );
AO31x2_ASAP7_75t_L g844 ( .A1(n_707), .A2(n_91), .A3(n_92), .B(n_93), .Y(n_844) );
OR2x2_ASAP7_75t_L g845 ( .A(n_713), .B(n_93), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_721), .Y(n_846) );
AOI21xp33_ASAP7_75t_L g847 ( .A1(n_704), .A2(n_94), .B(n_95), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_708), .B(n_95), .Y(n_848) );
O2A1O1Ixp33_ASAP7_75t_L g849 ( .A1(n_711), .A2(n_96), .B(n_97), .C(n_98), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_742), .A2(n_96), .B1(n_99), .B2(n_100), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_717), .A2(n_242), .B(n_291), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_717), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_660), .B(n_99), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_659), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_660), .B(n_101), .Y(n_855) );
AO31x2_ASAP7_75t_L g856 ( .A1(n_731), .A2(n_103), .A3(n_104), .B(n_105), .Y(n_856) );
INVxp67_ASAP7_75t_L g857 ( .A(n_642), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_689), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g859 ( .A1(n_735), .A2(n_105), .B(n_106), .C(n_107), .Y(n_859) );
INVx8_ASAP7_75t_L g860 ( .A(n_686), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_660), .B(n_109), .Y(n_861) );
INVx3_ASAP7_75t_L g862 ( .A(n_679), .Y(n_862) );
INVx2_ASAP7_75t_SL g863 ( .A(n_665), .Y(n_863) );
AO31x2_ASAP7_75t_L g864 ( .A1(n_731), .A2(n_110), .A3(n_111), .B(n_113), .Y(n_864) );
NOR2xp67_ASAP7_75t_L g865 ( .A(n_642), .B(n_110), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_689), .Y(n_866) );
AO31x2_ASAP7_75t_L g867 ( .A1(n_731), .A2(n_115), .A3(n_116), .B(n_117), .Y(n_867) );
AO22x2_ASAP7_75t_L g868 ( .A1(n_642), .A2(n_117), .B1(n_118), .B2(n_119), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_820), .B(n_119), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_759), .B(n_120), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_754), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g872 ( .A1(n_750), .A2(n_246), .B(n_281), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_858), .B(n_121), .Y(n_873) );
INVx4_ASAP7_75t_SL g874 ( .A(n_789), .Y(n_874) );
NAND2x1p5_ASAP7_75t_L g875 ( .A(n_774), .B(n_122), .Y(n_875) );
AOI21xp33_ASAP7_75t_SL g876 ( .A1(n_817), .A2(n_122), .B(n_124), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_857), .B(n_124), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_763), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_791), .Y(n_879) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_779), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_776), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_881) );
INVx3_ASAP7_75t_L g882 ( .A(n_779), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_798), .B(n_128), .Y(n_883) );
OR2x6_ASAP7_75t_L g884 ( .A(n_774), .B(n_128), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_802), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_810), .Y(n_886) );
INVx3_ASAP7_75t_L g887 ( .A(n_779), .Y(n_887) );
AO31x2_ASAP7_75t_L g888 ( .A1(n_811), .A2(n_129), .A3(n_130), .B(n_223), .Y(n_888) );
INVx2_ASAP7_75t_SL g889 ( .A(n_860), .Y(n_889) );
NAND2xp5_ASAP7_75t_SL g890 ( .A(n_796), .B(n_129), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_837), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_763), .Y(n_892) );
INVx3_ASAP7_75t_L g893 ( .A(n_862), .Y(n_893) );
BUFx4f_ASAP7_75t_L g894 ( .A(n_860), .Y(n_894) );
INVx6_ASAP7_75t_L g895 ( .A(n_758), .Y(n_895) );
AOI21xp5_ASAP7_75t_SL g896 ( .A1(n_837), .A2(n_226), .B(n_227), .Y(n_896) );
OR2x6_ASAP7_75t_L g897 ( .A(n_863), .B(n_228), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_793), .B(n_230), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_801), .A2(n_241), .B1(n_252), .B2(n_253), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_868), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_868), .Y(n_901) );
BUFx6f_ASAP7_75t_L g902 ( .A(n_745), .Y(n_902) );
NAND2x1p5_ASAP7_75t_L g903 ( .A(n_818), .B(n_263), .Y(n_903) );
AO21x2_ASAP7_75t_L g904 ( .A1(n_787), .A2(n_264), .B(n_266), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_803), .B(n_267), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_790), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_780), .Y(n_907) );
NAND2x1p5_ASAP7_75t_L g908 ( .A(n_846), .B(n_272), .Y(n_908) );
BUFx4f_ASAP7_75t_SL g909 ( .A(n_840), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_780), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_756), .B(n_813), .Y(n_911) );
OAI21x1_ASAP7_75t_SL g912 ( .A1(n_782), .A2(n_841), .B(n_809), .Y(n_912) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_745), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_795), .B(n_800), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_825), .Y(n_915) );
INVx3_ASAP7_75t_L g916 ( .A(n_862), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_825), .Y(n_917) );
INVx3_ASAP7_75t_L g918 ( .A(n_745), .Y(n_918) );
BUFx3_ASAP7_75t_L g919 ( .A(n_790), .Y(n_919) );
AND2x4_ASAP7_75t_L g920 ( .A(n_816), .B(n_838), .Y(n_920) );
AND2x4_ASAP7_75t_L g921 ( .A(n_816), .B(n_834), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_805), .A2(n_765), .B1(n_854), .B2(n_773), .Y(n_922) );
AO21x2_ASAP7_75t_L g923 ( .A1(n_771), .A2(n_799), .B(n_764), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_853), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_794), .A2(n_784), .B1(n_808), .B2(n_797), .Y(n_925) );
OAI21xp5_ASAP7_75t_L g926 ( .A1(n_859), .A2(n_757), .B(n_746), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_762), .Y(n_927) );
AOI21xp5_ASAP7_75t_SL g928 ( .A1(n_814), .A2(n_852), .B(n_831), .Y(n_928) );
AOI21xp5_ASAP7_75t_L g929 ( .A1(n_842), .A2(n_833), .B(n_819), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_855), .Y(n_930) );
AO21x2_ASAP7_75t_L g931 ( .A1(n_851), .A2(n_788), .B(n_783), .Y(n_931) );
OAI21xp5_ASAP7_75t_L g932 ( .A1(n_861), .A2(n_786), .B(n_845), .Y(n_932) );
AO21x2_ASAP7_75t_L g933 ( .A1(n_804), .A2(n_778), .B(n_785), .Y(n_933) );
AOI21xp33_ASAP7_75t_L g934 ( .A1(n_755), .A2(n_827), .B(n_812), .Y(n_934) );
BUFx8_ASAP7_75t_L g935 ( .A(n_766), .Y(n_935) );
AND2x4_ASAP7_75t_L g936 ( .A(n_835), .B(n_826), .Y(n_936) );
INVx4_ASAP7_75t_L g937 ( .A(n_822), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_824), .B(n_848), .Y(n_938) );
INVxp67_ASAP7_75t_SL g939 ( .A(n_836), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_767), .B(n_749), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_829), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_770), .Y(n_942) );
INVx3_ASAP7_75t_L g943 ( .A(n_775), .Y(n_943) );
A2O1A1Ixp33_ASAP7_75t_L g944 ( .A1(n_777), .A2(n_769), .B(n_747), .C(n_768), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_829), .Y(n_945) );
AND3x2_ASAP7_75t_L g946 ( .A(n_821), .B(n_839), .C(n_753), .Y(n_946) );
NAND2xp33_ASAP7_75t_R g947 ( .A(n_760), .B(n_758), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_792), .B(n_830), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_849), .A2(n_823), .B(n_847), .Y(n_949) );
OAI21x1_ASAP7_75t_L g950 ( .A1(n_815), .A2(n_850), .B(n_792), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_829), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_844), .Y(n_952) );
BUFx8_ASAP7_75t_L g953 ( .A(n_766), .Y(n_953) );
A2O1A1Ixp33_ASAP7_75t_L g954 ( .A1(n_843), .A2(n_781), .B(n_792), .C(n_772), .Y(n_954) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_856), .A2(n_864), .B(n_867), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_864), .A2(n_867), .B(n_806), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_772), .B(n_844), .Y(n_957) );
NAND2x1p5_ASAP7_75t_L g958 ( .A(n_781), .B(n_772), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_828), .Y(n_959) );
NOR2x1_ASAP7_75t_R g960 ( .A(n_781), .B(n_806), .Y(n_960) );
OA21x2_ASAP7_75t_L g961 ( .A1(n_828), .A2(n_748), .B(n_752), .Y(n_961) );
OA21x2_ASAP7_75t_L g962 ( .A1(n_748), .A2(n_752), .B(n_751), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_807), .Y(n_963) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_754), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_807), .B(n_820), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_807), .B(n_820), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_817), .A2(n_657), .B1(n_642), .B2(n_631), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_857), .B(n_613), .Y(n_968) );
INVx3_ASAP7_75t_L g969 ( .A(n_779), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_807), .B(n_820), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_857), .B(n_600), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_857), .B(n_600), .Y(n_972) );
AND2x4_ASAP7_75t_L g973 ( .A(n_858), .B(n_866), .Y(n_973) );
AOI21x1_ASAP7_75t_L g974 ( .A1(n_761), .A2(n_751), .B(n_748), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_807), .Y(n_975) );
OAI21x1_ASAP7_75t_L g976 ( .A1(n_752), .A2(n_751), .B(n_741), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_754), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_807), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_807), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_807), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_807), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_807), .Y(n_982) );
INVx4_ASAP7_75t_SL g983 ( .A(n_754), .Y(n_983) );
BUFx2_ASAP7_75t_L g984 ( .A(n_754), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_817), .A2(n_631), .B1(n_590), .B2(n_669), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_807), .B(n_820), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_754), .Y(n_987) );
BUFx6f_ASAP7_75t_L g988 ( .A(n_779), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_820), .B(n_568), .Y(n_989) );
INVx4_ASAP7_75t_SL g990 ( .A(n_754), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_807), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_807), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_807), .Y(n_993) );
INVx1_ASAP7_75t_SL g994 ( .A(n_846), .Y(n_994) );
A2O1A1Ixp33_ASAP7_75t_L g995 ( .A1(n_832), .A2(n_735), .B(n_590), .C(n_865), .Y(n_995) );
BUFx8_ASAP7_75t_SL g996 ( .A(n_789), .Y(n_996) );
INVx4_ASAP7_75t_L g997 ( .A(n_754), .Y(n_997) );
OA21x2_ASAP7_75t_L g998 ( .A1(n_748), .A2(n_752), .B(n_751), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_915), .B(n_917), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_968), .B(n_989), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_963), .B(n_978), .Y(n_1001) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_894), .Y(n_1002) );
AO21x2_ASAP7_75t_L g1003 ( .A1(n_955), .A2(n_956), .B(n_912), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_979), .B(n_982), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_879), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_965), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_885), .B(n_886), .Y(n_1007) );
OA21x2_ASAP7_75t_L g1008 ( .A1(n_976), .A2(n_957), .B(n_954), .Y(n_1008) );
OAI21xp5_ASAP7_75t_L g1009 ( .A1(n_995), .A2(n_944), .B(n_949), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_971), .B(n_972), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_919), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_975), .B(n_980), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_966), .B(n_970), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_981), .B(n_991), .Y(n_1014) );
AO21x2_ASAP7_75t_L g1015 ( .A1(n_957), .A2(n_974), .B(n_945), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_992), .B(n_993), .Y(n_1016) );
AOI21x1_ASAP7_75t_L g1017 ( .A1(n_962), .A2(n_998), .B(n_961), .Y(n_1017) );
NOR2xp33_ASAP7_75t_SL g1018 ( .A(n_997), .B(n_909), .Y(n_1018) );
INVx4_ASAP7_75t_SL g1019 ( .A(n_897), .Y(n_1019) );
AO21x2_ASAP7_75t_L g1020 ( .A1(n_941), .A2(n_952), .B(n_951), .Y(n_1020) );
INVx2_ASAP7_75t_SL g1021 ( .A(n_880), .Y(n_1021) );
AO21x2_ASAP7_75t_L g1022 ( .A1(n_948), .A2(n_923), .B(n_929), .Y(n_1022) );
OAI221xp5_ASAP7_75t_SL g1023 ( .A1(n_985), .A2(n_967), .B1(n_925), .B2(n_884), .C(n_922), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1024 ( .A(n_897), .B(n_927), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_986), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_959), .Y(n_1026) );
INVx3_ASAP7_75t_L g1027 ( .A(n_880), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_961), .Y(n_1028) );
INVx3_ASAP7_75t_L g1029 ( .A(n_880), .Y(n_1029) );
AO21x2_ASAP7_75t_L g1030 ( .A1(n_923), .A2(n_950), .B(n_933), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_877), .B(n_883), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_882), .B(n_887), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_936), .B(n_994), .Y(n_1033) );
BUFx3_ASAP7_75t_L g1034 ( .A(n_988), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_900), .A2(n_901), .B1(n_890), .B2(n_922), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_940), .B(n_907), .Y(n_1036) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_988), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_936), .B(n_878), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_937), .B(n_973), .Y(n_1039) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_891), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1041 ( .A(n_988), .Y(n_1041) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_882), .Y(n_1042) );
INVx3_ASAP7_75t_L g1043 ( .A(n_902), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_873), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_892), .B(n_910), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_924), .B(n_930), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_887), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_869), .Y(n_1048) );
NOR2x1_ASAP7_75t_L g1049 ( .A(n_884), .B(n_897), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_875), .Y(n_1050) );
OR2x6_ASAP7_75t_L g1051 ( .A(n_908), .B(n_896), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_969), .B(n_918), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_906), .Y(n_1053) );
OAI21xp5_ASAP7_75t_L g1054 ( .A1(n_934), .A2(n_932), .B(n_926), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_937), .B(n_938), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_902), .Y(n_1056) );
INVx3_ASAP7_75t_L g1057 ( .A(n_902), .Y(n_1057) );
CKINVDCx14_ASAP7_75t_R g1058 ( .A(n_984), .Y(n_1058) );
INVx2_ASAP7_75t_L g1059 ( .A(n_913), .Y(n_1059) );
AO21x2_ASAP7_75t_L g1060 ( .A1(n_933), .A2(n_931), .B(n_928), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_913), .Y(n_1061) );
BUFx12f_ASAP7_75t_L g1062 ( .A(n_889), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_913), .Y(n_1063) );
INVx3_ASAP7_75t_L g1064 ( .A(n_969), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_870), .Y(n_1065) );
INVx5_ASAP7_75t_SL g1066 ( .A(n_983), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_911), .B(n_942), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_987), .Y(n_1068) );
AO21x2_ASAP7_75t_L g1069 ( .A1(n_904), .A2(n_914), .B(n_872), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_911), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_876), .B(n_914), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_898), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_876), .B(n_958), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_893), .B(n_916), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_935), .A2(n_953), .B1(n_946), .B2(n_881), .Y(n_1075) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_895), .A2(n_947), .B1(n_977), .B2(n_964), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_905), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_920), .B(n_895), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_893), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1080 ( .A(n_871), .Y(n_1080) );
INVx3_ASAP7_75t_L g1081 ( .A(n_918), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_943), .B(n_920), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_943), .Y(n_1083) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_983), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_990), .Y(n_1085) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_990), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_874), .Y(n_1087) );
INVx4_ASAP7_75t_SL g1088 ( .A(n_888), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_921), .B(n_899), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_921), .B(n_888), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_939), .B(n_888), .Y(n_1091) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_1037), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1012), .B(n_960), .Y(n_1093) );
BUFx2_ASAP7_75t_SL g1094 ( .A(n_1085), .Y(n_1094) );
AND2x4_ASAP7_75t_L g1095 ( .A(n_1090), .B(n_935), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_999), .B(n_903), .Y(n_1096) );
BUFx2_ASAP7_75t_L g1097 ( .A(n_1024), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1026), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_999), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1020), .Y(n_1100) );
INVxp67_ASAP7_75t_L g1101 ( .A(n_1055), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1020), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_1000), .B(n_996), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_1049), .Y(n_1104) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1028), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_1013), .B(n_1033), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_1024), .B(n_1010), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1014), .B(n_1016), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_1024), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1016), .B(n_1001), .Y(n_1110) );
NAND2x1_ASAP7_75t_L g1111 ( .A(n_1024), .B(n_1089), .Y(n_1111) );
AO21x2_ASAP7_75t_L g1112 ( .A1(n_1054), .A2(n_1009), .B(n_1017), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1001), .B(n_1004), .Y(n_1113) );
BUFx2_ASAP7_75t_L g1114 ( .A(n_1019), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1067), .B(n_1007), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_1067), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1015), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1007), .B(n_1005), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1070), .B(n_1006), .Y(n_1119) );
BUFx3_ASAP7_75t_L g1120 ( .A(n_1062), .Y(n_1120) );
INVx4_ASAP7_75t_L g1121 ( .A(n_1019), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1073), .B(n_1003), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1025), .B(n_1046), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1046), .B(n_1071), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_1042), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1071), .B(n_1089), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1036), .B(n_1055), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_1062), .Y(n_1128) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_1019), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1073), .B(n_1008), .Y(n_1130) );
BUFx3_ASAP7_75t_L g1131 ( .A(n_1034), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1035), .B(n_1065), .Y(n_1132) );
BUFx3_ASAP7_75t_L g1133 ( .A(n_1034), .Y(n_1133) );
INVx4_ASAP7_75t_L g1134 ( .A(n_1051), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1008), .B(n_1040), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1038), .B(n_1035), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1137 ( .A(n_1003), .B(n_1091), .Y(n_1137) );
AND2x2_ASAP7_75t_SL g1138 ( .A(n_1075), .B(n_1091), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1040), .B(n_1053), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1048), .B(n_1031), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1141 ( .A(n_1072), .B(n_1077), .Y(n_1141) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1091), .B(n_1088), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_1061), .Y(n_1143) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_1037), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_1032), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_1002), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1126), .B(n_1030), .Y(n_1147) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1105), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1149 ( .A1(n_1101), .A2(n_1075), .B1(n_1050), .B2(n_1058), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1124), .B(n_1060), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1141), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1105), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1124), .B(n_1060), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1093), .B(n_1022), .Y(n_1154) );
INVx4_ASAP7_75t_L g1155 ( .A(n_1121), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1093), .B(n_1022), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1157 ( .A(n_1122), .B(n_1088), .Y(n_1157) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1116), .B(n_1039), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1108), .B(n_1044), .Y(n_1159) );
INVx4_ASAP7_75t_L g1160 ( .A(n_1121), .Y(n_1160) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_1114), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1110), .B(n_1082), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1130), .B(n_1069), .Y(n_1163) );
BUFx3_ASAP7_75t_L g1164 ( .A(n_1131), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1123), .B(n_1082), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1099), .B(n_1023), .Y(n_1166) );
BUFx2_ASAP7_75t_L g1167 ( .A(n_1114), .Y(n_1167) );
NOR2xp33_ASAP7_75t_SL g1168 ( .A(n_1120), .B(n_1018), .Y(n_1168) );
OAI21xp5_ASAP7_75t_L g1169 ( .A1(n_1132), .A2(n_1076), .B(n_1080), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1115), .B(n_1068), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1171 ( .A(n_1103), .B(n_1078), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1115), .B(n_1056), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1113), .B(n_1063), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1095), .B(n_1059), .Y(n_1174) );
NAND2x1p5_ASAP7_75t_L g1175 ( .A(n_1121), .B(n_1064), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_1125), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1118), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1119), .B(n_1083), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1119), .B(n_1011), .Y(n_1179) );
NAND2x1_ASAP7_75t_L g1180 ( .A(n_1121), .B(n_1051), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g1181 ( .A(n_1139), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1106), .B(n_1047), .Y(n_1182) );
AND2x4_ASAP7_75t_L g1183 ( .A(n_1122), .B(n_1057), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1107), .B(n_1045), .Y(n_1184) );
NAND2x1p5_ASAP7_75t_L g1185 ( .A(n_1155), .B(n_1086), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1186 ( .A(n_1157), .B(n_1137), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1150), .B(n_1135), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1176), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1181), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1151), .Y(n_1190) );
BUFx3_ASAP7_75t_L g1191 ( .A(n_1164), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1170), .B(n_1127), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1153), .B(n_1135), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1148), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1158), .B(n_1111), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1148), .Y(n_1196) );
INVx3_ASAP7_75t_L g1197 ( .A(n_1155), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1166), .B(n_1104), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1199 ( .A(n_1158), .B(n_1111), .Y(n_1199) );
INVxp67_ASAP7_75t_SL g1200 ( .A(n_1152), .Y(n_1200) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1166), .B(n_1096), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1177), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1172), .B(n_1138), .Y(n_1203) );
NAND2x1p5_ASAP7_75t_L g1204 ( .A(n_1160), .B(n_1129), .Y(n_1204) );
NAND2xp5_ASAP7_75t_SL g1205 ( .A(n_1160), .B(n_1129), .Y(n_1205) );
INVx2_ASAP7_75t_SL g1206 ( .A(n_1164), .Y(n_1206) );
NAND2xp5_ASAP7_75t_SL g1207 ( .A(n_1161), .B(n_1134), .Y(n_1207) );
INVx1_ASAP7_75t_SL g1208 ( .A(n_1179), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1178), .Y(n_1209) );
INVx3_ASAP7_75t_L g1210 ( .A(n_1180), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1173), .B(n_1098), .Y(n_1211) );
OR3x2_ASAP7_75t_L g1212 ( .A(n_1168), .B(n_1066), .C(n_1096), .Y(n_1212) );
INVxp67_ASAP7_75t_SL g1213 ( .A(n_1188), .Y(n_1213) );
AND2x4_ASAP7_75t_L g1214 ( .A(n_1186), .B(n_1157), .Y(n_1214) );
O2A1O1Ixp33_ASAP7_75t_L g1215 ( .A1(n_1205), .A2(n_1128), .B(n_1084), .C(n_1087), .Y(n_1215) );
INVx3_ASAP7_75t_L g1216 ( .A(n_1197), .Y(n_1216) );
AOI21xp33_ASAP7_75t_L g1217 ( .A1(n_1198), .A2(n_1169), .B(n_1171), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_1188), .Y(n_1218) );
INVx1_ASAP7_75t_SL g1219 ( .A(n_1191), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1220 ( .A1(n_1201), .A2(n_1140), .B1(n_1159), .B2(n_1165), .C(n_1162), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_1198), .A2(n_1149), .B1(n_1156), .B2(n_1154), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1222 ( .A(n_1211), .B(n_1147), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1194), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1209), .B(n_1154), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1189), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_1212), .A2(n_1134), .B1(n_1167), .B2(n_1094), .Y(n_1226) );
INVxp67_ASAP7_75t_L g1227 ( .A(n_1206), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g1228 ( .A1(n_1197), .A2(n_1097), .B1(n_1109), .B2(n_1094), .Y(n_1228) );
NOR2xp67_ASAP7_75t_SL g1229 ( .A(n_1210), .B(n_1146), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1196), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1202), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1190), .Y(n_1232) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1223), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_1217), .A2(n_1212), .B1(n_1208), .B2(n_1192), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1218), .B(n_1187), .Y(n_1235) );
INVxp33_ASAP7_75t_L g1236 ( .A(n_1229), .Y(n_1236) );
INVxp67_ASAP7_75t_L g1237 ( .A(n_1219), .Y(n_1237) );
AOI22xp5_ASAP7_75t_L g1238 ( .A1(n_1221), .A2(n_1203), .B1(n_1186), .B2(n_1199), .Y(n_1238) );
OAI221xp5_ASAP7_75t_L g1239 ( .A1(n_1215), .A2(n_1220), .B1(n_1228), .B2(n_1227), .C(n_1213), .Y(n_1239) );
OAI21xp33_ASAP7_75t_L g1240 ( .A1(n_1224), .A2(n_1195), .B(n_1193), .Y(n_1240) );
AOI31xp33_ASAP7_75t_L g1241 ( .A1(n_1226), .A2(n_1185), .A3(n_1204), .B(n_1207), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1232), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1231), .Y(n_1243) );
NOR2x1_ASAP7_75t_L g1244 ( .A(n_1216), .B(n_1214), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1225), .B(n_1163), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1242), .Y(n_1246) );
INVxp67_ASAP7_75t_L g1247 ( .A(n_1237), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1243), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g1249 ( .A1(n_1241), .A2(n_1200), .B(n_1230), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_1234), .A2(n_1222), .B1(n_1182), .B2(n_1175), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1235), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_1236), .A2(n_1066), .B1(n_1175), .B2(n_1184), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1245), .Y(n_1253) );
AOI211xp5_ASAP7_75t_L g1254 ( .A1(n_1236), .A2(n_1136), .B(n_1183), .C(n_1146), .Y(n_1254) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_1238), .B(n_1102), .C(n_1100), .Y(n_1255) );
INVxp67_ASAP7_75t_SL g1256 ( .A(n_1244), .Y(n_1256) );
A2O1A1Ixp33_ASAP7_75t_L g1257 ( .A1(n_1240), .A2(n_1133), .B(n_1145), .C(n_1142), .Y(n_1257) );
NOR2x1_ASAP7_75t_L g1258 ( .A(n_1233), .B(n_1133), .Y(n_1258) );
XOR2x2_ASAP7_75t_L g1259 ( .A(n_1239), .B(n_1174), .Y(n_1259) );
INVx1_ASAP7_75t_SL g1260 ( .A(n_1258), .Y(n_1260) );
O2A1O1Ixp33_ASAP7_75t_L g1261 ( .A1(n_1247), .A2(n_1250), .B(n_1256), .C(n_1252), .Y(n_1261) );
OAI221xp5_ASAP7_75t_L g1262 ( .A1(n_1249), .A2(n_1259), .B1(n_1257), .B2(n_1255), .C(n_1254), .Y(n_1262) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1251), .B(n_1253), .Y(n_1263) );
NOR3xp33_ASAP7_75t_L g1264 ( .A(n_1261), .B(n_1246), .C(n_1248), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1263), .B(n_1112), .Y(n_1265) );
AND2x4_ASAP7_75t_L g1266 ( .A(n_1260), .B(n_1174), .Y(n_1266) );
NOR2x1_ASAP7_75t_L g1267 ( .A(n_1262), .B(n_1064), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1265), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1264), .Y(n_1269) );
NAND2x1p5_ASAP7_75t_L g1270 ( .A(n_1267), .B(n_1021), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1269), .Y(n_1271) );
OAI22x1_ASAP7_75t_L g1272 ( .A1(n_1270), .A2(n_1266), .B1(n_1041), .B2(n_1052), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1268), .Y(n_1273) );
XOR2xp5_ASAP7_75t_L g1274 ( .A(n_1273), .B(n_1052), .Y(n_1274) );
OAI22x1_ASAP7_75t_SL g1275 ( .A1(n_1271), .A2(n_1041), .B1(n_1027), .B2(n_1029), .Y(n_1275) );
OA21x2_ASAP7_75t_L g1276 ( .A1(n_1274), .A2(n_1272), .B(n_1079), .Y(n_1276) );
AOI22x1_ASAP7_75t_L g1277 ( .A1(n_1275), .A2(n_1029), .B1(n_1074), .B2(n_1143), .Y(n_1277) );
OAI21xp5_ASAP7_75t_L g1278 ( .A1(n_1277), .A2(n_1043), .B(n_1081), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1278), .B(n_1276), .Y(n_1279) );
AOI21xp5_ASAP7_75t_L g1280 ( .A1(n_1279), .A2(n_1092), .B(n_1144), .Y(n_1280) );
AOI21xp5_ASAP7_75t_L g1281 ( .A1(n_1280), .A2(n_1081), .B(n_1117), .Y(n_1281) );
endmodule