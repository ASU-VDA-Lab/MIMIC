module real_jpeg_8922_n_16 (n_5, n_4, n_8, n_0, n_12, n_303, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_303;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_300;
wire n_292;
wire n_286;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_197;
wire n_173;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_293;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_128;
wire n_295;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx24_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_7),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_66),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_66),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_8),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_143),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_143),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_8),
.A2(n_40),
.B1(n_50),
.B2(n_143),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_9),
.A2(n_58),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_58),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_9),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_9),
.A2(n_27),
.B1(n_33),
.B2(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_52),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_42),
.B(n_46),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_9),
.A2(n_40),
.B1(n_50),
.B2(n_161),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_40),
.B1(n_50),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_10),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_101),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_101),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_101),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_36),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_12),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_12),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_13),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_152),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_152),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_13),
.A2(n_40),
.B1(n_50),
.B2(n_152),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_14),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_40),
.B1(n_50),
.B2(n_75),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_75),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_40),
.B1(n_50),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_15),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_20),
.B(n_109),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_21),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_21),
.B(n_294),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_71),
.CI(n_90),
.CON(n_21),
.SN(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_55),
.B2(n_70),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_25),
.A2(n_38),
.B(n_70),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_25),
.A2(n_26),
.B1(n_56),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_27),
.A2(n_33),
.B1(n_142),
.B2(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_27),
.A2(n_95),
.B(n_145),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_27),
.A2(n_34),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_27),
.A2(n_33),
.B1(n_208),
.B2(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_27),
.A2(n_194),
.B(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_28),
.B(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_28),
.A2(n_32),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_29),
.A2(n_30),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_29),
.B(n_64),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_29),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_30),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_32),
.B(n_94),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_33),
.B(n_161),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_33),
.A2(n_93),
.B(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_48),
.B(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_39),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_39),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_39),
.A2(n_44),
.B1(n_244),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_39),
.A2(n_44),
.B1(n_100),
.B2(n_253),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_40),
.A2(n_41),
.B(n_161),
.C(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_44),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_77),
.B(n_79),
.C(n_80),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_77),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_46),
.B(n_161),
.CON(n_186),
.SN(n_186)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_52),
.A2(n_117),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_56),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_65),
.B(n_67),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_63),
.B1(n_65),
.B2(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_57),
.A2(n_63),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_57),
.A2(n_63),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_57),
.A2(n_63),
.B1(n_151),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_57),
.A2(n_63),
.B1(n_176),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_57),
.A2(n_83),
.B(n_184),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_59),
.B1(n_77),
.B2(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_58),
.B(n_77),
.Y(n_192)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_59),
.A2(n_79),
.B1(n_186),
.B2(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_63),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_63),
.A2(n_86),
.B(n_97),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_68),
.A2(n_85),
.B(n_88),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_82),
.B(n_89),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_82),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_76),
.A2(n_80),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_76),
.A2(n_124),
.B(n_256),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_80),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_111),
.B1(n_112),
.B2(n_129),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_89),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.C(n_103),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_91),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_92),
.B(n_96),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_105),
.A2(n_121),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_105),
.A2(n_121),
.B1(n_204),
.B2(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_130),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_121),
.A2(n_240),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI321xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_281),
.A3(n_293),
.B1(n_295),
.B2(n_301),
.C(n_303),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_246),
.C(n_277),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_220),
.B(n_245),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_197),
.B(n_219),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_179),
.B(n_196),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_170),
.B(n_178),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_158),
.B(n_169),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_153),
.B2(n_157),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_157),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_180),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.CI(n_177),
.CON(n_173),
.SN(n_173)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_190),
.B2(n_195),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_189),
.C(n_195),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_213),
.B2(n_214),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_216),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_205),
.B1(n_206),
.B2(n_212),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_209),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_210),
.C(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_222),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_233),
.C(n_234),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_229),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_241),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_238),
.C(n_241),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_246),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_264),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_264),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_258),
.C(n_262),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_251),
.C(n_257),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_257),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_254),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_261),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_273),
.C(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_269),
.C(n_272),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_296),
.B(n_300),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_284),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_290),
.C(n_292),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B(n_299),
.Y(n_296)
);


endmodule