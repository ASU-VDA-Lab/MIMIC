module real_aes_16500_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_841, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_841;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g115 ( .A(n_0), .B(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_1), .A2(n_4), .B1(n_143), .B2(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_2), .A2(n_42), .B1(n_150), .B2(n_186), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_3), .A2(n_24), .B1(n_186), .B2(n_228), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_5), .A2(n_16), .B1(n_140), .B2(n_217), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_6), .A2(n_62), .B1(n_200), .B2(n_230), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_7), .A2(n_17), .B1(n_150), .B2(n_171), .Y(n_621) );
INVx1_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_9), .A2(n_473), .B(n_830), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_10), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_11), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_12), .A2(n_18), .B1(n_199), .B2(n_202), .Y(n_198) );
OR2x2_ASAP7_75t_L g108 ( .A(n_13), .B(n_37), .Y(n_108) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_15), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_19), .A2(n_101), .B1(n_140), .B2(n_143), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_20), .A2(n_38), .B1(n_175), .B2(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_21), .B(n_141), .Y(n_172) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_22), .A2(n_58), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_23), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_25), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_26), .B(n_147), .Y(n_541) );
INVx4_ASAP7_75t_R g589 ( .A(n_27), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_28), .A2(n_47), .B1(n_188), .B2(n_189), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_29), .A2(n_55), .B1(n_140), .B2(n_189), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_30), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_31), .B(n_175), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_32), .Y(n_251) );
INVx1_ASAP7_75t_L g520 ( .A(n_33), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_34), .B(n_186), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_SL g532 ( .A1(n_35), .A2(n_146), .B(n_150), .C(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_36), .A2(n_56), .B1(n_150), .B2(n_189), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_39), .A2(n_88), .B1(n_150), .B2(n_227), .Y(n_226) );
XOR2x2_ASAP7_75t_L g823 ( .A(n_40), .B(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_41), .A2(n_45), .B1(n_150), .B2(n_171), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_43), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_44), .A2(n_60), .B1(n_140), .B2(n_149), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_46), .A2(n_74), .B1(n_825), .B2(n_826), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_46), .Y(n_826) );
INVx1_ASAP7_75t_L g544 ( .A(n_48), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_49), .B(n_150), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_50), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_51), .Y(n_561) );
INVx2_ASAP7_75t_L g481 ( .A(n_52), .Y(n_481) );
INVx1_ASAP7_75t_L g111 ( .A(n_53), .Y(n_111) );
BUFx3_ASAP7_75t_L g490 ( .A(n_53), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_54), .A2(n_119), .B(n_469), .Y(n_118) );
AOI31xp33_ASAP7_75t_L g469 ( .A1(n_54), .A2(n_470), .A3(n_472), .B(n_473), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_57), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_59), .A2(n_89), .B1(n_150), .B2(n_189), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_61), .A2(n_69), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_61), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_63), .A2(n_77), .B1(n_149), .B2(n_188), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_64), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_65), .A2(n_79), .B1(n_150), .B2(n_171), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_66), .A2(n_100), .B1(n_140), .B2(n_202), .Y(n_248) );
AND2x4_ASAP7_75t_L g136 ( .A(n_67), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g159 ( .A(n_68), .Y(n_159) );
INVx1_ASAP7_75t_L g122 ( .A(n_69), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_70), .A2(n_92), .B1(n_188), .B2(n_189), .Y(n_516) );
AO22x1_ASAP7_75t_L g578 ( .A1(n_71), .A2(n_78), .B1(n_214), .B2(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g137 ( .A(n_72), .Y(n_137) );
AND2x2_ASAP7_75t_L g536 ( .A(n_73), .B(n_181), .Y(n_536) );
INVx1_ASAP7_75t_L g825 ( .A(n_74), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_75), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_76), .B(n_230), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_80), .B(n_186), .Y(n_562) );
INVx2_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_82), .B(n_181), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_83), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_84), .A2(n_99), .B1(n_189), .B2(n_230), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_85), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_86), .B(n_157), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_87), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_90), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_91), .B(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_93), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_94), .B(n_181), .Y(n_558) );
INVx1_ASAP7_75t_L g114 ( .A(n_95), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_95), .B(n_467), .Y(n_466) );
NAND2xp33_ASAP7_75t_L g177 ( .A(n_96), .B(n_141), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_97), .A2(n_205), .B(n_230), .C(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g591 ( .A(n_98), .B(n_592), .Y(n_591) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_102), .B(n_176), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_117), .B(n_837), .Y(n_103) );
CKINVDCx11_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx6_ASAP7_75t_L g839 ( .A(n_105), .Y(n_839) );
NAND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g468 ( .A(n_108), .Y(n_468) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_108), .B(n_490), .Y(n_836) );
NOR2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g467 ( .A(n_111), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g496 ( .A(n_114), .Y(n_496) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_477), .B(n_482), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_463), .Y(n_119) );
INVx1_ASAP7_75t_L g472 ( .A(n_120), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
INVx2_ASAP7_75t_L g497 ( .A(n_124), .Y(n_497) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_366), .Y(n_124) );
NAND4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_290), .C(n_321), .D(n_350), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_257), .Y(n_126) );
OAI322xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_193), .A3(n_222), .B1(n_235), .B2(n_243), .C1(n_252), .C2(n_254), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_129), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_163), .Y(n_129) );
AND2x2_ASAP7_75t_L g287 ( .A(n_130), .B(n_288), .Y(n_287) );
INVx4_ASAP7_75t_L g323 ( .A(n_130), .Y(n_323) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g298 ( .A(n_131), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g301 ( .A(n_131), .B(n_195), .Y(n_301) );
AND2x2_ASAP7_75t_L g318 ( .A(n_131), .B(n_211), .Y(n_318) );
AND2x2_ASAP7_75t_L g416 ( .A(n_131), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g239 ( .A(n_132), .Y(n_239) );
AND2x4_ASAP7_75t_L g422 ( .A(n_132), .B(n_417), .Y(n_422) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .A3(n_154), .B(n_160), .Y(n_132) );
AO31x2_ASAP7_75t_L g246 ( .A1(n_133), .A2(n_206), .A3(n_247), .B(n_250), .Y(n_246) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_134), .A2(n_584), .B(n_587), .Y(n_583) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AO31x2_ASAP7_75t_L g183 ( .A1(n_135), .A2(n_184), .A3(n_190), .B(n_191), .Y(n_183) );
AO31x2_ASAP7_75t_L g196 ( .A1(n_135), .A2(n_197), .A3(n_206), .B(n_208), .Y(n_196) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_135), .A2(n_212), .A3(n_219), .B(n_220), .Y(n_211) );
AO31x2_ASAP7_75t_L g619 ( .A1(n_135), .A2(n_162), .A3(n_620), .B(n_623), .Y(n_619) );
BUFx10_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
BUFx10_ASAP7_75t_L g511 ( .A(n_136), .Y(n_511) );
INVx1_ASAP7_75t_L g535 ( .A(n_136), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B1(n_148), .B2(n_151), .Y(n_138) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_141), .Y(n_579) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g144 ( .A(n_142), .Y(n_144) );
INVx3_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g201 ( .A(n_142), .Y(n_201) );
INVx1_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
INVx1_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
INVx2_ASAP7_75t_L g228 ( .A(n_142), .Y(n_228) );
INVx1_ASAP7_75t_L g230 ( .A(n_142), .Y(n_230) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_144), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_145), .A2(n_174), .B(n_177), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_145), .A2(n_151), .B1(n_185), .B2(n_187), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_145), .A2(n_198), .B1(n_203), .B2(n_204), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_145), .A2(n_151), .B1(n_213), .B2(n_216), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_145), .A2(n_226), .B1(n_229), .B2(n_231), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_145), .A2(n_204), .B1(n_248), .B2(n_249), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_145), .A2(n_151), .B1(n_267), .B2(n_268), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_145), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_145), .A2(n_231), .B1(n_516), .B2(n_517), .Y(n_515) );
OAI22x1_ASAP7_75t_L g620 ( .A1(n_145), .A2(n_231), .B1(n_621), .B2(n_622), .Y(n_620) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
O2A1O1Ixp5_ASAP7_75t_L g169 ( .A1(n_146), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_146), .A2(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_146), .B(n_578), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_146), .A2(n_574), .B(n_578), .C(n_581), .Y(n_635) );
BUFx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
INVx1_ASAP7_75t_L g531 ( .A(n_147), .Y(n_531) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g510 ( .A(n_152), .Y(n_510) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g564 ( .A(n_153), .Y(n_564) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_154), .A2(n_232), .A3(n_266), .B(n_269), .Y(n_265) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_154), .A2(n_583), .B(n_591), .Y(n_582) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_SL g208 ( .A(n_156), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_156), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
INVx2_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_157), .A2(n_535), .B(n_576), .Y(n_581) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_162), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g427 ( .A(n_163), .B(n_328), .Y(n_427) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g256 ( .A(n_164), .Y(n_256) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_164), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_182), .Y(n_164) );
AND2x2_ASAP7_75t_L g244 ( .A(n_165), .B(n_183), .Y(n_244) );
INVx1_ASAP7_75t_L g285 ( .A(n_165), .Y(n_285) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_180), .Y(n_165) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_166), .A2(n_168), .B(n_180), .Y(n_280) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g181 ( .A(n_167), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_167), .B(n_192), .Y(n_191) );
BUFx3_ASAP7_75t_L g219 ( .A(n_167), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_167), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_167), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g548 ( .A(n_167), .B(n_511), .Y(n_548) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_178), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_171), .A2(n_561), .B(n_562), .C(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g188 ( .A(n_176), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_176), .A2(n_218), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_SL g232 ( .A(n_179), .Y(n_232) );
INVx2_ASAP7_75t_L g190 ( .A(n_181), .Y(n_190) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_181), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g276 ( .A(n_182), .Y(n_276) );
AND2x2_ASAP7_75t_L g340 ( .A(n_182), .B(n_279), .Y(n_340) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g294 ( .A(n_183), .Y(n_294) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_183), .Y(n_347) );
OR2x2_ASAP7_75t_L g418 ( .A(n_183), .B(n_224), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_186), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g518 ( .A(n_189), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_189), .B(n_543), .Y(n_542) );
AO31x2_ASAP7_75t_L g506 ( .A1(n_190), .A2(n_507), .A3(n_511), .B(n_512), .Y(n_506) );
NAND4xp25_ASAP7_75t_L g296 ( .A(n_193), .B(n_297), .C(n_300), .D(n_302), .Y(n_296) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g434 ( .A(n_194), .B(n_422), .Y(n_434) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_210), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_195), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g288 ( .A(n_195), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g308 ( .A(n_195), .Y(n_308) );
INVx1_ASAP7_75t_L g325 ( .A(n_195), .Y(n_325) );
INVx1_ASAP7_75t_L g333 ( .A(n_195), .Y(n_333) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_195), .Y(n_447) );
INVx4_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_196), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g365 ( .A(n_196), .B(n_265), .Y(n_365) );
AND2x2_ASAP7_75t_L g373 ( .A(n_196), .B(n_211), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_196), .B(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g438 ( .A(n_196), .Y(n_438) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_201), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
AO31x2_ASAP7_75t_L g514 ( .A1(n_206), .A2(n_232), .A3(n_515), .B(n_519), .Y(n_514) );
AOI21x1_ASAP7_75t_L g523 ( .A1(n_206), .A2(n_524), .B(n_536), .Y(n_523) );
BUFx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_207), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_207), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g592 ( .A(n_207), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_207), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g242 ( .A(n_211), .Y(n_242) );
OR2x2_ASAP7_75t_L g303 ( .A(n_211), .B(n_265), .Y(n_303) );
INVx2_ASAP7_75t_L g310 ( .A(n_211), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_211), .B(n_263), .Y(n_334) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_211), .Y(n_421) );
OAI21xp33_ASAP7_75t_SL g540 ( .A1(n_214), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_219), .A2(n_225), .A3(n_232), .B(n_233), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_222), .B(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g245 ( .A(n_224), .B(n_246), .Y(n_245) );
BUFx2_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
INVx2_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
AND2x4_ASAP7_75t_L g305 ( .A(n_224), .B(n_277), .Y(n_305) );
OR2x2_ASAP7_75t_L g385 ( .A(n_224), .B(n_285), .Y(n_385) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_228), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_231), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_237), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g302 ( .A(n_237), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_237), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_238), .B(n_308), .Y(n_316) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
OR2x2_ASAP7_75t_L g354 ( .A(n_239), .B(n_264), .Y(n_354) );
INVx1_ASAP7_75t_L g281 ( .A(n_240), .Y(n_281) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g253 ( .A(n_241), .Y(n_253) );
INVx1_ASAP7_75t_L g289 ( .A(n_242), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
OAI322xp33_ASAP7_75t_L g257 ( .A1(n_244), .A2(n_258), .A3(n_271), .B1(n_274), .B2(n_281), .C1(n_282), .C2(n_286), .Y(n_257) );
AND2x4_ASAP7_75t_L g304 ( .A(n_244), .B(n_305), .Y(n_304) );
AOI211xp5_ASAP7_75t_SL g335 ( .A1(n_244), .A2(n_336), .B(n_337), .C(n_341), .Y(n_335) );
AND2x2_ASAP7_75t_L g355 ( .A(n_244), .B(n_245), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_244), .B(n_272), .Y(n_361) );
AND2x4_ASAP7_75t_SL g283 ( .A(n_245), .B(n_284), .Y(n_283) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_245), .B(n_301), .C(n_329), .Y(n_374) );
AND2x2_ASAP7_75t_L g405 ( .A(n_245), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g272 ( .A(n_246), .B(n_273), .Y(n_272) );
INVx3_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
BUFx2_ASAP7_75t_L g345 ( .A(n_246), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_255), .B(n_279), .Y(n_278) );
NAND2x1_ASAP7_75t_L g319 ( .A(n_255), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g338 ( .A(n_255), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_256), .B(n_272), .Y(n_403) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g346 ( .A(n_261), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_265), .Y(n_299) );
AND2x4_ASAP7_75t_L g309 ( .A(n_265), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g396 ( .A(n_265), .Y(n_396) );
INVx2_ASAP7_75t_L g417 ( .A(n_265), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_271), .A2(n_430), .B1(n_432), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g341 ( .A(n_272), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g295 ( .A(n_273), .B(n_279), .Y(n_295) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x4_ASAP7_75t_L g284 ( .A(n_276), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g406 ( .A(n_276), .Y(n_406) );
INVx2_ASAP7_75t_L g292 ( .A(n_277), .Y(n_292) );
AND2x2_ASAP7_75t_L g320 ( .A(n_277), .B(n_279), .Y(n_320) );
INVx3_ASAP7_75t_L g328 ( .A(n_277), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_277), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g329 ( .A(n_280), .Y(n_329) );
OAI222xp33_ASAP7_75t_L g452 ( .A1(n_282), .A2(n_442), .B1(n_453), .B2(n_456), .C1(n_458), .C2(n_460), .Y(n_452) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g393 ( .A(n_284), .Y(n_393) );
AND2x2_ASAP7_75t_L g457 ( .A(n_284), .B(n_327), .Y(n_457) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_287), .B(n_378), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_296), .B1(n_304), .B2(n_306), .C(n_311), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g379 ( .A(n_292), .Y(n_379) );
INVx2_ASAP7_75t_L g441 ( .A(n_293), .Y(n_441) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g342 ( .A(n_294), .Y(n_342) );
AND2x2_ASAP7_75t_L g378 ( .A(n_294), .B(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g344 ( .A(n_295), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g370 ( .A(n_295), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g459 ( .A(n_295), .Y(n_459) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g408 ( .A(n_299), .Y(n_408) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g431 ( .A(n_301), .B(n_309), .Y(n_431) );
AND2x2_ASAP7_75t_L g454 ( .A(n_301), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g315 ( .A(n_303), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g450 ( .A(n_303), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_304), .A2(n_358), .B1(n_392), .B2(n_394), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_304), .A2(n_420), .B(n_423), .Y(n_419) );
INVxp67_ASAP7_75t_L g336 ( .A(n_305), .Y(n_336) );
INVx2_ASAP7_75t_SL g440 ( .A(n_305), .Y(n_440) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
OR2x2_ASAP7_75t_L g353 ( .A(n_307), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g451 ( .A(n_307), .B(n_450), .Y(n_451) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g324 ( .A(n_309), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_309), .B(n_333), .Y(n_349) );
INVx2_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_317), .B2(n_319), .Y(n_311) );
NOR2xp33_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_313), .A2(n_387), .B1(n_400), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g409 ( .A(n_318), .B(n_410), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_326), .B(n_330), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g390 ( .A(n_323), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_323), .B(n_373), .Y(n_401) );
INVx1_ASAP7_75t_L g359 ( .A(n_325), .Y(n_359) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_327), .B(n_340), .Y(n_432) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_328), .A2(n_446), .B(n_448), .Y(n_445) );
OAI21xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_335), .B(n_343), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g389 ( .A(n_334), .Y(n_389) );
INVx1_ASAP7_75t_L g455 ( .A(n_334), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g428 ( .A(n_338), .Y(n_428) );
OR2x2_ASAP7_75t_L g439 ( .A(n_339), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .C(n_348), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_344), .A2(n_405), .B1(n_407), .B2(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_346), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_349), .B(n_353), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_349), .A2(n_412), .B1(n_415), .B2(n_418), .C(n_419), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B(n_356), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g360 ( .A(n_354), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B1(n_362), .B2(n_841), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g443 ( .A(n_365), .B(n_421), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_397), .C(n_424), .D(n_444), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_380), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B1(n_374), .B2(n_375), .C(n_377), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_370), .A2(n_427), .B1(n_449), .B2(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_373), .B(n_416), .Y(n_415) );
NAND2x1_ASAP7_75t_L g460 ( .A(n_373), .B(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_375), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g382 ( .A(n_379), .B(n_383), .Y(n_382) );
OAI21xp33_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_386), .B(n_391), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g410 ( .A(n_396), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g424 ( .A1(n_396), .A2(n_425), .B(n_429), .C(n_435), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_411), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g458 ( .A(n_406), .B(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx3_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp33_ASAP7_75t_R g435 ( .A1(n_436), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g449 ( .A(n_438), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .Y(n_444) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx5_ASAP7_75t_L g471 ( .A(n_465), .Y(n_471) );
INVx5_ASAP7_75t_L g476 ( .A(n_465), .Y(n_476) );
AND2x6_ASAP7_75t_SL g465 ( .A(n_466), .B(n_468), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_468), .B(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx8_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g487 ( .A(n_481), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_481), .B(n_834), .Y(n_833) );
OAI321xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_491), .A3(n_822), .B1(n_827), .B2(n_828), .C(n_829), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_484), .B(n_822), .Y(n_828) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx6_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x6_ASAP7_75t_SL g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g827 ( .A(n_491), .Y(n_827) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_495), .Y(n_498) );
BUFx8_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g835 ( .A(n_496), .B(n_836), .Y(n_835) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_714), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_501), .B(n_656), .Y(n_500) );
NAND3xp33_ASAP7_75t_SL g501 ( .A(n_502), .B(n_593), .C(n_638), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_549), .B(n_570), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_503), .A2(n_594), .B1(n_613), .B2(n_625), .Y(n_593) );
AOI22x1_ASAP7_75t_L g718 ( .A1(n_503), .A2(n_719), .B1(n_723), .B2(n_724), .Y(n_718) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_521), .Y(n_504) );
OR2x2_ASAP7_75t_L g679 ( .A(n_505), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
OR2x2_ASAP7_75t_L g554 ( .A(n_506), .B(n_514), .Y(n_554) );
AND2x2_ASAP7_75t_L g597 ( .A(n_506), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g605 ( .A(n_506), .Y(n_605) );
BUFx2_ASAP7_75t_L g655 ( .A(n_506), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_510), .A2(n_546), .B(n_547), .Y(n_545) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_510), .A2(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
AND2x2_ASAP7_75t_L g600 ( .A(n_514), .B(n_537), .Y(n_600) );
INVx1_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
INVx1_ASAP7_75t_L g612 ( .A(n_514), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_514), .B(n_605), .Y(n_674) );
INVx1_ASAP7_75t_L g695 ( .A(n_514), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_514), .B(n_598), .Y(n_765) );
INVx1_ASAP7_75t_L g658 ( .A(n_521), .Y(n_658) );
OR2x2_ASAP7_75t_L g710 ( .A(n_521), .B(n_674), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_537), .Y(n_521) );
AND2x2_ASAP7_75t_L g555 ( .A(n_522), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g603 ( .A(n_522), .B(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_522), .B(n_552), .Y(n_686) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g598 ( .A(n_523), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_532), .B(n_535), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_528), .B(n_530), .Y(n_525) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_531), .B(n_544), .Y(n_543) );
INVx3_ASAP7_75t_L g552 ( .A(n_537), .Y(n_552) );
INVx1_ASAP7_75t_L g652 ( .A(n_537), .Y(n_652) );
AND2x2_ASAP7_75t_L g654 ( .A(n_537), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g672 ( .A(n_537), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g694 ( .A(n_537), .B(n_695), .Y(n_694) );
NAND2x1p5_ASAP7_75t_SL g705 ( .A(n_537), .B(n_681), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_537), .B(n_612), .Y(n_795) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_545), .B(n_548), .Y(n_539) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_550), .A2(n_734), .B1(n_735), .B2(n_737), .Y(n_733) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_551), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_551), .B(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_L g812 ( .A(n_551), .B(n_670), .Y(n_812) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g611 ( .A(n_552), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_552), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g700 ( .A(n_552), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g651 ( .A(n_553), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g741 ( .A(n_554), .Y(n_741) );
OR2x2_ASAP7_75t_L g815 ( .A(n_554), .B(n_742), .Y(n_815) );
INVx1_ASAP7_75t_L g646 ( .A(n_555), .Y(n_646) );
INVx3_ASAP7_75t_L g650 ( .A(n_556), .Y(n_650) );
BUFx2_ASAP7_75t_L g661 ( .A(n_556), .Y(n_661) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g631 ( .A(n_557), .B(n_582), .Y(n_631) );
INVx2_ASAP7_75t_L g677 ( .A(n_557), .Y(n_677) );
INVx1_ASAP7_75t_L g709 ( .A(n_557), .Y(n_709) );
AND2x2_ASAP7_75t_L g722 ( .A(n_557), .B(n_619), .Y(n_722) );
AND2x2_ASAP7_75t_L g744 ( .A(n_557), .B(n_643), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_565), .B(n_568), .Y(n_559) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g735 ( .A(n_571), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_571), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g760 ( .A(n_571), .B(n_628), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_571), .B(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_582), .Y(n_571) );
INVx2_ASAP7_75t_L g617 ( .A(n_572), .Y(n_617) );
AND2x2_ASAP7_75t_L g644 ( .A(n_572), .B(n_645), .Y(n_644) );
AOI21x1_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B(n_580), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g618 ( .A(n_582), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g637 ( .A(n_582), .Y(n_637) );
INVx2_ASAP7_75t_L g645 ( .A(n_582), .Y(n_645) );
OR2x2_ASAP7_75t_L g665 ( .A(n_582), .B(n_619), .Y(n_665) );
AND2x2_ASAP7_75t_L g676 ( .A(n_582), .B(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B1(n_601), .B2(n_606), .C(n_608), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI32xp33_ASAP7_75t_L g706 ( .A1(n_596), .A2(n_610), .A3(n_707), .B1(n_710), .B2(n_711), .Y(n_706) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g696 ( .A(n_597), .Y(n_696) );
AND2x2_ASAP7_75t_L g732 ( .A(n_597), .B(n_611), .Y(n_732) );
INVx1_ASAP7_75t_L g796 ( .A(n_597), .Y(n_796) );
OR2x2_ASAP7_75t_L g670 ( .A(n_598), .B(n_605), .Y(n_670) );
INVx2_ASAP7_75t_L g681 ( .A(n_598), .Y(n_681) );
BUFx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g820 ( .A(n_600), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g807 ( .A(n_603), .Y(n_807) );
INVx1_ASAP7_75t_L g821 ( .A(n_603), .Y(n_821) );
OR2x2_ASAP7_75t_L g701 ( .A(n_604), .B(n_681), .Y(n_701) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_606), .B(n_701), .Y(n_723) );
INVx1_ASAP7_75t_L g754 ( .A(n_606), .Y(n_754) );
BUFx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g788 ( .A(n_607), .Y(n_788) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2x1_ASAP7_75t_L g757 ( .A(n_609), .B(n_758), .Y(n_757) );
OAI21xp5_ASAP7_75t_SL g779 ( .A1(n_610), .A2(n_780), .B(n_785), .Y(n_779) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
AND2x2_ASAP7_75t_L g689 ( .A(n_615), .B(n_631), .Y(n_689) );
INVxp67_ASAP7_75t_SL g819 ( .A(n_615), .Y(n_819) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g721 ( .A(n_616), .Y(n_721) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g703 ( .A(n_617), .B(n_677), .Y(n_703) );
AND2x2_ASAP7_75t_L g774 ( .A(n_617), .B(n_645), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_618), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g702 ( .A(n_618), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g781 ( .A(n_618), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g630 ( .A(n_619), .Y(n_630) );
INVx2_ASAP7_75t_L g643 ( .A(n_619), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_619), .B(n_634), .Y(n_691) );
AND2x2_ASAP7_75t_L g751 ( .A(n_619), .B(n_645), .Y(n_751) );
NAND2xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_632), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g726 ( .A(n_629), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_629), .B(n_709), .Y(n_801) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g633 ( .A(n_630), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g762 ( .A(n_630), .B(n_677), .Y(n_762) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_636), .Y(n_632) );
OR2x2_ASAP7_75t_L g707 ( .A(n_633), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g664 ( .A(n_634), .Y(n_664) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g690 ( .A(n_637), .B(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_646), .B(n_647), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g653 ( .A(n_641), .B(n_650), .Y(n_653) );
BUFx2_ASAP7_75t_L g671 ( .A(n_641), .Y(n_671) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g682 ( .A(n_642), .Y(n_682) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g697 ( .A(n_644), .B(n_661), .Y(n_697) );
INVx2_ASAP7_75t_L g713 ( .A(n_644), .Y(n_713) );
AND2x2_ASAP7_75t_L g755 ( .A(n_644), .B(n_677), .Y(n_755) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g730 ( .A(n_650), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g777 ( .A(n_651), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g808 ( .A(n_652), .Y(n_808) );
INVx2_ASAP7_75t_L g747 ( .A(n_655), .Y(n_747) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_666), .C(n_683), .D(n_698), .Y(n_656) );
NAND2xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_659), .A2(n_737), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_752) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g734 ( .A(n_663), .Y(n_734) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx2_ASAP7_75t_L g727 ( .A(n_664), .Y(n_727) );
INVx2_ASAP7_75t_L g799 ( .A(n_665), .Y(n_799) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B1(n_672), .B2(n_675), .C1(n_678), .C2(n_682), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g753 ( .A(n_669), .B(n_754), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_669), .A2(n_781), .B(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g792 ( .A(n_670), .B(n_736), .Y(n_792) );
OAI21xp33_ASAP7_75t_SL g766 ( .A1(n_671), .A2(n_692), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g685 ( .A(n_674), .B(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_674), .Y(n_737) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx2_ASAP7_75t_L g736 ( .A(n_677), .Y(n_736) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g742 ( .A(n_681), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_687), .B1(n_692), .B2(n_697), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_689), .A2(n_699), .B1(n_702), .B2(n_704), .C(n_706), .Y(n_698) );
INVx3_ASAP7_75t_R g813 ( .A(n_690), .Y(n_813) );
INVx1_ASAP7_75t_L g731 ( .A(n_691), .Y(n_731) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_694), .Y(n_748) );
INVx1_ASAP7_75t_L g758 ( .A(n_694), .Y(n_758) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_703), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g776 ( .A(n_703), .Y(n_776) );
AND2x2_ASAP7_75t_L g804 ( .A(n_703), .B(n_751), .Y(n_804) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g798 ( .A(n_708), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_770), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_752), .C(n_766), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_728), .C(n_738), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g729 ( .A1(n_719), .A2(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g769 ( .A(n_721), .Y(n_769) );
AND2x2_ASAP7_75t_L g810 ( .A(n_721), .B(n_799), .Y(n_810) );
NAND2x1_ASAP7_75t_L g768 ( .A(n_722), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g790 ( .A(n_727), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g782 ( .A(n_736), .Y(n_782) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_743), .B1(n_745), .B2(n_749), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g778 ( .A(n_742), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_744), .B(n_774), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g817 ( .A(n_750), .Y(n_817) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI22xp33_ASAP7_75t_SL g756 ( .A1(n_757), .A2(n_759), .B1(n_761), .B2(n_763), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_797), .Y(n_770) );
O2A1O1Ixp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_775), .B(n_777), .C(n_779), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_773), .A2(n_787), .B(n_789), .Y(n_786) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
O2A1O1Ixp5_ASAP7_75t_SL g797 ( .A1(n_777), .A2(n_798), .B(n_800), .C(n_802), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_781), .A2(n_786), .B1(n_791), .B2(n_793), .Y(n_785) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OAI211xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B(n_809), .C(n_816), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_813), .B2(n_814), .Y(n_809) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI21xp5_ASAP7_75t_SL g816 ( .A1(n_817), .A2(n_818), .B(n_820), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx10_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_R g837 ( .A(n_838), .B(n_839), .Y(n_837) );
endmodule