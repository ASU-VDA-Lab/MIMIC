module fake_jpeg_16553_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_41),
.B1(n_29),
.B2(n_43),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_25),
.B1(n_40),
.B2(n_17),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_52),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_25),
.B(n_30),
.C(n_22),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_32),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_59),
.B1(n_57),
.B2(n_56),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_29),
.B1(n_32),
.B2(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_25),
.B1(n_18),
.B2(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_29),
.B1(n_32),
.B2(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_40),
.Y(n_95)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_73),
.B1(n_89),
.B2(n_68),
.Y(n_98)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_30),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_22),
.B(n_21),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_90),
.B1(n_96),
.B2(n_57),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_0),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_91),
.B1(n_97),
.B2(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_31),
.B1(n_28),
.B2(n_19),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_99),
.B1(n_69),
.B2(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_108),
.B1(n_122),
.B2(n_93),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_47),
.B1(n_62),
.B2(n_67),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_67),
.B1(n_62),
.B2(n_47),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_118),
.B1(n_122),
.B2(n_75),
.Y(n_128)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_47),
.B1(n_58),
.B2(n_65),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_123),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_74),
.B(n_81),
.C(n_85),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_97),
.B(n_19),
.C(n_24),
.D(n_28),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_58),
.B1(n_65),
.B2(n_14),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_83),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_148),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_85),
.B1(n_115),
.B2(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_132),
.B1(n_140),
.B2(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_138),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_96),
.B1(n_90),
.B2(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_137),
.Y(n_158)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_80),
.B(n_78),
.C(n_84),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_93),
.B1(n_88),
.B2(n_92),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_91),
.B1(n_95),
.B2(n_86),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_143),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_89),
.B(n_70),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_70),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_1),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_1),
.B(n_2),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_99),
.A2(n_65),
.B1(n_58),
.B2(n_13),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_127),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_31),
.B1(n_28),
.B2(n_19),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_107),
.C(n_105),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_166),
.C(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_116),
.C(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_104),
.Y(n_171)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_139),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_148),
.B(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_106),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_109),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_149),
.B(n_142),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_203),
.B(n_156),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_129),
.B1(n_145),
.B2(n_133),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_186),
.B1(n_192),
.B2(n_198),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_199),
.B(n_205),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_159),
.B1(n_175),
.B2(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_169),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_166),
.C(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_160),
.B1(n_168),
.B2(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_194),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_145),
.C(n_148),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_128),
.B1(n_148),
.B2(n_136),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_144),
.B(n_147),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_164),
.B(n_169),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_162),
.A2(n_137),
.B1(n_136),
.B2(n_102),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_178),
.B1(n_164),
.B2(n_176),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_206),
.A2(n_209),
.B1(n_217),
.B2(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_213),
.C(n_221),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_153),
.B1(n_170),
.B2(n_161),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_227),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_166),
.C(n_176),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_155),
.B1(n_173),
.B2(n_158),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_155),
.B1(n_137),
.B2(n_152),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_102),
.B1(n_119),
.B2(n_147),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_109),
.C(n_126),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_24),
.C(n_31),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_202),
.C(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_124),
.B1(n_114),
.B2(n_113),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_226),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_24),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_179),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_200),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_242),
.C(n_244),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_203),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_239),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_229),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_185),
.C(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_241),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_221),
.C(n_222),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_206),
.B(n_179),
.CI(n_197),
.CON(n_243),
.SN(n_243)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_243),
.B(n_13),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_183),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_204),
.C(n_188),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_250),
.C(n_252),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_202),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_183),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_204),
.C(n_189),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_212),
.B1(n_218),
.B2(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_231),
.C(n_233),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_227),
.B1(n_220),
.B2(n_180),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_266),
.B1(n_269),
.B2(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_209),
.B1(n_197),
.B2(n_215),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_268),
.B1(n_271),
.B2(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_226),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_228),
.B(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_248),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_236),
.B1(n_239),
.B2(n_238),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_281),
.B(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_282),
.C(n_283),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_277),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_244),
.B(n_234),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_231),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_3),
.C(n_4),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_5),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_285),
.Y(n_295)
);

XOR2x2_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_5),
.Y(n_286)
);

XOR2x1_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_271),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_253),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_293),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_261),
.Y(n_293)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_254),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_267),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_266),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_5),
.B(n_7),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_263),
.B1(n_7),
.B2(n_8),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_256),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_283),
.C(n_282),
.Y(n_303)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_299),
.B(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_294),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_311),
.C(n_312),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_284),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_308),
.B(n_7),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_273),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_9),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_5),
.Y(n_311)
);

AO21x1_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_10),
.B(n_11),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_292),
.B(n_289),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_298),
.B(n_9),
.C(n_10),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_7),
.B(n_9),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_9),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_309),
.B(n_303),
.C(n_311),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_10),
.B(n_11),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_324),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_327),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_326),
.A2(n_318),
.B(n_11),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_323),
.B(n_11),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.C(n_328),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_321),
.B(n_10),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_R g334 ( 
.A(n_333),
.B(n_12),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_12),
.B(n_322),
.Y(n_335)
);


endmodule