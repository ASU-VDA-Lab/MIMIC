module real_aes_17121_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_1404;
wire n_402;
wire n_733;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_0), .A2(n_6), .B1(n_446), .B2(n_981), .Y(n_980) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_0), .A2(n_238), .B1(n_902), .B2(n_1016), .Y(n_1015) );
OAI22xp33_ASAP7_75t_SL g759 ( .A1(n_1), .A2(n_125), .B1(n_619), .B2(n_671), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g772 ( .A1(n_1), .A2(n_31), .B1(n_363), .B2(n_384), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_2), .A2(n_32), .B1(n_401), .B2(n_412), .Y(n_800) );
OAI22xp5_ASAP7_75t_SL g808 ( .A1(n_2), .A2(n_130), .B1(n_363), .B2(n_386), .Y(n_808) );
INVx1_ASAP7_75t_L g1131 ( .A(n_3), .Y(n_1131) );
INVx1_ASAP7_75t_L g688 ( .A(n_4), .Y(n_688) );
INVx1_ASAP7_75t_L g905 ( .A(n_5), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_6), .A2(n_240), .B1(n_350), .B2(n_1016), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_7), .A2(n_257), .B1(n_451), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_7), .A2(n_185), .B1(n_335), .B2(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_8), .A2(n_261), .B1(n_902), .B2(n_955), .Y(n_1078) );
INVxp33_ASAP7_75t_SL g1109 ( .A(n_8), .Y(n_1109) );
OAI211xp5_ASAP7_75t_L g474 ( .A1(n_9), .A2(n_475), .B(n_479), .C(n_480), .Y(n_474) );
INVx1_ASAP7_75t_L g494 ( .A(n_9), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_10), .Y(n_803) );
AOI22xp5_ASAP7_75t_SL g1201 ( .A1(n_11), .A2(n_260), .B1(n_1184), .B2(n_1192), .Y(n_1201) );
INVx1_ASAP7_75t_L g888 ( .A(n_12), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g944 ( .A1(n_13), .A2(n_237), .B1(n_451), .B2(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_13), .A2(n_221), .B1(n_318), .B2(n_966), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g1403 ( .A1(n_14), .A2(n_88), .B1(n_1404), .B2(n_1407), .Y(n_1403) );
OAI22xp33_ASAP7_75t_L g1470 ( .A1(n_14), .A2(n_45), .B1(n_1471), .B2(n_1474), .Y(n_1470) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_15), .Y(n_779) );
INVx1_ASAP7_75t_L g295 ( .A(n_16), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_16), .B(n_305), .Y(n_444) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_16), .B(n_406), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_16), .B(n_228), .Y(n_1402) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_17), .A2(n_206), .B1(n_297), .B2(n_487), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_17), .A2(n_206), .B1(n_626), .B2(n_628), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_18), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_19), .Y(n_717) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_20), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_21), .A2(n_232), .B1(n_451), .B2(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_21), .A2(n_64), .B1(n_353), .B2(n_867), .Y(n_866) );
OAI222xp33_ASAP7_75t_L g822 ( .A1(n_22), .A2(n_209), .B1(n_402), .B2(n_755), .C1(n_823), .C2(n_824), .Y(n_822) );
OAI222xp33_ASAP7_75t_L g853 ( .A1(n_22), .A2(n_147), .B1(n_209), .B2(n_854), .C1(n_855), .C2(n_856), .Y(n_853) );
INVx1_ASAP7_75t_L g500 ( .A(n_23), .Y(n_500) );
INVx1_ASAP7_75t_L g379 ( .A(n_24), .Y(n_379) );
INVx1_ASAP7_75t_L g997 ( .A(n_25), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_25), .A2(n_41), .B1(n_810), .B2(n_855), .Y(n_1007) );
INVx1_ASAP7_75t_L g1002 ( .A(n_26), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1119 ( .A1(n_27), .A2(n_187), .B1(n_297), .B2(n_671), .Y(n_1119) );
OAI22xp33_ASAP7_75t_L g1158 ( .A1(n_27), .A2(n_187), .B1(n_626), .B2(n_650), .Y(n_1158) );
INVx2_ASAP7_75t_L g1179 ( .A(n_28), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_28), .B(n_1180), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_28), .B(n_117), .Y(n_1187) );
OAI22xp33_ASAP7_75t_SL g1125 ( .A1(n_29), .A2(n_30), .B1(n_618), .B2(n_1126), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1162 ( .A1(n_29), .A2(n_30), .B1(n_641), .B2(n_1105), .Y(n_1162) );
OAI22xp33_ASAP7_75t_SL g756 ( .A1(n_31), .A2(n_239), .B1(n_401), .B2(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_32), .B(n_365), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g906 ( .A1(n_33), .A2(n_217), .B1(n_363), .B2(n_907), .Y(n_906) );
OAI22xp33_ASAP7_75t_L g918 ( .A1(n_33), .A2(n_272), .B1(n_401), .B2(n_487), .Y(n_918) );
AOI22xp5_ASAP7_75t_SL g1215 ( .A1(n_34), .A2(n_138), .B1(n_1184), .B2(n_1192), .Y(n_1215) );
INVx1_ASAP7_75t_L g1142 ( .A(n_35), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_36), .A2(n_207), .B1(n_1052), .B2(n_1056), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_36), .A2(n_235), .B1(n_370), .B2(n_966), .Y(n_1064) );
AOI22xp5_ASAP7_75t_SL g1210 ( .A1(n_37), .A2(n_250), .B1(n_1181), .B2(n_1186), .Y(n_1210) );
INVx1_ASAP7_75t_L g838 ( .A(n_38), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_38), .A2(n_232), .B1(n_323), .B2(n_867), .Y(n_873) );
XOR2xp5_ASAP7_75t_L g712 ( .A(n_39), .B(n_713), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_40), .Y(n_789) );
INVx1_ASAP7_75t_L g1000 ( .A(n_41), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_42), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_43), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_44), .A2(n_120), .B1(n_492), .B2(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1114 ( .A(n_44), .Y(n_1114) );
OAI211xp5_ASAP7_75t_L g1390 ( .A1(n_45), .A2(n_1391), .B(n_1396), .C(n_1424), .Y(n_1390) );
INVx1_ASAP7_75t_L g678 ( .A(n_46), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_47), .A2(n_177), .B1(n_1176), .B2(n_1181), .Y(n_1175) );
INVx1_ASAP7_75t_L g1003 ( .A(n_48), .Y(n_1003) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_49), .A2(n_129), .B1(n_411), .B2(n_412), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_49), .A2(n_61), .B1(n_384), .B2(n_386), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_50), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_51), .A2(n_111), .B1(n_1184), .B2(n_1231), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_52), .A2(n_180), .B1(n_384), .B2(n_386), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_52), .A2(n_53), .B1(n_411), .B2(n_412), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_53), .A2(n_277), .B1(n_363), .B2(n_365), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_54), .A2(n_179), .B1(n_1184), .B2(n_1186), .Y(n_1183) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_55), .A2(n_100), .B1(n_1176), .B2(n_1184), .Y(n_1193) );
INVx1_ASAP7_75t_L g927 ( .A(n_56), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_57), .A2(n_90), .B1(n_1052), .B2(n_1054), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_57), .A2(n_102), .B1(n_1063), .B2(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g321 ( .A(n_58), .Y(n_321) );
INVx1_ASAP7_75t_L g329 ( .A(n_58), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_59), .A2(n_137), .B1(n_626), .B2(n_650), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_59), .A2(n_137), .B1(n_297), .B2(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g1034 ( .A(n_60), .Y(n_1034) );
OAI221xp5_ASAP7_75t_L g1043 ( .A1(n_60), .A2(n_116), .B1(n_531), .B2(n_1044), .C(n_1045), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_61), .A2(n_203), .B1(n_401), .B2(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g578 ( .A(n_62), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_63), .Y(n_781) );
INVx1_ASAP7_75t_L g839 ( .A(n_64), .Y(n_839) );
XOR2xp5_ASAP7_75t_L g874 ( .A(n_65), .B(n_875), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_65), .A2(n_270), .B1(n_1176), .B2(n_1181), .Y(n_1195) );
INVx1_ASAP7_75t_L g562 ( .A(n_66), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_67), .A2(n_89), .B1(n_446), .B2(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g1014 ( .A(n_67), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1451 ( .A1(n_68), .A2(n_245), .B1(n_1452), .B2(n_1456), .Y(n_1451) );
INVxp67_ASAP7_75t_SL g1481 ( .A(n_68), .Y(n_1481) );
INVx1_ASAP7_75t_L g288 ( .A(n_69), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_70), .A2(n_225), .B1(n_666), .B2(n_1093), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_70), .A2(n_225), .B1(n_1103), .B2(n_1105), .Y(n_1102) );
INVx2_ASAP7_75t_L g344 ( .A(n_71), .Y(n_344) );
XNOR2x2_ASAP7_75t_L g550 ( .A(n_72), .B(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_73), .A2(n_241), .B1(n_318), .B2(n_323), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_73), .A2(n_183), .B1(n_454), .B2(n_456), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_74), .A2(n_227), .B1(n_618), .B2(n_620), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_74), .A2(n_227), .B1(n_640), .B2(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g880 ( .A(n_75), .Y(n_880) );
INVx1_ASAP7_75t_L g1144 ( .A(n_76), .Y(n_1144) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_77), .A2(n_82), .B1(n_1176), .B2(n_1184), .Y(n_1211) );
INVx1_ASAP7_75t_L g375 ( .A(n_78), .Y(n_375) );
INVx1_ASAP7_75t_L g484 ( .A(n_79), .Y(n_484) );
INVx1_ASAP7_75t_L g369 ( .A(n_80), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g1522 ( .A1(n_81), .A2(n_267), .B1(n_365), .B2(n_386), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1528 ( .A1(n_81), .A2(n_267), .B1(n_411), .B2(n_412), .Y(n_1528) );
INVx1_ASAP7_75t_L g1081 ( .A(n_83), .Y(n_1081) );
INVx1_ASAP7_75t_L g564 ( .A(n_84), .Y(n_564) );
INVx1_ASAP7_75t_L g508 ( .A(n_85), .Y(n_508) );
OAI22xp33_ASAP7_75t_SL g1517 ( .A1(n_86), .A2(n_276), .B1(n_363), .B2(n_384), .Y(n_1517) );
OAI22xp33_ASAP7_75t_L g1524 ( .A1(n_86), .A2(n_276), .B1(n_401), .B2(n_487), .Y(n_1524) );
INVx1_ASAP7_75t_L g993 ( .A(n_87), .Y(n_993) );
OAI221xp5_ASAP7_75t_L g1444 ( .A1(n_88), .A2(n_124), .B1(n_1445), .B2(n_1447), .C(n_1449), .Y(n_1444) );
INVxp67_ASAP7_75t_SL g1018 ( .A(n_89), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_90), .A2(n_192), .B1(n_1061), .B2(n_1063), .Y(n_1060) );
XOR2xp5_ASAP7_75t_L g814 ( .A(n_91), .B(n_815), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_92), .A2(n_274), .B1(n_331), .B2(n_335), .C(n_340), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_92), .A2(n_135), .B1(n_462), .B2(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g1502 ( .A(n_93), .Y(n_1502) );
INVx1_ASAP7_75t_L g1090 ( .A(n_94), .Y(n_1090) );
INVx1_ASAP7_75t_L g752 ( .A(n_95), .Y(n_752) );
OAI211xp5_ASAP7_75t_SL g763 ( .A1(n_95), .A2(n_632), .B(n_764), .C(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g932 ( .A(n_96), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_96), .A2(n_243), .B1(n_719), .B2(n_938), .C(n_939), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_97), .A2(n_162), .B1(n_411), .B2(n_412), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_97), .A2(n_162), .B1(n_365), .B2(n_386), .Y(n_936) );
INVx1_ASAP7_75t_L g998 ( .A(n_98), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g1191 ( .A1(n_99), .A2(n_190), .B1(n_1181), .B2(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1499 ( .A(n_101), .Y(n_1499) );
AOI22xp33_ASAP7_75t_SL g1057 ( .A1(n_102), .A2(n_192), .B1(n_989), .B2(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g556 ( .A(n_103), .Y(n_556) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_104), .A2(n_606), .B(n_609), .C(n_615), .Y(n_605) );
INVx1_ASAP7_75t_L g638 ( .A(n_104), .Y(n_638) );
INVx1_ASAP7_75t_L g1421 ( .A(n_105), .Y(n_1421) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_106), .A2(n_272), .B1(n_365), .B2(n_384), .C(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g916 ( .A(n_106), .Y(n_916) );
INVx1_ASAP7_75t_L g684 ( .A(n_107), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_108), .A2(n_210), .B1(n_411), .B2(n_412), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_108), .A2(n_210), .B1(n_365), .B2(n_386), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_109), .Y(n_290) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_109), .B(n_288), .Y(n_1177) );
OAI211xp5_ASAP7_75t_L g817 ( .A1(n_110), .A2(n_818), .B(n_819), .C(n_828), .Y(n_817) );
INVx1_ASAP7_75t_L g860 ( .A(n_110), .Y(n_860) );
INVx1_ASAP7_75t_L g882 ( .A(n_112), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g950 ( .A1(n_113), .A2(n_221), .B1(n_821), .B2(n_947), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_113), .A2(n_237), .B1(n_955), .B2(n_957), .Y(n_954) );
INVx1_ASAP7_75t_L g1123 ( .A(n_114), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g1233 ( .A1(n_115), .A2(n_163), .B1(n_1176), .B2(n_1181), .Y(n_1233) );
INVx1_ASAP7_75t_L g1485 ( .A(n_115), .Y(n_1485) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_115), .A2(n_1490), .B1(n_1492), .B2(n_1529), .Y(n_1489) );
INVx1_ASAP7_75t_L g1038 ( .A(n_116), .Y(n_1038) );
INVx1_ASAP7_75t_L g1180 ( .A(n_117), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_117), .B(n_1179), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_118), .A2(n_186), .B1(n_1176), .B2(n_1181), .Y(n_1202) );
INVx1_ASAP7_75t_L g883 ( .A(n_119), .Y(n_883) );
INVx1_ASAP7_75t_L g1110 ( .A(n_120), .Y(n_1110) );
INVx2_ASAP7_75t_L g342 ( .A(n_121), .Y(n_342) );
INVx1_ASAP7_75t_L g359 ( .A(n_121), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_121), .B(n_344), .Y(n_1455) );
INVx1_ASAP7_75t_L g516 ( .A(n_122), .Y(n_516) );
INVx1_ASAP7_75t_L g1508 ( .A(n_123), .Y(n_1508) );
INVxp67_ASAP7_75t_SL g1429 ( .A(n_124), .Y(n_1429) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_125), .A2(n_239), .B1(n_365), .B2(n_386), .Y(n_762) );
OAI22xp33_ASAP7_75t_SL g805 ( .A1(n_126), .A2(n_130), .B1(n_411), .B2(n_487), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_126), .A2(n_134), .B1(n_769), .B2(n_770), .Y(n_812) );
XNOR2xp5_ASAP7_75t_L g1116 ( .A(n_127), .B(n_1117), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1422 ( .A1(n_128), .A2(n_142), .B1(n_442), .B2(n_1417), .C(n_1423), .Y(n_1422) );
AOI221xp5_ASAP7_75t_L g1466 ( .A1(n_128), .A2(n_157), .B1(n_869), .B2(n_966), .C(n_1467), .Y(n_1466) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_129), .A2(n_203), .B1(n_363), .B2(n_365), .Y(n_489) );
INVx1_ASAP7_75t_L g693 ( .A(n_131), .Y(n_693) );
INVx1_ASAP7_75t_L g521 ( .A(n_132), .Y(n_521) );
INVx1_ASAP7_75t_L g1419 ( .A(n_133), .Y(n_1419) );
AOI221xp5_ASAP7_75t_L g1459 ( .A1(n_133), .A2(n_279), .B1(n_331), .B2(n_869), .C(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g804 ( .A(n_134), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_135), .A2(n_218), .B1(n_331), .B2(n_335), .C(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g1506 ( .A(n_136), .Y(n_1506) );
INVx1_ASAP7_75t_L g1229 ( .A(n_139), .Y(n_1229) );
INVx1_ASAP7_75t_L g1076 ( .A(n_140), .Y(n_1076) );
INVx1_ASAP7_75t_L g827 ( .A(n_141), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_141), .A2(n_226), .B1(n_365), .B2(n_386), .Y(n_857) );
INVx1_ASAP7_75t_L g1462 ( .A(n_142), .Y(n_1462) );
INVx1_ASAP7_75t_L g518 ( .A(n_143), .Y(n_518) );
AOI31xp33_ASAP7_75t_L g315 ( .A1(n_144), .A2(n_316), .A3(n_361), .B(n_397), .Y(n_315) );
NAND2xp33_ASAP7_75t_SL g439 ( .A(n_144), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_144), .Y(n_468) );
INVx1_ASAP7_75t_L g1028 ( .A(n_145), .Y(n_1028) );
INVx1_ASAP7_75t_L g1137 ( .A(n_146), .Y(n_1137) );
INVx1_ASAP7_75t_L g820 ( .A(n_147), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_148), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g1234 ( .A1(n_149), .A2(n_184), .B1(n_1184), .B2(n_1231), .Y(n_1234) );
INVx1_ASAP7_75t_L g1521 ( .A(n_150), .Y(n_1521) );
OAI211xp5_ASAP7_75t_L g1525 ( .A1(n_150), .A2(n_479), .B(n_512), .C(n_1526), .Y(n_1525) );
BUFx3_ASAP7_75t_L g322 ( .A(n_151), .Y(n_322) );
OAI211xp5_ASAP7_75t_SL g801 ( .A1(n_152), .A2(n_479), .B(n_750), .C(n_802), .Y(n_801) );
OAI211xp5_ASAP7_75t_SL g809 ( .A1(n_152), .A2(n_632), .B(n_810), .C(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g1500 ( .A(n_153), .Y(n_1500) );
INVx1_ASAP7_75t_L g979 ( .A(n_154), .Y(n_979) );
INVx1_ASAP7_75t_L g506 ( .A(n_155), .Y(n_506) );
INVx1_ASAP7_75t_L g676 ( .A(n_156), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g1415 ( .A1(n_157), .A2(n_204), .B1(n_990), .B2(n_1416), .C(n_1417), .Y(n_1415) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_158), .A2(n_254), .B1(n_297), .B2(n_671), .Y(n_1087) );
OAI22xp33_ASAP7_75t_L g1095 ( .A1(n_158), .A2(n_254), .B1(n_650), .B2(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1503 ( .A(n_159), .Y(n_1503) );
CKINVDCx5p33_ASAP7_75t_R g1520 ( .A(n_160), .Y(n_1520) );
INVx1_ASAP7_75t_L g558 ( .A(n_161), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_164), .A2(n_220), .B1(n_1184), .B2(n_1192), .Y(n_1196) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_165), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_166), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_167), .Y(n_834) );
INVx1_ASAP7_75t_L g904 ( .A(n_168), .Y(n_904) );
INVx1_ASAP7_75t_L g1082 ( .A(n_169), .Y(n_1082) );
INVx1_ASAP7_75t_L g1140 ( .A(n_170), .Y(n_1140) );
XOR2x2_ASAP7_75t_L g470 ( .A(n_171), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g682 ( .A(n_172), .Y(n_682) );
INVx1_ASAP7_75t_L g1091 ( .A(n_173), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g1097 ( .A1(n_173), .A2(n_632), .B(n_1098), .C(n_1099), .Y(n_1097) );
INVx1_ASAP7_75t_L g354 ( .A(n_174), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_174), .A2(n_241), .B1(n_446), .B2(n_451), .Y(n_445) );
INVx1_ASAP7_75t_L g571 ( .A(n_175), .Y(n_571) );
INVx1_ASAP7_75t_L g653 ( .A(n_176), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_178), .Y(n_721) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_180), .Y(n_403) );
INVx1_ASAP7_75t_L g994 ( .A(n_181), .Y(n_994) );
INVx1_ASAP7_75t_L g891 ( .A(n_182), .Y(n_891) );
INVx1_ASAP7_75t_L g351 ( .A(n_183), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_185), .A2(n_247), .B1(n_947), .B2(n_949), .Y(n_946) );
INVx1_ASAP7_75t_L g1130 ( .A(n_188), .Y(n_1130) );
INVx1_ASAP7_75t_L g832 ( .A(n_189), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_189), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g523 ( .A(n_191), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_193), .B(n_343), .Y(n_903) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_193), .Y(n_912) );
OAI211xp5_ASAP7_75t_SL g651 ( .A1(n_194), .A2(n_631), .B(n_632), .C(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g664 ( .A(n_194), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_195), .Y(n_734) );
INVx1_ASAP7_75t_L g926 ( .A(n_196), .Y(n_926) );
OAI211xp5_ASAP7_75t_L g749 ( .A1(n_197), .A2(n_479), .B(n_750), .C(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g771 ( .A(n_197), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_198), .A2(n_264), .B1(n_640), .B2(n_641), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_198), .A2(n_264), .B1(n_666), .B2(n_667), .Y(n_665) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_199), .Y(n_301) );
INVx1_ASAP7_75t_L g931 ( .A(n_200), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_201), .Y(n_718) );
INVx1_ASAP7_75t_L g481 ( .A(n_202), .Y(n_481) );
INVx1_ASAP7_75t_L g1461 ( .A(n_204), .Y(n_1461) );
INVx1_ASAP7_75t_L g1425 ( .A(n_205), .Y(n_1425) );
AOI221xp5_ASAP7_75t_L g1067 ( .A1(n_207), .A2(n_262), .B1(n_340), .B2(n_350), .C(n_966), .Y(n_1067) );
INVx1_ASAP7_75t_L g886 ( .A(n_208), .Y(n_886) );
OAI211xp5_ASAP7_75t_L g1088 ( .A1(n_211), .A2(n_658), .B(n_661), .C(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1101 ( .A(n_211), .Y(n_1101) );
XNOR2xp5_ASAP7_75t_L g1493 ( .A(n_212), .B(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1505 ( .A(n_213), .Y(n_1505) );
INVx1_ASAP7_75t_L g614 ( .A(n_214), .Y(n_614) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_214), .A2(n_631), .B(n_632), .C(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g514 ( .A(n_215), .Y(n_514) );
OA22x2_ASAP7_75t_L g922 ( .A1(n_216), .A2(n_923), .B1(n_968), .B2(n_969), .Y(n_922) );
INVxp67_ASAP7_75t_SL g969 ( .A(n_216), .Y(n_969) );
INVxp67_ASAP7_75t_SL g914 ( .A(n_217), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_218), .A2(n_274), .B1(n_454), .B2(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g1124 ( .A(n_219), .Y(n_1124) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_219), .A2(n_631), .B(n_632), .C(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1029 ( .A(n_222), .Y(n_1029) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_223), .Y(n_790) );
XOR2xp5_ASAP7_75t_L g774 ( .A(n_224), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g829 ( .A(n_226), .Y(n_829) );
BUFx3_ASAP7_75t_L g305 ( .A(n_228), .Y(n_305) );
INVx1_ASAP7_75t_L g406 ( .A(n_228), .Y(n_406) );
INVx1_ASAP7_75t_L g611 ( .A(n_229), .Y(n_611) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_230), .B(n_647), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_231), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_233), .Y(n_783) );
INVx1_ASAP7_75t_L g879 ( .A(n_234), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_235), .A2(n_262), .B1(n_465), .B2(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g689 ( .A(n_236), .Y(n_689) );
INVxp67_ASAP7_75t_SL g984 ( .A(n_238), .Y(n_984) );
INVxp67_ASAP7_75t_SL g985 ( .A(n_240), .Y(n_985) );
INVx2_ASAP7_75t_L g346 ( .A(n_242), .Y(n_346) );
INVx1_ASAP7_75t_L g396 ( .A(n_242), .Y(n_396) );
INVx1_ASAP7_75t_L g598 ( .A(n_242), .Y(n_598) );
OAI211xp5_ASAP7_75t_L g929 ( .A1(n_243), .A2(n_430), .B(n_837), .C(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g978 ( .A(n_244), .Y(n_978) );
INVxp67_ASAP7_75t_SL g1432 ( .A(n_245), .Y(n_1432) );
INVx1_ASAP7_75t_L g1509 ( .A(n_246), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_247), .A2(n_257), .B1(n_959), .B2(n_961), .Y(n_958) );
XNOR2x1_ASAP7_75t_L g1070 ( .A(n_248), .B(n_1071), .Y(n_1070) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_249), .A2(n_268), .B1(n_1176), .B2(n_1181), .Y(n_1214) );
XNOR2xp5_ASAP7_75t_L g1024 ( .A(n_251), .B(n_1025), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_252), .Y(n_728) );
XNOR2xp5_ASAP7_75t_L g974 ( .A(n_253), .B(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g1227 ( .A(n_253), .Y(n_1227) );
INVx1_ASAP7_75t_L g1134 ( .A(n_255), .Y(n_1134) );
INVx1_ASAP7_75t_L g890 ( .A(n_256), .Y(n_890) );
INVx1_ASAP7_75t_L g579 ( .A(n_258), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_259), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_261), .Y(n_1113) );
INVx1_ASAP7_75t_L g1077 ( .A(n_263), .Y(n_1077) );
INVx1_ASAP7_75t_L g692 ( .A(n_265), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g843 ( .A1(n_266), .A2(n_454), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g863 ( .A(n_266), .Y(n_863) );
INVx1_ASAP7_75t_L g654 ( .A(n_269), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_269), .A2(n_658), .B(n_661), .C(n_662), .Y(n_657) );
NAND2xp33_ASAP7_75t_SL g1413 ( .A(n_271), .B(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1468 ( .A(n_271), .Y(n_1468) );
OAI211xp5_ASAP7_75t_L g1120 ( .A1(n_273), .A2(n_615), .B(n_1121), .C(n_1122), .Y(n_1120) );
INVx1_ASAP7_75t_L g1161 ( .A(n_273), .Y(n_1161) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_275), .Y(n_825) );
INVx1_ASAP7_75t_L g399 ( .A(n_277), .Y(n_399) );
INVx1_ASAP7_75t_L g569 ( .A(n_278), .Y(n_569) );
INVx1_ASAP7_75t_L g1411 ( .A(n_279), .Y(n_1411) );
OAI211xp5_ASAP7_75t_L g1518 ( .A1(n_280), .A2(n_372), .B(n_1143), .C(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1527 ( .A(n_280), .Y(n_1527) );
INVx1_ASAP7_75t_L g1135 ( .A(n_281), .Y(n_1135) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_306), .B(n_1166), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1488 ( .A(n_285), .B(n_294), .Y(n_1488) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1491 ( .A(n_287), .B(n_290), .Y(n_1491) );
INVx1_ASAP7_75t_L g1533 ( .A(n_287), .Y(n_1533) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g1535 ( .A(n_290), .B(n_1533), .Y(n_1535) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g433 ( .A(n_294), .B(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_SL g816 ( .A1(n_294), .A2(n_817), .B(n_830), .Y(n_816) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g460 ( .A(n_295), .B(n_305), .Y(n_460) );
AND2x4_ASAP7_75t_L g845 ( .A(n_295), .B(n_304), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_296), .A2(n_404), .B1(n_926), .B2(n_927), .Y(n_925) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_296), .A2(n_404), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
AND2x4_ASAP7_75t_SL g1487 ( .A(n_296), .B(n_1488), .Y(n_1487) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
OR2x2_ASAP7_75t_L g411 ( .A(n_298), .B(n_405), .Y(n_411) );
OR2x6_ASAP7_75t_L g619 ( .A(n_298), .B(n_405), .Y(n_619) );
INVx1_ASAP7_75t_L g746 ( .A(n_298), .Y(n_746) );
BUFx4f_ASAP7_75t_L g833 ( .A(n_298), .Y(n_833) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g402 ( .A(n_299), .Y(n_402) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_299), .Y(n_502) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g407 ( .A(n_301), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g416 ( .A(n_301), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_301), .Y(n_423) );
AND2x2_ASAP7_75t_L g429 ( .A(n_301), .B(n_302), .Y(n_429) );
INVx2_ASAP7_75t_L g449 ( .A(n_301), .Y(n_449) );
NAND2x1_ASAP7_75t_L g478 ( .A(n_301), .B(n_302), .Y(n_478) );
INVx2_ASAP7_75t_L g408 ( .A(n_302), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_302), .B(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g420 ( .A(n_302), .Y(n_420) );
INVx1_ASAP7_75t_L g450 ( .A(n_302), .Y(n_450) );
AND2x2_ASAP7_75t_L g452 ( .A(n_302), .B(n_416), .Y(n_452) );
OR2x2_ASAP7_75t_L g511 ( .A(n_302), .B(n_449), .Y(n_511) );
OR2x6_ASAP7_75t_L g401 ( .A(n_303), .B(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_303), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_824) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g413 ( .A(n_304), .Y(n_413) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g421 ( .A(n_305), .B(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g483 ( .A(n_305), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_919), .B2(n_1165), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
XOR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_709), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_548), .B2(n_708), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
XNOR2x1_ASAP7_75t_L g313 ( .A(n_314), .B(n_470), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_436), .Y(n_314) );
INVx1_ASAP7_75t_L g438 ( .A(n_316), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_330), .B(n_347), .Y(n_316) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx3_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
INVx2_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
AND2x4_ASAP7_75t_L g373 ( .A(n_319), .B(n_360), .Y(n_373) );
BUFx2_ASAP7_75t_L g492 ( .A(n_319), .Y(n_492) );
BUFx2_ASAP7_75t_L g867 ( .A(n_319), .Y(n_867) );
BUFx2_ASAP7_75t_L g902 ( .A(n_319), .Y(n_902) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_319), .B(n_1473), .Y(n_1475) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g339 ( .A(n_320), .Y(n_339) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g382 ( .A(n_321), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_321), .B(n_322), .Y(n_388) );
INVx2_ASAP7_75t_L g326 ( .A(n_322), .Y(n_326) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_322), .Y(n_338) );
OR2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_328), .Y(n_364) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx8_ASAP7_75t_L g966 ( .A(n_324), .Y(n_966) );
INVx3_ASAP7_75t_L g1016 ( .A(n_324), .Y(n_1016) );
INVx8_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
BUFx3_ASAP7_75t_L g956 ( .A(n_325), .Y(n_956) );
NAND2x1p5_ASAP7_75t_L g1441 ( .A(n_325), .B(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_325), .B(n_1473), .Y(n_1472) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x4_ASAP7_75t_L g333 ( .A(n_326), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_L g334 ( .A(n_329), .Y(n_334) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g385 ( .A(n_332), .B(n_366), .Y(n_385) );
INVx2_ASAP7_75t_L g540 ( .A(n_332), .Y(n_540) );
AND2x4_ASAP7_75t_L g629 ( .A(n_332), .B(n_366), .Y(n_629) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_332), .Y(n_865) );
INVx2_ASAP7_75t_L g960 ( .A(n_332), .Y(n_960) );
INVx1_ASAP7_75t_L g964 ( .A(n_332), .Y(n_964) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_333), .Y(n_535) );
BUFx8_ASAP7_75t_L g723 ( .A(n_333), .Y(n_723) );
INVx2_ASAP7_75t_L g872 ( .A(n_333), .Y(n_872) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_R g961 ( .A(n_336), .Y(n_961) );
INVx5_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g869 ( .A(n_337), .Y(n_869) );
BUFx12f_ASAP7_75t_L g1063 ( .A(n_337), .Y(n_1063) );
AND2x4_ASAP7_75t_L g1457 ( .A(n_337), .B(n_1454), .Y(n_1457) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
BUFx2_ASAP7_75t_L g378 ( .A(n_338), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_338), .B(n_382), .Y(n_532) );
INVx2_ASAP7_75t_L g770 ( .A(n_338), .Y(n_770) );
INVx1_ASAP7_75t_L g768 ( .A(n_339), .Y(n_768) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI33xp33_ASAP7_75t_L g953 ( .A1(n_341), .A2(n_954), .A3(n_958), .B1(n_962), .B2(n_965), .B3(n_967), .Y(n_953) );
AND3x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .C(n_345), .Y(n_341) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_342), .Y(n_391) );
NAND2xp33_ASAP7_75t_SL g527 ( .A(n_342), .B(n_344), .Y(n_527) );
INVx1_ASAP7_75t_L g1443 ( .A(n_342), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_342), .B(n_343), .Y(n_1469) );
INVx3_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
AND2x2_ASAP7_75t_L g767 ( .A(n_343), .B(n_768), .Y(n_767) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx3_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
INVx1_ASAP7_75t_L g1479 ( .A(n_345), .Y(n_1479) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g357 ( .A(n_346), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_346), .B(n_1402), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_352), .B2(n_354), .C(n_355), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AOI32xp33_ASAP7_75t_L g1059 ( .A1(n_355), .A2(n_1060), .A3(n_1064), .B1(n_1065), .B2(n_1067), .Y(n_1059) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI33xp33_ASAP7_75t_L g877 ( .A1(n_356), .A2(n_674), .A3(n_878), .B1(n_881), .B2(n_884), .B3(n_889), .Y(n_877) );
INVx1_ASAP7_75t_L g967 ( .A(n_356), .Y(n_967) );
OR2x6_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x4_ASAP7_75t_L g443 ( .A(n_357), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g542 ( .A(n_357), .B(n_358), .Y(n_542) );
INVx1_ASAP7_75t_L g849 ( .A(n_357), .Y(n_849) );
INVx3_ASAP7_75t_L g1465 ( .A(n_358), .Y(n_1465) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND3x1_ASAP7_75t_L g596 ( .A(n_359), .B(n_360), .C(n_597), .Y(n_596) );
OR2x4_ASAP7_75t_L g363 ( .A(n_360), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_360), .Y(n_366) );
OR2x6_ASAP7_75t_L g386 ( .A(n_360), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g1442 ( .A(n_360), .B(n_1443), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_361), .B(n_397), .Y(n_437) );
OAI31xp33_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_367), .A3(n_383), .B(n_389), .Y(n_361) );
INVx2_ASAP7_75t_SL g627 ( .A(n_363), .Y(n_627) );
INVx1_ASAP7_75t_L g859 ( .A(n_363), .Y(n_859) );
INVx2_ASAP7_75t_SL g941 ( .A(n_363), .Y(n_941) );
OR2x4_ASAP7_75t_L g365 ( .A(n_364), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g530 ( .A(n_364), .Y(n_530) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_364), .Y(n_544) );
BUFx3_ASAP7_75t_L g585 ( .A(n_364), .Y(n_585) );
BUFx3_ASAP7_75t_L g677 ( .A(n_364), .Y(n_677) );
BUFx3_ASAP7_75t_L g640 ( .A(n_365), .Y(n_640) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_365), .Y(n_1011) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_365), .Y(n_1106) );
NAND3xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_372), .C(n_374), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_369), .A2(n_375), .B1(n_419), .B2(n_421), .Y(n_418) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g957 ( .A(n_371), .Y(n_957) );
INVx2_ASAP7_75t_L g1006 ( .A(n_371), .Y(n_1006) );
NAND3xp33_ASAP7_75t_SL g490 ( .A(n_372), .B(n_491), .C(n_493), .Y(n_490) );
CKINVDCx8_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
CKINVDCx8_ASAP7_75t_R g632 ( .A(n_373), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g852 ( .A(n_373), .B(n_853), .C(n_857), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g935 ( .A(n_373), .B(n_936), .C(n_937), .Y(n_935) );
AOI211xp5_ASAP7_75t_L g1005 ( .A1(n_373), .A2(n_998), .B(n_1006), .C(n_1007), .Y(n_1005) );
NOR3xp33_ASAP7_75t_L g1042 ( .A(n_373), .B(n_1043), .C(n_1046), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_379), .B2(n_380), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_376), .A2(n_380), .B1(n_481), .B2(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_376), .A2(n_767), .B1(n_803), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g855 ( .A(n_376), .Y(n_855) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_376), .A2(n_380), .B1(n_902), .B2(n_903), .C1(n_904), .C2(n_905), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_376), .B(n_931), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_376), .B(n_1033), .Y(n_1045) );
AOI22xp33_ASAP7_75t_SL g1519 ( .A1(n_376), .A2(n_380), .B1(n_1520), .B2(n_1521), .Y(n_1519) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g380 ( .A(n_377), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g635 ( .A(n_377), .B(n_378), .Y(n_635) );
AND2x4_ASAP7_75t_L g637 ( .A(n_377), .B(n_381), .Y(n_637) );
AND2x4_ASAP7_75t_L g765 ( .A(n_377), .B(n_378), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_379), .B(n_425), .Y(n_424) );
AOI32xp33_ASAP7_75t_L g766 ( .A1(n_380), .A2(n_753), .A3(n_767), .B1(n_769), .B2(n_771), .Y(n_766) );
INVxp67_ASAP7_75t_L g810 ( .A(n_380), .Y(n_810) );
INVxp67_ASAP7_75t_L g856 ( .A(n_380), .Y(n_856) );
INVx1_ASAP7_75t_L g1044 ( .A(n_380), .Y(n_1044) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_385), .A2(n_825), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_385), .A2(n_941), .B1(n_1028), .B2(n_1029), .Y(n_1041) );
INVx1_ASAP7_75t_L g642 ( .A(n_386), .Y(n_642) );
INVx2_ASAP7_75t_L g908 ( .A(n_386), .Y(n_908) );
INVx1_ASAP7_75t_L g1104 ( .A(n_386), .Y(n_1104) );
BUFx3_ASAP7_75t_L g593 ( .A(n_387), .Y(n_593) );
INVx1_ASAP7_75t_L g725 ( .A(n_387), .Y(n_725) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g538 ( .A(n_388), .Y(n_538) );
OAI31xp33_ASAP7_75t_SL g488 ( .A1(n_389), .A2(n_489), .A3(n_490), .B(n_495), .Y(n_488) );
INVx1_ASAP7_75t_L g942 ( .A(n_389), .Y(n_942) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
AND2x2_ASAP7_75t_SL g644 ( .A(n_390), .B(n_392), .Y(n_644) );
AND2x2_ASAP7_75t_L g773 ( .A(n_390), .B(n_392), .Y(n_773) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_394), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g526 ( .A(n_394), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g575 ( .A(n_394), .Y(n_575) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AO21x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_409), .B(n_432), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_403), .B2(n_404), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_400), .A2(n_404), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx3_ASAP7_75t_L g577 ( .A(n_402), .Y(n_577) );
BUFx3_ASAP7_75t_L g793 ( .A(n_402), .Y(n_793) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_402), .Y(n_898) );
INVx4_ASAP7_75t_L g487 ( .A(n_404), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g671 ( .A(n_404), .Y(n_671) );
INVx3_ASAP7_75t_SL g818 ( .A(n_404), .Y(n_818) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g917 ( .A(n_412), .Y(n_917) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
AND2x2_ASAP7_75t_L g419 ( .A(n_413), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g431 ( .A(n_413), .B(n_427), .Y(n_431) );
AND2x2_ASAP7_75t_L g616 ( .A(n_413), .B(n_457), .Y(n_616) );
INVx8_ASAP7_75t_L g505 ( .A(n_414), .Y(n_505) );
OR2x2_ASAP7_75t_L g622 ( .A(n_414), .B(n_483), .Y(n_622) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_424), .C(n_430), .Y(n_417) );
INVx1_ASAP7_75t_L g823 ( .A(n_419), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_419), .A2(n_754), .B1(n_931), .B2(n_932), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_419), .A2(n_754), .B1(n_997), .B2(n_998), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_419), .A2(n_421), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
AND2x4_ASAP7_75t_L g482 ( .A(n_420), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g663 ( .A(n_420), .B(n_483), .Y(n_663) );
INVx1_ASAP7_75t_L g1406 ( .A(n_420), .Y(n_1406) );
BUFx3_ASAP7_75t_L g485 ( .A(n_421), .Y(n_485) );
INVx2_ASAP7_75t_L g613 ( .A(n_421), .Y(n_613) );
INVx2_ASAP7_75t_L g755 ( .A(n_421), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_421), .A2(n_663), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_422), .B(n_1402), .Y(n_1408) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_428), .Y(n_1037) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_429), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g995 ( .A(n_430), .B(n_996), .C(n_999), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_430), .B(n_1032), .C(n_1035), .Y(n_1031) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
AO21x1_ASAP7_75t_L g924 ( .A1(n_432), .A2(n_925), .B(n_928), .Y(n_924) );
AOI21xp33_ASAP7_75t_L g991 ( .A1(n_432), .A2(n_992), .B(n_1001), .Y(n_991) );
AO21x1_ASAP7_75t_L g1026 ( .A1(n_432), .A2(n_1027), .B(n_1030), .Y(n_1026) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_433), .A2(n_473), .A3(n_474), .B(n_486), .Y(n_472) );
BUFx3_ASAP7_75t_L g623 ( .A(n_433), .Y(n_623) );
BUFx2_ASAP7_75t_L g760 ( .A(n_433), .Y(n_760) );
OAI31xp33_ASAP7_75t_L g799 ( .A1(n_433), .A2(n_800), .A3(n_801), .B(n_805), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g909 ( .A1(n_433), .A2(n_910), .B(n_918), .Y(n_909) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g1393 ( .A(n_435), .Y(n_1393) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_435), .B(n_1408), .Y(n_1407) );
OAI31xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .A3(n_439), .B(n_467), .Y(n_436) );
INVx1_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
AOI33xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_445), .A3(n_453), .B1(n_458), .B2(n_459), .B3(n_461), .Y(n_440) );
AOI33xp33_ASAP7_75t_L g943 ( .A1(n_441), .A2(n_459), .A3(n_944), .B1(n_946), .B2(n_950), .B3(n_951), .Y(n_943) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_442), .Y(n_1048) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
INVx2_ASAP7_75t_L g554 ( .A(n_443), .Y(n_554) );
INVx2_ASAP7_75t_L g736 ( .A(n_443), .Y(n_736) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g847 ( .A(n_447), .Y(n_847) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_447), .Y(n_1050) );
INVx1_ASAP7_75t_L g1058 ( .A(n_447), .Y(n_1058) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_448), .Y(n_464) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_448), .B(n_1395), .Y(n_1394) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_448), .B(n_1402), .Y(n_1437) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
BUFx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g466 ( .A(n_452), .Y(n_466) );
BUFx6f_ASAP7_75t_L g989 ( .A(n_452), .Y(n_989) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g948 ( .A(n_455), .Y(n_948) );
INVx2_ASAP7_75t_L g1053 ( .A(n_455), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_455), .B(n_1395), .Y(n_1484) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g821 ( .A(n_457), .Y(n_821) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_457), .Y(n_949) );
INVx2_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
INVx2_ASAP7_75t_L g747 ( .A(n_459), .Y(n_747) );
AOI33xp33_ASAP7_75t_L g1047 ( .A1(n_459), .A2(n_1048), .A3(n_1049), .B1(n_1051), .B2(n_1055), .B3(n_1057), .Y(n_1047) );
AND2x4_ASAP7_75t_L g573 ( .A(n_460), .B(n_574), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g836 ( .A1(n_460), .A2(n_699), .B1(n_837), .B2(n_838), .C(n_839), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_460), .B(n_574), .Y(n_990) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g952 ( .A(n_463), .Y(n_952) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g915 ( .A(n_464), .B(n_483), .Y(n_915) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_464), .Y(n_945) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g981 ( .A(n_466), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NAND3xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_488), .C(n_496), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_475), .A2(n_566), .B1(n_1134), .B2(n_1137), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_475), .A2(n_1131), .B1(n_1144), .B2(n_1150), .Y(n_1149) );
INVx5_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_477), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_561) );
BUFx2_ASAP7_75t_SL g570 ( .A(n_477), .Y(n_570) );
BUFx3_ASAP7_75t_L g660 ( .A(n_477), .Y(n_660) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_477), .B(n_1428), .Y(n_1431) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_478), .Y(n_513) );
NAND3xp33_ASAP7_75t_SL g910 ( .A(n_479), .B(n_911), .C(n_913), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_484), .B2(n_485), .Y(n_480) );
BUFx3_ASAP7_75t_L g610 ( .A(n_482), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_482), .A2(n_485), .B1(n_803), .B2(n_804), .Y(n_802) );
O2A1O1Ixp33_ASAP7_75t_L g819 ( .A1(n_483), .A2(n_820), .B(n_821), .C(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g826 ( .A(n_483), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_484), .B(n_492), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g911 ( .A1(n_485), .A2(n_663), .B1(n_821), .B2(n_904), .C1(n_905), .C2(n_912), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_524), .Y(n_496) );
OAI33xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .A3(n_507), .B1(n_515), .B2(n_519), .B3(n_520), .Y(n_497) );
OAI33xp33_ASAP7_75t_L g791 ( .A1(n_498), .A2(n_747), .A3(n_792), .B1(n_794), .B2(n_795), .B3(n_798), .Y(n_791) );
BUFx6f_ASAP7_75t_L g982 ( .A(n_498), .Y(n_982) );
OAI33xp33_ASAP7_75t_L g1145 ( .A1(n_498), .A2(n_572), .A3(n_1146), .B1(n_1148), .B2(n_1149), .B3(n_1152), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_503), .B2(n_506), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_500), .A2(n_516), .B1(n_529), .B2(n_531), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_501), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_501), .A2(n_717), .B1(n_733), .B2(n_738), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g1511 ( .A1(n_501), .A2(n_1156), .B1(n_1502), .B2(n_1505), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g1515 ( .A1(n_501), .A2(n_738), .B1(n_1500), .B2(n_1509), .Y(n_1515) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g557 ( .A(n_502), .Y(n_557) );
BUFx6f_ASAP7_75t_L g1154 ( .A(n_502), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_503), .A2(n_779), .B1(n_789), .B2(n_793), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_503), .A2(n_883), .B1(n_888), .B2(n_898), .Y(n_897) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVxp33_ASAP7_75t_L g1423 ( .A(n_504), .Y(n_1423) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g522 ( .A(n_505), .Y(n_522) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_505), .Y(n_560) );
INVx4_ASAP7_75t_L g738 ( .A(n_505), .Y(n_738) );
INVx1_ASAP7_75t_L g1147 ( .A(n_505), .Y(n_1147) );
INVx1_ASAP7_75t_L g1156 ( .A(n_505), .Y(n_1156) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_506), .A2(n_518), .B1(n_544), .B2(n_545), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_512), .B2(n_514), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_508), .A2(n_521), .B1(n_534), .B2(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_509), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_515) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g563 ( .A(n_510), .Y(n_563) );
BUFx2_ASAP7_75t_L g700 ( .A(n_510), .Y(n_700) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g568 ( .A(n_511), .Y(n_568) );
INVx1_ASAP7_75t_L g741 ( .A(n_511), .Y(n_741) );
BUFx3_ASAP7_75t_L g796 ( .A(n_511), .Y(n_796) );
BUFx2_ASAP7_75t_L g1513 ( .A(n_511), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_512), .A2(n_880), .B1(n_891), .B2(n_896), .Y(n_895) );
OAI221xp5_ASAP7_75t_L g983 ( .A1(n_512), .A2(n_566), .B1(n_984), .B2(n_985), .C(n_986), .Y(n_983) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx4f_ASAP7_75t_L g517 ( .A(n_513), .Y(n_517) );
BUFx4f_ASAP7_75t_L g608 ( .A(n_513), .Y(n_608) );
INVx4_ASAP7_75t_L g702 ( .A(n_513), .Y(n_702) );
BUFx4f_ASAP7_75t_L g750 ( .A(n_513), .Y(n_750) );
BUFx4f_ASAP7_75t_L g842 ( .A(n_513), .Y(n_842) );
OR2x6_ASAP7_75t_L g1398 ( .A(n_513), .B(n_1399), .Y(n_1398) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_514), .A2(n_523), .B1(n_540), .B2(n_541), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_517), .A2(n_740), .B1(n_783), .B2(n_786), .Y(n_794) );
OAI221xp5_ASAP7_75t_L g977 ( .A1(n_517), .A2(n_896), .B1(n_978), .B2(n_979), .C(n_980), .Y(n_977) );
OAI221xp5_ASAP7_75t_L g1418 ( .A1(n_517), .A2(n_1419), .B1(n_1420), .B2(n_1421), .C(n_1422), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1512 ( .A1(n_517), .A2(n_1499), .B1(n_1508), .B2(n_1513), .Y(n_1512) );
OAI33xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_528), .A3(n_533), .B1(n_539), .B2(n_542), .B3(n_543), .Y(n_524) );
OAI33xp33_ASAP7_75t_L g715 ( .A1(n_525), .A2(n_542), .A3(n_716), .B1(n_720), .B2(n_727), .B3(n_732), .Y(n_715) );
OAI33xp33_ASAP7_75t_L g777 ( .A1(n_525), .A2(n_542), .A3(n_778), .B1(n_782), .B2(n_785), .B3(n_788), .Y(n_777) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_525), .Y(n_1079) );
OAI33xp33_ASAP7_75t_L g1128 ( .A1(n_525), .A2(n_594), .A3(n_1129), .B1(n_1133), .B2(n_1136), .B3(n_1141), .Y(n_1128) );
OAI33xp33_ASAP7_75t_L g1497 ( .A1(n_525), .A2(n_542), .A3(n_1498), .B1(n_1501), .B2(n_1504), .B3(n_1507), .Y(n_1497) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx4f_ASAP7_75t_L g581 ( .A(n_526), .Y(n_581) );
BUFx2_ASAP7_75t_L g674 ( .A(n_526), .Y(n_674) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g587 ( .A(n_531), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_531), .A2(n_544), .B1(n_733), .B2(n_734), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_531), .A2(n_544), .B1(n_789), .B2(n_790), .Y(n_788) );
BUFx6f_ASAP7_75t_L g1143 ( .A(n_531), .Y(n_1143) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_531), .A2(n_544), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_532), .Y(n_547) );
BUFx2_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
INVx2_ASAP7_75t_L g687 ( .A(n_534), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_534), .A2(n_728), .B1(n_729), .B2(n_731), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g1498 ( .A1(n_534), .A2(n_541), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx5_ASAP7_75t_L g589 ( .A(n_535), .Y(n_589) );
INVx2_ASAP7_75t_SL g592 ( .A(n_535), .Y(n_592) );
INVx2_ASAP7_75t_SL g1062 ( .A(n_535), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_536), .A2(n_540), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g541 ( .A(n_537), .Y(n_541) );
CKINVDCx8_ASAP7_75t_R g590 ( .A(n_537), .Y(n_590) );
INVx3_ASAP7_75t_L g887 ( .A(n_537), .Y(n_887) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g730 ( .A(n_538), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_540), .A2(n_541), .B1(n_979), .B2(n_1018), .C(n_1019), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_540), .A2(n_593), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_541), .A2(n_592), .B1(n_786), .B2(n_787), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_544), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_544), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g878 ( .A1(n_544), .A2(n_854), .B1(n_879), .B2(n_880), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_544), .A2(n_719), .B1(n_890), .B2(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g1464 ( .A(n_544), .Y(n_1464) );
OAI22xp5_ASAP7_75t_SL g1501 ( .A1(n_544), .A2(n_780), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g631 ( .A(n_546), .Y(n_631) );
INVx2_ASAP7_75t_L g854 ( .A(n_546), .Y(n_854) );
INVx1_ASAP7_75t_L g1098 ( .A(n_546), .Y(n_1098) );
INVx1_ASAP7_75t_L g1132 ( .A(n_546), .Y(n_1132) );
INVx4_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g680 ( .A(n_547), .Y(n_680) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_547), .Y(n_719) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_645), .B(n_707), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g708 ( .A1(n_549), .A2(n_645), .B(n_707), .Y(n_708) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g707 ( .A(n_550), .B(n_646), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_603), .C(n_624), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_580), .Y(n_552) );
OAI33xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .A3(n_561), .B1(n_565), .B2(n_572), .B3(n_576), .Y(n_553) );
OAI33xp33_ASAP7_75t_L g694 ( .A1(n_554), .A2(n_695), .A3(n_698), .B1(n_703), .B2(n_705), .B3(n_706), .Y(n_694) );
OAI22xp5_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_556), .A2(n_569), .B1(n_583), .B2(n_586), .Y(n_582) );
INVx2_ASAP7_75t_SL g697 ( .A(n_557), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_558), .A2(n_571), .B1(n_583), .B2(n_600), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_559), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_559), .A2(n_676), .B1(n_692), .B2(n_696), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_559), .A2(n_684), .B1(n_689), .B2(n_696), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_559), .A2(n_577), .B1(n_1077), .B2(n_1082), .Y(n_1115) );
INVx6_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx5_ASAP7_75t_L g835 ( .A(n_560), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_562), .A2(n_578), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g1151 ( .A(n_563), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_564), .A2(n_579), .B1(n_592), .B2(n_593), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_566), .A2(n_570), .B1(n_1076), .B2(n_1081), .Y(n_1111) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_573), .Y(n_705) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI33xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .A3(n_588), .B1(n_591), .B2(n_594), .B3(n_599), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_583), .A2(n_1130), .B1(n_1131), .B2(n_1132), .Y(n_1129) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx3_ASAP7_75t_L g683 ( .A(n_589), .Y(n_683) );
INVx8_ASAP7_75t_L g1139 ( .A(n_589), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_590), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g870 ( .A1(n_590), .A2(n_834), .B1(n_841), .B2(n_871), .C(n_873), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g1507 ( .A1(n_592), .A2(n_724), .B1(n_1508), .B2(n_1509), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_593), .A2(n_686), .B1(n_688), .B2(n_689), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_593), .A2(n_960), .B1(n_978), .B2(n_1014), .C(n_1015), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_593), .A2(n_1075), .B1(n_1076), .B2(n_1077), .C(n_1078), .Y(n_1074) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_593), .A2(n_864), .B1(n_1081), .B2(n_1082), .C(n_1083), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_593), .A2(n_1137), .B1(n_1138), .B2(n_1140), .Y(n_1136) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_595), .Y(n_690) );
INVx2_ASAP7_75t_L g1085 ( .A(n_595), .Y(n_1085) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g1022 ( .A(n_596), .Y(n_1022) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_598), .B(n_1395), .Y(n_1428) );
INVx1_ASAP7_75t_L g1435 ( .A(n_598), .Y(n_1435) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_600), .A2(n_677), .B1(n_692), .B2(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x6_ASAP7_75t_L g1449 ( .A(n_602), .B(n_1450), .Y(n_1449) );
OAI31xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .A3(n_617), .B(n_623), .Y(n_603) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_612), .B2(n_614), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_610), .A2(n_754), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_611), .A2(n_634), .B1(n_636), .B2(n_638), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_612), .A2(n_653), .B1(n_663), .B2(n_664), .Y(n_662) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g661 ( .A(n_616), .Y(n_661) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g666 ( .A(n_619), .Y(n_666) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g1093 ( .A(n_621), .Y(n_1093) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g669 ( .A(n_622), .Y(n_669) );
INVx1_ASAP7_75t_L g758 ( .A(n_622), .Y(n_758) );
OAI31xp33_ASAP7_75t_L g656 ( .A1(n_623), .A2(n_657), .A3(n_665), .B(n_670), .Y(n_656) );
OAI31xp33_ASAP7_75t_L g1118 ( .A1(n_623), .A2(n_1119), .A3(n_1120), .B(n_1125), .Y(n_1118) );
OAI31xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_630), .A3(n_639), .B(n_643), .Y(n_624) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_627), .A2(n_629), .B1(n_1002), .B2(n_1003), .Y(n_1008) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g650 ( .A(n_629), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_629), .A2(n_926), .B1(n_927), .B2(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_634), .A2(n_636), .B1(n_653), .B2(n_654), .Y(n_652) );
BUFx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_635), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_636), .A2(n_1090), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_636), .A2(n_1100), .B1(n_1123), .B2(n_1161), .Y(n_1160) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g938 ( .A(n_637), .Y(n_938) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI31xp33_ASAP7_75t_L g648 ( .A1(n_643), .A2(n_649), .A3(n_651), .B(n_655), .Y(n_648) );
BUFx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_644), .A2(n_851), .B(n_861), .Y(n_850) );
OAI31xp33_ASAP7_75t_L g1094 ( .A1(n_644), .A2(n_1095), .A3(n_1097), .B(n_1102), .Y(n_1094) );
OAI31xp33_ASAP7_75t_L g1157 ( .A1(n_644), .A2(n_1158), .A3(n_1159), .B(n_1162), .Y(n_1157) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_656), .C(n_672), .Y(n_647) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_660), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_663), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_663), .A2(n_754), .B1(n_1520), .B2(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_668), .A2(n_915), .B1(n_993), .B2(n_994), .C(n_995), .Y(n_992) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g1126 ( .A(n_669), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_694), .Y(n_672) );
OAI33xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .A3(n_681), .B1(n_685), .B2(n_690), .B3(n_691), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_674), .A2(n_690), .B1(n_862), .B2(n_870), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_674), .A2(n_1013), .B1(n_1017), .B2(n_1020), .Y(n_1012) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g1141 ( .A1(n_677), .A2(n_1142), .B1(n_1143), .B2(n_1144), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_678), .A2(n_693), .B1(n_699), .B2(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx3_ASAP7_75t_L g780 ( .A(n_680), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_682), .A2(n_688), .B1(n_699), .B2(n_701), .Y(n_698) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g1146 ( .A1(n_696), .A2(n_1130), .B1(n_1142), .B2(n_1147), .Y(n_1146) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_699), .A2(n_750), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
INVx4_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_702), .Y(n_704) );
INVx2_ASAP7_75t_L g742 ( .A(n_702), .Y(n_742) );
INVx2_ASAP7_75t_L g797 ( .A(n_702), .Y(n_797) );
INVx1_ASAP7_75t_L g837 ( .A(n_702), .Y(n_837) );
OA33x2_ASAP7_75t_L g1107 ( .A1(n_705), .A2(n_982), .A3(n_1108), .B1(n_1111), .B2(n_1112), .B3(n_1115), .Y(n_1107) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
XNOR2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_813), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_774), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_748), .C(n_761), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g714 ( .A(n_715), .B(n_735), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_718), .A2(n_734), .B1(n_740), .B2(n_742), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_724), .B2(n_726), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_721), .A2(n_728), .B1(n_740), .B2(n_742), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g1467 ( .A1(n_722), .A2(n_854), .B1(n_1421), .B2(n_1468), .C(n_1469), .Y(n_1467) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g885 ( .A(n_723), .Y(n_885) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_726), .A2(n_731), .B1(n_738), .B2(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_729), .A2(n_871), .B1(n_882), .B2(n_883), .Y(n_881) );
BUFx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .A3(n_739), .B1(n_743), .B2(n_744), .B3(n_747), .Y(n_735) );
OAI33xp33_ASAP7_75t_L g892 ( .A1(n_736), .A2(n_747), .A3(n_893), .B1(n_894), .B2(n_895), .B3(n_897), .Y(n_892) );
OAI33xp33_ASAP7_75t_L g1510 ( .A1(n_736), .A2(n_747), .A3(n_1511), .B1(n_1512), .B2(n_1514), .B3(n_1515), .Y(n_1510) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_738), .A2(n_784), .B1(n_787), .B2(n_793), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_738), .A2(n_793), .B1(n_879), .B2(n_890), .Y(n_893) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_738), .Y(n_1412) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_740), .A2(n_742), .B1(n_1503), .B2(n_1506), .Y(n_1514) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g896 ( .A(n_741), .Y(n_896) );
INVx1_ASAP7_75t_L g1416 ( .A(n_742), .Y(n_1416) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI31xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_756), .A3(n_759), .B(n_760), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_750), .A2(n_796), .B1(n_882), .B2(n_886), .Y(n_894) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g828 ( .A(n_758), .B(n_829), .Y(n_828) );
OAI31xp33_ASAP7_75t_SL g1086 ( .A1(n_760), .A2(n_1087), .A3(n_1088), .B(n_1092), .Y(n_1086) );
OAI31xp33_ASAP7_75t_SL g1523 ( .A1(n_760), .A2(n_1524), .A3(n_1525), .B(n_1528), .Y(n_1523) );
OAI31xp33_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_763), .A3(n_772), .B(n_773), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_768), .B(n_1442), .Y(n_1448) );
AND2x6_ASAP7_75t_L g1446 ( .A(n_769), .B(n_1442), .Y(n_1446) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI31xp33_ASAP7_75t_SL g806 ( .A1(n_773), .A2(n_807), .A3(n_808), .B(n_809), .Y(n_806) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_773), .A2(n_900), .B(n_906), .Y(n_899) );
OAI31xp33_ASAP7_75t_L g1516 ( .A1(n_773), .A2(n_1517), .A3(n_1518), .B(n_1522), .Y(n_1516) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_799), .C(n_806), .Y(n_775) );
NOR2xp33_ASAP7_75t_SL g776 ( .A(n_777), .B(n_791), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_781), .A2(n_790), .B1(n_796), .B2(n_797), .Y(n_795) );
INVx2_ASAP7_75t_L g1414 ( .A(n_796), .Y(n_1414) );
XOR2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_874), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_848), .B(n_850), .Y(n_815) );
OAI21xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_836), .B(n_840), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_833), .A2(n_835), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
OAI211xp5_ASAP7_75t_SL g840 ( .A1(n_841), .A2(n_842), .B(n_843), .C(n_846), .Y(n_840) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
BUFx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_852), .B(n_858), .Y(n_851) );
OAI221xp5_ASAP7_75t_L g1460 ( .A1(n_854), .A2(n_1461), .B1(n_1462), .B2(n_1463), .C(n_1465), .Y(n_1460) );
OAI211xp5_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_864), .B(n_866), .C(n_868), .Y(n_862) );
INVx2_ASAP7_75t_SL g864 ( .A(n_865), .Y(n_864) );
BUFx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx3_ASAP7_75t_L g1066 ( .A(n_872), .Y(n_1066) );
OR2x6_ASAP7_75t_SL g1452 ( .A(n_872), .B(n_1453), .Y(n_1452) );
NAND3xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_899), .C(n_909), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_892), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_884) );
INVx2_ASAP7_75t_L g1417 ( .A(n_898), .Y(n_1417) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_908), .A2(n_993), .B1(n_994), .B2(n_1010), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_916), .B2(n_917), .Y(n_913) );
INVx1_ASAP7_75t_L g1165 ( .A(n_919), .Y(n_1165) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_1068), .B1(n_1163), .B2(n_1164), .Y(n_919) );
INVx1_ASAP7_75t_L g1164 ( .A(n_920), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_922), .B1(n_970), .B2(n_971), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g968 ( .A(n_923), .Y(n_968) );
NAND4xp75_ASAP7_75t_L g923 ( .A(n_924), .B(n_934), .C(n_943), .D(n_953), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_933), .Y(n_928) );
AO21x1_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_940), .B(n_942), .Y(n_934) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_941), .Y(n_1096) );
AOI31xp33_ASAP7_75t_L g1004 ( .A1(n_942), .A2(n_1005), .A3(n_1008), .B(n_1009), .Y(n_1004) );
AO21x1_ASAP7_75t_L g1040 ( .A1(n_942), .A2(n_1041), .B(n_1042), .Y(n_1040) );
INVx2_ASAP7_75t_SL g947 ( .A(n_948), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_949), .B(n_1000), .Y(n_999) );
BUFx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_966), .Y(n_1084) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
XNOR2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_1023), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NOR4xp25_ASAP7_75t_L g975 ( .A(n_976), .B(n_991), .C(n_1004), .D(n_1012), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_982), .B1(n_983), .B2(n_990), .Y(n_976) );
AND2x4_ASAP7_75t_L g1426 ( .A(n_981), .B(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
NAND4xp75_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1040), .C(n_1047), .D(n_1059), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1039), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1038), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1037), .Y(n_1054) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1037), .Y(n_1056) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1066), .Y(n_1075) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1068), .Y(n_1163) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
XNOR2x1_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1116), .Y(n_1069) );
NAND4xp75_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1086), .C(n_1094), .D(n_1107), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1079), .B1(n_1080), .B2(n_1085), .Y(n_1073) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
AND3x1_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1127), .C(n_1157), .Y(n_1117) );
NOR2xp33_ASAP7_75t_SL g1127 ( .A(n_1128), .B(n_1145), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_1135), .A2(n_1140), .B1(n_1153), .B2(n_1155), .Y(n_1152) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1385), .B1(n_1387), .B2(n_1486), .C(n_1489), .Y(n_1166) );
AND3x1_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1314), .C(n_1350), .Y(n_1167) );
NOR3xp33_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1245), .C(n_1303), .Y(n_1168) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1172), .B1(n_1222), .B2(n_1235), .C(n_1238), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1197), .B1(n_1203), .B2(n_1212), .C(n_1216), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1188), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1173), .B(n_1263), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1298 ( .A(n_1173), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1173), .B(n_1317), .Y(n_1316) );
OAI211xp5_ASAP7_75t_SL g1351 ( .A1(n_1173), .A2(n_1352), .B(n_1355), .C(n_1367), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1173), .B(n_1249), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1382 ( .A(n_1173), .B(n_1383), .Y(n_1382) );
INVx4_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx4_ASAP7_75t_L g1205 ( .A(n_1174), .Y(n_1205) );
NAND2xp5_ASAP7_75t_SL g1220 ( .A(n_1174), .B(n_1221), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1174), .B(n_1221), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1174), .B(n_1306), .Y(n_1305) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_1174), .B(n_1237), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1174), .B(n_1273), .Y(n_1360) );
AND2x4_ASAP7_75t_SL g1174 ( .A(n_1175), .B(n_1183), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
AND2x6_ASAP7_75t_L g1181 ( .A(n_1177), .B(n_1182), .Y(n_1181) );
AND2x6_ASAP7_75t_L g1184 ( .A(n_1177), .B(n_1185), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1177), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1177), .B(n_1187), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1177), .B(n_1178), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1177), .B(n_1187), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1181), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1532 ( .A(n_1182), .Y(n_1532) );
INVxp67_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1189), .B(n_1205), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1194), .Y(n_1189) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1190), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1190), .B(n_1213), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1190), .B(n_1221), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1190), .B(n_1212), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1190), .B(n_1213), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1359 ( .A(n_1190), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1190), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1193), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1194), .B(n_1218), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1194), .B(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1194), .B(n_1271), .Y(n_1295) );
AOI222xp33_ASAP7_75t_L g1381 ( .A1(n_1194), .A2(n_1317), .B1(n_1323), .B2(n_1331), .C1(n_1382), .C2(n_1384), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1195), .B(n_1196), .Y(n_1221) );
OAI321xp33_ASAP7_75t_L g1303 ( .A1(n_1197), .A2(n_1304), .A3(n_1307), .B1(n_1308), .B2(n_1309), .C(n_1310), .Y(n_1303) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1198), .B(n_1232), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1198), .B(n_1205), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g1340 ( .A(n_1198), .B(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1199), .B(n_1208), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1199), .B(n_1209), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1199), .B(n_1240), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1199), .B(n_1250), .Y(n_1257) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1199), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1199), .B(n_1232), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1199), .B(n_1232), .Y(n_1362) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1200), .B(n_1250), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
NOR2xp33_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1206), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1204), .B(n_1236), .Y(n_1259) );
NAND3xp33_ASAP7_75t_L g1266 ( .A(n_1204), .B(n_1264), .C(n_1267), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1204), .B(n_1208), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1204), .B(n_1207), .Y(n_1384) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_1205), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1205), .B(n_1208), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1205), .B(n_1225), .Y(n_1297) );
NAND2x1_ASAP7_75t_L g1374 ( .A(n_1205), .B(n_1375), .Y(n_1374) );
NOR2xp33_ASAP7_75t_L g1216 ( .A(n_1206), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1207), .B(n_1306), .Y(n_1309) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1208), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1208), .B(n_1240), .Y(n_1319) );
OAI31xp33_ASAP7_75t_L g1365 ( .A1(n_1208), .A2(n_1213), .A3(n_1258), .B(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1209), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1212), .B(n_1264), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1212), .B(n_1221), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1212), .B(n_1221), .Y(n_1346) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1213), .B(n_1219), .Y(n_1218) );
NAND2x1p5_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1215), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1220), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1218), .B(n_1270), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1218), .B(n_1264), .Y(n_1318) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1218), .Y(n_1353) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1220), .Y(n_1282) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1221), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1221), .B(n_1370), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1221), .B(n_1277), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1221), .B(n_1370), .Y(n_1383) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
NOR2xp33_ASAP7_75t_SL g1223 ( .A(n_1224), .B(n_1232), .Y(n_1223) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1224), .Y(n_1285) );
A2O1A1Ixp33_ASAP7_75t_L g1291 ( .A1(n_1224), .A2(n_1273), .B(n_1292), .C(n_1294), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1224), .B(n_1239), .Y(n_1372) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
OAI221xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1227), .B1(n_1228), .B2(n_1229), .C(n_1230), .Y(n_1225) );
CKINVDCx20_ASAP7_75t_R g1386 ( .A(n_1228), .Y(n_1386) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1232), .Y(n_1236) );
INVx3_ASAP7_75t_L g1240 ( .A(n_1232), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1235), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
NAND3xp33_ASAP7_75t_L g1366 ( .A(n_1236), .B(n_1243), .C(n_1271), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1241), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1239), .B(n_1271), .C(n_1364), .Y(n_1363) );
CKINVDCx14_ASAP7_75t_R g1239 ( .A(n_1240), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1240), .B(n_1249), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1240), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1240), .B(n_1323), .Y(n_1322) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1244), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND3xp33_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1272), .C(n_1287), .Y(n_1245) );
AOI21xp5_ASAP7_75t_L g1246 ( .A1(n_1247), .A2(n_1255), .B(n_1256), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1251), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1248), .B(n_1280), .Y(n_1279) );
O2A1O1Ixp33_ASAP7_75t_L g1344 ( .A1(n_1248), .A2(n_1345), .B(n_1347), .C(n_1349), .Y(n_1344) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1249), .B(n_1255), .Y(n_1265) );
OAI22xp5_ASAP7_75t_SL g1296 ( .A1(n_1249), .A2(n_1284), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
OAI221xp5_ASAP7_75t_L g1373 ( .A1(n_1249), .A2(n_1374), .B1(n_1376), .B2(n_1377), .C(n_1381), .Y(n_1373) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
AOI222xp33_ASAP7_75t_L g1367 ( .A1(n_1251), .A2(n_1267), .B1(n_1295), .B2(n_1322), .C1(n_1368), .C2(n_1369), .Y(n_1367) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1254), .Y(n_1252) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1253), .Y(n_1290) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1254), .Y(n_1281) );
OAI211xp5_ASAP7_75t_SL g1320 ( .A1(n_1254), .A2(n_1321), .B(n_1324), .C(n_1326), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1254), .B(n_1264), .Y(n_1328) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1255), .Y(n_1349) );
OAI322xp33_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1258), .A3(n_1260), .B1(n_1261), .B2(n_1265), .C1(n_1266), .C2(n_1268), .Y(n_1256) );
CKINVDCx5p33_ASAP7_75t_R g1323 ( .A(n_1257), .Y(n_1323) );
CKINVDCx14_ASAP7_75t_R g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1260), .Y(n_1342) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1264), .B(n_1281), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1264), .B(n_1271), .Y(n_1306) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1271), .B(n_1290), .Y(n_1330) );
A2O1A1Ixp33_ASAP7_75t_R g1272 ( .A1(n_1273), .A2(n_1274), .B(n_1278), .C(n_1283), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1273), .B(n_1325), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1273), .B(n_1294), .Y(n_1338) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1273), .Y(n_1376) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
AOI21xp33_ASAP7_75t_SL g1315 ( .A1(n_1275), .A2(n_1316), .B(n_1319), .Y(n_1315) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1277), .B(n_1290), .Y(n_1289) );
AOI211xp5_ASAP7_75t_L g1355 ( .A1(n_1277), .A2(n_1356), .B(n_1357), .C(n_1365), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1277), .B(n_1282), .Y(n_1380) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
INVx2_ASAP7_75t_L g1308 ( .A(n_1285), .Y(n_1308) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1286), .Y(n_1368) );
AOI222xp33_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1291), .B1(n_1295), .B2(n_1296), .C1(n_1299), .C2(n_1300), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
OAI21xp5_ASAP7_75t_L g1310 ( .A1(n_1295), .A2(n_1311), .B(n_1313), .Y(n_1310) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1295), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1298), .B(n_1299), .Y(n_1325) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1299), .Y(n_1334) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g1331 ( .A(n_1302), .Y(n_1331) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AOI22xp5_ASAP7_75t_L g1350 ( .A1(n_1307), .A2(n_1351), .B1(n_1371), .B2(n_1373), .Y(n_1350) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
OAI31xp33_ASAP7_75t_L g1314 ( .A1(n_1308), .A2(n_1315), .A3(n_1320), .B(n_1332), .Y(n_1314) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_1318), .A2(n_1333), .B1(n_1336), .B2(n_1338), .C(n_1339), .Y(n_1332) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
OAI21xp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1329), .B(n_1331), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1328), .B(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1335), .Y(n_1333) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1338), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1344), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
CKINVDCx14_ASAP7_75t_R g1345 ( .A(n_1346), .Y(n_1345) );
INVxp67_ASAP7_75t_SL g1347 ( .A(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1354), .Y(n_1352) );
OAI21xp33_ASAP7_75t_L g1357 ( .A1(n_1358), .A2(n_1361), .B(n_1363), .Y(n_1357) );
INVxp33_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
CKINVDCx20_ASAP7_75t_R g1385 ( .A(n_1386), .Y(n_1385) );
HB1xp67_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
XOR2x2_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1485), .Y(n_1388) );
NOR2x1_ASAP7_75t_SL g1389 ( .A(n_1390), .B(n_1438), .Y(n_1389) );
INVx3_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
AND2x4_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1394), .Y(n_1392) );
AND2x4_ASAP7_75t_L g1483 ( .A(n_1393), .B(n_1484), .Y(n_1483) );
NOR3xp33_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1403), .C(n_1409), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g1397 ( .A(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
NAND2x2_ASAP7_75t_L g1404 ( .A(n_1400), .B(n_1405), .Y(n_1404) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx2_ASAP7_75t_SL g1405 ( .A(n_1406), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1418), .Y(n_1409) );
OAI211xp5_ASAP7_75t_L g1410 ( .A1(n_1411), .A2(n_1412), .B(n_1413), .C(n_1415), .Y(n_1410) );
INVx3_ASAP7_75t_L g1420 ( .A(n_1414), .Y(n_1420) );
AOI222xp33_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1426), .B1(n_1429), .B2(n_1430), .C1(n_1432), .C2(n_1433), .Y(n_1424) );
AOI211xp5_ASAP7_75t_SL g1439 ( .A1(n_1425), .A2(n_1440), .B(n_1444), .C(n_1451), .Y(n_1439) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
AND2x4_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1436), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
A2O1A1Ixp33_ASAP7_75t_SL g1438 ( .A1(n_1439), .A2(n_1458), .B(n_1476), .C(n_1480), .Y(n_1438) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1442), .Y(n_1450) );
INVx4_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
INVx2_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1455), .Y(n_1473) );
INVx3_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NOR3xp33_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1466), .C(n_1470), .Y(n_1458) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx2_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
BUFx2_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1482), .Y(n_1480) );
HB1xp67_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
HB1xp67_ASAP7_75t_SL g1490 ( .A(n_1491), .Y(n_1490) );
INVxp33_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
HB1xp67_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
AND3x1_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1516), .C(n_1523), .Y(n_1495) );
NOR2xp33_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1510), .Y(n_1496) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
OAI21xp5_ASAP7_75t_L g1531 ( .A1(n_1532), .A2(n_1533), .B(n_1534), .Y(n_1531) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
endmodule