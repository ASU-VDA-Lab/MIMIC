module fake_jpeg_8671_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_22),
.B1(n_27),
.B2(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_27),
.B1(n_22),
.B2(n_31),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_66),
.B1(n_57),
.B2(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_21),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_24),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_32),
.B1(n_25),
.B2(n_29),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_32),
.B1(n_19),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_28),
.B1(n_33),
.B2(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_34),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_73),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_43),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_77),
.B1(n_84),
.B2(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_51),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_30),
.B1(n_33),
.B2(n_20),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_36),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_64),
.B(n_57),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_82),
.Y(n_89)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_14),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_65),
.B1(n_51),
.B2(n_52),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_13),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_95),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_77),
.B1(n_74),
.B2(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_108),
.B1(n_74),
.B2(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_63),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_73),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_58),
.B1(n_33),
.B2(n_43),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_83),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_115),
.B(n_124),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_92),
.B(n_107),
.C(n_103),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_128),
.B(n_120),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_80),
.C(n_87),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_109),
.C(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_122),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_68),
.B(n_67),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_99),
.B(n_33),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_128),
.A3(n_94),
.B1(n_127),
.B2(n_115),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_58),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_73),
.B1(n_82),
.B2(n_33),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_91),
.B1(n_95),
.B2(n_89),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_41),
.C(n_54),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_104),
.C(n_90),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_137),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_126),
.B(n_113),
.C(n_112),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_133),
.B1(n_145),
.B2(n_20),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_91),
.B1(n_89),
.B2(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_94),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_146),
.C(n_112),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_106),
.B(n_101),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_122),
.C(n_33),
.Y(n_156)
);

AOI21x1_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_138),
.B(n_139),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_142),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_20),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_20),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_54),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_124),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_152),
.C(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_125),
.C(n_122),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_122),
.C(n_110),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_159),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_85),
.C(n_50),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_39),
.B1(n_50),
.B2(n_3),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_50),
.C(n_2),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_167),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_131),
.B1(n_138),
.B2(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_171),
.B1(n_174),
.B2(n_152),
.Y(n_180)
);

OAI321xp33_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_135),
.A3(n_138),
.B1(n_136),
.B2(n_5),
.C(n_6),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_85),
.B(n_39),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_1),
.B(n_5),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_85),
.B1(n_50),
.B2(n_3),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_154),
.B1(n_147),
.B2(n_153),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_172),
.B1(n_163),
.B2(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_179),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_147),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_182),
.C(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_185),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_177),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_189),
.B(n_182),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_187),
.A2(n_183),
.B1(n_181),
.B2(n_179),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_188),
.A2(n_171),
.B(n_168),
.C(n_9),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_169),
.B(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_194),
.C(n_7),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_190),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_6),
.B(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_193),
.C(n_10),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_11),
.C(n_198),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_11),
.Y(n_200)
);


endmodule