module fake_jpeg_20403_n_77 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_16),
.C(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_8),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_21),
.B(n_10),
.C(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_31),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_20),
.C(n_19),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_22),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_11),
.B(n_14),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_50),
.B(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_14),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_37),
.B1(n_17),
.B2(n_33),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_56),
.B1(n_13),
.B2(n_19),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_37),
.B1(n_13),
.B2(n_41),
.Y(n_56)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_19),
.B(n_13),
.C(n_9),
.D(n_3),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.C(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_65),
.C(n_56),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.C(n_71),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_65),
.B1(n_5),
.B2(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_0),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_66),
.C(n_29),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_1),
.B(n_2),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_3),
.B(n_4),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_72),
.B1(n_6),
.B2(n_5),
.C(n_29),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_19),
.Y(n_77)
);


endmodule