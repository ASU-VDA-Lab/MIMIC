module real_jpeg_12238_n_8 (n_46, n_5, n_4, n_0, n_1, n_47, n_51, n_2, n_48, n_6, n_50, n_7, n_3, n_49, n_52, n_8);

input n_46;
input n_5;
input n_4;
input n_0;
input n_1;
input n_47;
input n_51;
input n_2;
input n_48;
input n_6;
input n_50;
input n_7;
input n_3;
input n_49;
input n_52;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_16),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_28),
.C(n_38),
.Y(n_27)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g8 ( 
.A(n_5),
.B(n_9),
.CI(n_13),
.CON(n_8),
.SN(n_8)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_22),
.C(n_41),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

A2O1A1Ixp33_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_20),
.B(n_21),
.C(n_43),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_26),
.B(n_27),
.C(n_40),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.C(n_34),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_46),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_47),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_48),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_49),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_50),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_51),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_52),
.Y(n_42)
);


endmodule