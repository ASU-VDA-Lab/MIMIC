module real_aes_18121_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_1404;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1280;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI211xp5_ASAP7_75t_L g1347 ( .A1(n_0), .A2(n_688), .B(n_1279), .C(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1361 ( .A(n_0), .Y(n_1361) );
INVx1_ASAP7_75t_L g548 ( .A(n_1), .Y(n_548) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_1), .A2(n_612), .B(n_614), .C(n_623), .Y(n_611) );
INVx1_ASAP7_75t_L g343 ( .A(n_2), .Y(n_343) );
AND2x2_ASAP7_75t_L g390 ( .A(n_2), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g480 ( .A(n_2), .B(n_236), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_2), .B(n_353), .Y(n_700) );
INVx1_ASAP7_75t_L g1127 ( .A(n_3), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_4), .A2(n_139), .B1(n_666), .B2(n_1269), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1282 ( .A1(n_4), .A2(n_139), .B1(n_684), .B2(n_694), .Y(n_1282) );
OAI22xp33_ASAP7_75t_L g1271 ( .A1(n_5), .A2(n_258), .B1(n_345), .B2(n_880), .Y(n_1271) );
OAI22xp33_ASAP7_75t_L g1277 ( .A1(n_5), .A2(n_258), .B1(n_683), .B2(n_1215), .Y(n_1277) );
INVx1_ASAP7_75t_L g1418 ( .A(n_6), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_7), .A2(n_74), .B1(n_590), .B2(n_591), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_7), .A2(n_20), .B1(n_829), .B2(n_1154), .C(n_1156), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1439 ( .A1(n_8), .A2(n_43), .B1(n_1440), .B2(n_1442), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1449 ( .A1(n_8), .A2(n_43), .B1(n_880), .B2(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g364 ( .A(n_9), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_10), .A2(n_160), .B1(n_600), .B2(n_602), .Y(n_599) );
INVx1_ASAP7_75t_L g615 ( .A(n_10), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_11), .A2(n_198), .B1(n_1519), .B2(n_1533), .Y(n_1545) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_12), .A2(n_25), .B1(n_519), .B2(n_1112), .Y(n_1466) );
INVx1_ASAP7_75t_L g1494 ( .A(n_12), .Y(n_1494) );
OAI211xp5_ASAP7_75t_L g785 ( .A1(n_13), .A2(n_688), .B(n_786), .C(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g799 ( .A(n_13), .Y(n_799) );
INVx1_ASAP7_75t_L g1185 ( .A(n_14), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_15), .A2(n_91), .B1(n_1519), .B2(n_1521), .Y(n_1537) );
INVx1_ASAP7_75t_L g1235 ( .A(n_16), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1634 ( .A1(n_17), .A2(n_319), .B1(n_1511), .B2(n_1516), .Y(n_1634) );
OAI22xp33_ASAP7_75t_L g1397 ( .A1(n_18), .A2(n_152), .B1(n_1214), .B2(n_1215), .Y(n_1397) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_18), .A2(n_152), .B1(n_345), .B2(n_806), .Y(n_1399) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_19), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_20), .A2(n_223), .B1(n_1112), .B2(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g765 ( .A(n_21), .Y(n_765) );
INVx2_ASAP7_75t_L g376 ( .A(n_22), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_23), .A2(n_328), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g514 ( .A(n_23), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g1206 ( .A1(n_24), .A2(n_267), .B1(n_345), .B2(n_676), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_24), .A2(n_267), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
AOI221xp5_ASAP7_75t_L g1478 ( .A1(n_25), .A2(n_42), .B1(n_493), .B2(n_1479), .C(n_1481), .Y(n_1478) );
INVx1_ASAP7_75t_L g1135 ( .A(n_26), .Y(n_1135) );
AOI22xp5_ASAP7_75t_L g1542 ( .A1(n_27), .A2(n_204), .B1(n_1511), .B2(n_1516), .Y(n_1542) );
OA222x2_ASAP7_75t_L g1728 ( .A1(n_28), .A2(n_81), .B1(n_232), .B2(n_1729), .C1(n_1732), .C2(n_1736), .Y(n_1728) );
INVx1_ASAP7_75t_L g1780 ( .A(n_28), .Y(n_1780) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_29), .Y(n_338) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_29), .B(n_336), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_30), .A2(n_184), .B1(n_1519), .B2(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g971 ( .A(n_31), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_32), .A2(n_308), .B1(n_621), .B2(n_622), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_32), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_33), .A2(n_193), .B1(n_1519), .B2(n_1521), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_34), .A2(n_190), .B1(n_460), .B2(n_462), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_34), .A2(n_248), .B1(n_533), .B2(n_535), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_35), .A2(n_200), .B1(n_852), .B2(n_1343), .Y(n_1467) );
INVx1_ASAP7_75t_L g1483 ( .A(n_35), .Y(n_1483) );
INVx1_ASAP7_75t_L g404 ( .A(n_36), .Y(n_404) );
INVx1_ASAP7_75t_L g1419 ( .A(n_37), .Y(n_1419) );
INVx1_ASAP7_75t_L g1192 ( .A(n_38), .Y(n_1192) );
CKINVDCx5p33_ASAP7_75t_R g1018 ( .A(n_39), .Y(n_1018) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_40), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g888 ( .A(n_41), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g1469 ( .A1(n_42), .A2(n_298), .B1(n_1112), .B2(n_1470), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_44), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_44), .A2(n_159), .B1(n_949), .B2(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g897 ( .A(n_45), .Y(n_897) );
INVx1_ASAP7_75t_L g1374 ( .A(n_46), .Y(n_1374) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_47), .A2(n_650), .B(n_653), .C(n_656), .Y(n_649) );
INVx1_ASAP7_75t_L g691 ( .A(n_47), .Y(n_691) );
INVx1_ASAP7_75t_L g1231 ( .A(n_48), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1207 ( .A1(n_49), .A2(n_797), .B(n_874), .C(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1218 ( .A(n_49), .Y(n_1218) );
CKINVDCx5p33_ASAP7_75t_R g1749 ( .A(n_50), .Y(n_1749) );
INVx1_ASAP7_75t_L g1148 ( .A(n_51), .Y(n_1148) );
INVx1_ASAP7_75t_L g584 ( .A(n_52), .Y(n_584) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_52), .A2(n_625), .B(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_53), .A2(n_243), .B1(n_621), .B2(n_1085), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_53), .A2(n_227), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
INVx1_ASAP7_75t_L g1394 ( .A(n_54), .Y(n_1394) );
AOI22xp5_ASAP7_75t_L g1527 ( .A1(n_55), .A2(n_158), .B1(n_1519), .B2(n_1521), .Y(n_1527) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_56), .Y(n_1131) );
INVx1_ASAP7_75t_L g1174 ( .A(n_57), .Y(n_1174) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_58), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g1468 ( .A1(n_59), .A2(n_72), .B1(n_1124), .B2(n_1138), .Y(n_1468) );
INVx1_ASAP7_75t_L g1482 ( .A(n_59), .Y(n_1482) );
INVx1_ASAP7_75t_L g712 ( .A(n_60), .Y(n_712) );
INVx1_ASAP7_75t_L g1370 ( .A(n_61), .Y(n_1370) );
OAI22xp33_ASAP7_75t_SL g1073 ( .A1(n_62), .A2(n_234), .B1(n_722), .B2(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1113 ( .A(n_62), .Y(n_1113) );
INVx1_ASAP7_75t_L g568 ( .A(n_63), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_63), .A2(n_290), .B1(n_608), .B2(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g975 ( .A(n_64), .Y(n_975) );
INVx1_ASAP7_75t_L g1287 ( .A(n_65), .Y(n_1287) );
AOI21xp33_ASAP7_75t_L g837 ( .A1(n_66), .A2(n_457), .B(n_838), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_66), .A2(n_250), .B1(n_852), .B2(n_860), .C(n_862), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_67), .Y(n_1462) );
INVx1_ASAP7_75t_L g1188 ( .A(n_68), .Y(n_1188) );
OAI222xp33_ASAP7_75t_L g814 ( .A1(n_69), .A2(n_79), .B1(n_86), .B2(n_366), .C1(n_815), .C2(n_816), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g1036 ( .A1(n_70), .A2(n_112), .B1(n_345), .B2(n_806), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1050 ( .A1(n_70), .A2(n_112), .B1(n_683), .B2(n_794), .Y(n_1050) );
AOI21xp33_ASAP7_75t_L g487 ( .A1(n_71), .A2(n_488), .B(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_71), .A2(n_190), .B1(n_516), .B2(n_519), .Y(n_515) );
INVx1_ASAP7_75t_L g1498 ( .A(n_72), .Y(n_1498) );
INVx1_ASAP7_75t_L g1254 ( .A(n_73), .Y(n_1254) );
OAI211xp5_ASAP7_75t_L g1258 ( .A1(n_73), .A2(n_574), .B(n_857), .C(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1173 ( .A(n_74), .Y(n_1173) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_75), .A2(n_80), .B1(n_882), .B2(n_883), .Y(n_881) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_75), .A2(n_80), .B1(n_694), .B2(n_931), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_76), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_77), .Y(n_443) );
INVx1_ASAP7_75t_L g1230 ( .A(n_78), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1765 ( .A1(n_81), .A2(n_181), .B1(n_1766), .B2(n_1768), .C(n_1770), .Y(n_1765) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_82), .A2(n_281), .B1(n_673), .B2(n_949), .Y(n_1487) );
INVx1_ASAP7_75t_L g1500 ( .A(n_82), .Y(n_1500) );
INVx1_ASAP7_75t_L g1743 ( .A(n_83), .Y(n_1743) );
AOI22xp33_ASAP7_75t_L g1795 ( .A1(n_83), .A2(n_124), .B1(n_531), .B2(n_533), .Y(n_1795) );
INVx1_ASAP7_75t_L g906 ( .A(n_84), .Y(n_906) );
XOR2x2_ASAP7_75t_L g937 ( .A(n_85), .B(n_938), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_86), .A2(n_325), .B1(n_610), .B2(n_846), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_87), .A2(n_157), .B1(n_802), .B2(n_946), .Y(n_1211) );
OAI22xp33_ASAP7_75t_L g1219 ( .A1(n_87), .A2(n_157), .B1(n_1057), .B2(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g943 ( .A(n_88), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_89), .A2(n_149), .B1(n_462), .B2(n_492), .Y(n_839) );
INVx1_ASAP7_75t_L g854 ( .A(n_89), .Y(n_854) );
XNOR2xp5_ASAP7_75t_L g1221 ( .A(n_90), .B(n_1222), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_92), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_93), .A2(n_303), .B1(n_1138), .B2(n_1140), .Y(n_1137) );
AOI221xp5_ASAP7_75t_L g1170 ( .A1(n_93), .A2(n_197), .B1(n_493), .B2(n_621), .C(n_1171), .Y(n_1170) );
OAI211xp5_ASAP7_75t_L g1272 ( .A1(n_94), .A2(n_650), .B(n_653), .C(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1281 ( .A(n_94), .Y(n_1281) );
INVx1_ASAP7_75t_L g1371 ( .A(n_95), .Y(n_1371) );
AOI22xp5_ASAP7_75t_L g1510 ( .A1(n_96), .A2(n_203), .B1(n_1511), .B2(n_1516), .Y(n_1510) );
OAI22xp33_ASAP7_75t_L g1346 ( .A1(n_97), .A2(n_147), .B1(n_570), .B2(n_794), .Y(n_1346) );
OAI22xp33_ASAP7_75t_L g1355 ( .A1(n_97), .A2(n_147), .B1(n_345), .B2(n_676), .Y(n_1355) );
INVx1_ASAP7_75t_L g1501 ( .A(n_98), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_99), .A2(n_138), .B1(n_879), .B2(n_880), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_99), .A2(n_138), .B1(n_923), .B2(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g1209 ( .A(n_100), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_101), .A2(n_169), .B1(n_694), .B2(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_101), .A2(n_205), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g1325 ( .A(n_102), .Y(n_1325) );
INVx1_ASAP7_75t_L g598 ( .A(n_103), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_103), .A2(n_238), .B1(n_621), .B2(n_622), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_104), .Y(n_437) );
INVx1_ASAP7_75t_L g336 ( .A(n_105), .Y(n_336) );
INVx1_ASAP7_75t_L g761 ( .A(n_106), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g940 ( .A1(n_107), .A2(n_653), .B(n_941), .C(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g957 ( .A(n_107), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_108), .A2(n_326), .B1(n_666), .B2(n_670), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_108), .A2(n_116), .B1(n_683), .B2(n_684), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_109), .A2(n_146), .B1(n_802), .B2(n_946), .Y(n_1255) );
OAI22xp33_ASAP7_75t_L g1261 ( .A1(n_109), .A2(n_146), .B1(n_1220), .B2(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1275 ( .A(n_110), .Y(n_1275) );
OAI211xp5_ASAP7_75t_L g1278 ( .A1(n_110), .A2(n_574), .B(n_1279), .C(n_1280), .Y(n_1278) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_111), .A2(n_143), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_111), .B(n_684), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1475 ( .A(n_113), .Y(n_1475) );
INVx1_ASAP7_75t_L g1335 ( .A(n_114), .Y(n_1335) );
INVx1_ASAP7_75t_L g1189 ( .A(n_115), .Y(n_1189) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_116), .A2(n_302), .B1(n_345), .B2(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g983 ( .A(n_117), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g1531 ( .A1(n_118), .A2(n_299), .B1(n_1511), .B2(n_1516), .Y(n_1531) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_119), .A2(n_260), .B1(n_589), .B2(n_591), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_119), .A2(n_489), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g1373 ( .A(n_120), .Y(n_1373) );
INVx1_ASAP7_75t_L g1253 ( .A(n_121), .Y(n_1253) );
INVx1_ASAP7_75t_L g1446 ( .A(n_122), .Y(n_1446) );
OAI211xp5_ASAP7_75t_L g1452 ( .A1(n_122), .A2(n_718), .B(n_1357), .C(n_1453), .Y(n_1452) );
OAI211xp5_ASAP7_75t_L g1392 ( .A1(n_123), .A2(n_574), .B(n_786), .C(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1407 ( .A(n_123), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1750 ( .A1(n_124), .A2(n_166), .B1(n_496), .B2(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1226 ( .A(n_125), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1541 ( .A1(n_126), .A2(n_208), .B1(n_1519), .B2(n_1521), .Y(n_1541) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_127), .A2(n_314), .B1(n_802), .B2(n_946), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_127), .A2(n_314), .B1(n_684), .B2(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g1380 ( .A(n_128), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1756 ( .A1(n_129), .A2(n_181), .B1(n_1757), .B2(n_1760), .Y(n_1756) );
INVx1_ASAP7_75t_L g1781 ( .A(n_129), .Y(n_1781) );
INVx1_ASAP7_75t_L g1327 ( .A(n_130), .Y(n_1327) );
INVx1_ASAP7_75t_L g1329 ( .A(n_131), .Y(n_1329) );
OAI211xp5_ASAP7_75t_L g1037 ( .A1(n_132), .A2(n_653), .B(n_1038), .C(n_1040), .Y(n_1037) );
INVx1_ASAP7_75t_L g1055 ( .A(n_132), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_133), .A2(n_173), .B1(n_806), .B2(n_948), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g958 ( .A1(n_133), .A2(n_173), .B1(n_570), .B2(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g1424 ( .A(n_134), .Y(n_1424) );
INVx1_ASAP7_75t_L g900 ( .A(n_135), .Y(n_900) );
INVx1_ASAP7_75t_L g769 ( .A(n_136), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g1546 ( .A1(n_137), .A2(n_217), .B1(n_1511), .B2(n_1516), .Y(n_1546) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_140), .A2(n_310), .B1(n_941), .B2(n_1089), .C(n_1090), .Y(n_1088) );
INVx1_ASAP7_75t_L g1108 ( .A(n_140), .Y(n_1108) );
INVx1_ASAP7_75t_L g1077 ( .A(n_141), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_141), .A2(n_243), .B1(n_1098), .B2(n_1104), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_142), .Y(n_1081) );
INVx1_ASAP7_75t_L g1111 ( .A(n_143), .Y(n_1111) );
INVx1_ASAP7_75t_L g792 ( .A(n_144), .Y(n_792) );
OAI211xp5_ASAP7_75t_SL g796 ( .A1(n_144), .A2(n_653), .B(n_797), .C(n_798), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_145), .A2(n_205), .B1(n_683), .B2(n_784), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_145), .A2(n_169), .B1(n_345), .B2(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g1274 ( .A(n_148), .Y(n_1274) );
INVxp67_ASAP7_75t_SL g863 ( .A(n_149), .Y(n_863) );
INVx1_ASAP7_75t_L g1349 ( .A(n_150), .Y(n_1349) );
INVx1_ASAP7_75t_L g1377 ( .A(n_151), .Y(n_1377) );
INVx1_ASAP7_75t_L g1195 ( .A(n_153), .Y(n_1195) );
INVx1_ASAP7_75t_L g1238 ( .A(n_154), .Y(n_1238) );
INVx1_ASAP7_75t_L g1332 ( .A(n_155), .Y(n_1332) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_156), .A2(n_316), .B1(n_452), .B2(n_454), .C(n_457), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_156), .A2(n_328), .B1(n_529), .B2(n_530), .Y(n_528) );
XOR2x2_ASAP7_75t_L g1411 ( .A(n_158), .B(n_1412), .Y(n_1411) );
INVxp67_ASAP7_75t_SL g1150 ( .A(n_159), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_160), .A2(n_260), .B1(n_621), .B2(n_622), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g1748 ( .A(n_161), .Y(n_1748) );
INVx1_ASAP7_75t_L g1445 ( .A(n_162), .Y(n_1445) );
INVx1_ASAP7_75t_L g1427 ( .A(n_163), .Y(n_1427) );
INVx1_ASAP7_75t_L g1063 ( .A(n_164), .Y(n_1063) );
INVx1_ASAP7_75t_L g706 ( .A(n_165), .Y(n_706) );
INVx1_ASAP7_75t_L g1791 ( .A(n_166), .Y(n_1791) );
XNOR2xp5_ASAP7_75t_L g1178 ( .A(n_167), .B(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g657 ( .A(n_168), .Y(n_657) );
INVx1_ASAP7_75t_L g974 ( .A(n_170), .Y(n_974) );
INVx1_ASAP7_75t_L g1237 ( .A(n_171), .Y(n_1237) );
INVx1_ASAP7_75t_L g944 ( .A(n_172), .Y(n_944) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_172), .A2(n_688), .B(n_954), .C(n_956), .Y(n_953) );
OAI22xp33_ASAP7_75t_L g1396 ( .A1(n_174), .A2(n_318), .B1(n_694), .B2(n_784), .Y(n_1396) );
OAI22xp33_ASAP7_75t_L g1400 ( .A1(n_174), .A2(n_318), .B1(n_666), .B2(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g836 ( .A(n_175), .Y(n_836) );
AOI221x1_ASAP7_75t_SL g851 ( .A1(n_175), .A2(n_246), .B1(n_777), .B2(n_852), .C(n_853), .Y(n_851) );
AOI221x1_ASAP7_75t_SL g1738 ( .A1(n_176), .A2(n_241), .B1(n_1739), .B2(n_1741), .C(n_1742), .Y(n_1738) );
AOI21xp33_ASAP7_75t_L g1793 ( .A1(n_176), .A2(n_743), .B(n_1794), .Y(n_1793) );
AOI21xp33_ASAP7_75t_L g843 ( .A1(n_177), .A2(n_488), .B(n_489), .Y(n_843) );
INVx1_ASAP7_75t_L g864 ( .A(n_177), .Y(n_864) );
INVx2_ASAP7_75t_L g1514 ( .A(n_178), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_178), .B(n_1515), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_178), .B(n_279), .Y(n_1522) );
INVx1_ASAP7_75t_L g717 ( .A(n_179), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g1526 ( .A1(n_180), .A2(n_255), .B1(n_1511), .B2(n_1516), .Y(n_1526) );
OAI22xp33_ASAP7_75t_L g1447 ( .A1(n_182), .A2(n_240), .B1(n_952), .B2(n_1352), .Y(n_1447) );
OAI22xp33_ASAP7_75t_L g1455 ( .A1(n_182), .A2(n_240), .B1(n_802), .B2(n_883), .Y(n_1455) );
INVx1_ASAP7_75t_L g723 ( .A(n_183), .Y(n_723) );
INVx1_ASAP7_75t_L g876 ( .A(n_185), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_186), .A2(n_362), .B1(n_541), .B2(n_542), .Y(n_361) );
INVxp67_ASAP7_75t_L g542 ( .A(n_186), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g1532 ( .A1(n_186), .A2(n_288), .B1(n_1519), .B2(n_1533), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g1744 ( .A(n_187), .Y(n_1744) );
INVx1_ASAP7_75t_L g732 ( .A(n_188), .Y(n_732) );
OAI211xp5_ASAP7_75t_L g873 ( .A1(n_189), .A2(n_763), .B(n_874), .C(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g929 ( .A(n_189), .Y(n_929) );
XOR2x2_ASAP7_75t_L g1264 ( .A(n_191), .B(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1350 ( .A(n_192), .Y(n_1350) );
OAI211xp5_ASAP7_75t_L g1356 ( .A1(n_192), .A2(n_831), .B(n_1357), .C(n_1360), .Y(n_1356) );
XOR2x2_ASAP7_75t_L g994 ( .A(n_193), .B(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1183 ( .A(n_194), .Y(n_1183) );
OAI221xp5_ASAP7_75t_SL g419 ( .A1(n_195), .A2(n_274), .B1(n_420), .B2(n_428), .C(n_436), .Y(n_419) );
INVx1_ASAP7_75t_L g474 ( .A(n_195), .Y(n_474) );
XOR2xp5_ASAP7_75t_L g1805 ( .A(n_196), .B(n_1806), .Y(n_1805) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_197), .A2(n_285), .B1(n_777), .B2(n_1124), .Y(n_1123) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_198), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g1421 ( .A(n_199), .Y(n_1421) );
INVx1_ASAP7_75t_L g1496 ( .A(n_200), .Y(n_1496) );
INVx1_ASAP7_75t_L g1422 ( .A(n_201), .Y(n_1422) );
INVx2_ASAP7_75t_L g378 ( .A(n_202), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_202), .B(n_376), .Y(n_403) );
INVx1_ASAP7_75t_L g540 ( .A(n_202), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_206), .A2(n_214), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_206), .A2(n_214), .B1(n_784), .B2(n_1057), .Y(n_1056) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_207), .Y(n_1008) );
INVx1_ASAP7_75t_L g791 ( .A(n_209), .Y(n_791) );
INVx1_ASAP7_75t_L g812 ( .A(n_210), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g1536 ( .A1(n_211), .A2(n_296), .B1(n_1511), .B2(n_1516), .Y(n_1536) );
INVx1_ASAP7_75t_L g735 ( .A(n_212), .Y(n_735) );
INVx1_ASAP7_75t_L g768 ( .A(n_213), .Y(n_768) );
OAI22xp33_ASAP7_75t_L g1250 ( .A1(n_215), .A2(n_239), .B1(n_345), .B2(n_676), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_215), .A2(n_239), .B1(n_959), .B2(n_1214), .Y(n_1257) );
BUFx3_ASAP7_75t_L g370 ( .A(n_216), .Y(n_370) );
INVx1_ASAP7_75t_L g384 ( .A(n_218), .Y(n_384) );
INVx1_ASAP7_75t_L g1429 ( .A(n_219), .Y(n_1429) );
INVx1_ASAP7_75t_L g1395 ( .A(n_220), .Y(n_1395) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_220), .A2(n_874), .B(n_1404), .C(n_1406), .Y(n_1403) );
INVx1_ASAP7_75t_L g1191 ( .A(n_221), .Y(n_1191) );
OAI22xp5_ASAP7_75t_SL g824 ( .A1(n_222), .A2(n_261), .B1(n_439), .B2(n_445), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_222), .Y(n_834) );
INVx1_ASAP7_75t_L g1172 ( .A(n_223), .Y(n_1172) );
INVx1_ASAP7_75t_L g966 ( .A(n_224), .Y(n_966) );
INVx1_ASAP7_75t_L g1210 ( .A(n_225), .Y(n_1210) );
OAI211xp5_ASAP7_75t_SL g1216 ( .A1(n_225), .A2(n_688), .B(n_857), .C(n_1217), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_226), .Y(n_1004) );
AOI21xp33_ASAP7_75t_L g1078 ( .A1(n_227), .A2(n_488), .B(n_489), .Y(n_1078) );
INVx1_ASAP7_75t_L g1290 ( .A(n_228), .Y(n_1290) );
INVx1_ASAP7_75t_L g896 ( .A(n_229), .Y(n_896) );
INVx1_ASAP7_75t_L g766 ( .A(n_230), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g1518 ( .A1(n_231), .A2(n_244), .B1(n_1519), .B2(n_1521), .Y(n_1518) );
INVx1_ASAP7_75t_L g1771 ( .A(n_232), .Y(n_1771) );
INVx1_ASAP7_75t_L g561 ( .A(n_233), .Y(n_561) );
INVx1_ASAP7_75t_L g1116 ( .A(n_234), .Y(n_1116) );
INVx1_ASAP7_75t_L g702 ( .A(n_235), .Y(n_702) );
BUFx3_ASAP7_75t_L g353 ( .A(n_236), .Y(n_353) );
INVx1_ASAP7_75t_L g391 ( .A(n_236), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g1351 ( .A1(n_237), .A2(n_283), .B1(n_1262), .B2(n_1352), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_237), .A2(n_283), .B1(n_802), .B2(n_946), .Y(n_1362) );
INVx1_ASAP7_75t_L g587 ( .A(n_238), .Y(n_587) );
INVx1_ASAP7_75t_L g1790 ( .A(n_241), .Y(n_1790) );
INVx1_ASAP7_75t_L g758 ( .A(n_242), .Y(n_758) );
INVx1_ASAP7_75t_L g1726 ( .A(n_244), .Y(n_1726) );
AOI22xp33_ASAP7_75t_L g1800 ( .A1(n_244), .A2(n_1801), .B1(n_1804), .B2(n_1807), .Y(n_1800) );
INVx1_ASAP7_75t_L g759 ( .A(n_245), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_246), .A2(n_250), .B1(n_462), .B2(n_492), .Y(n_844) );
INVx1_ASAP7_75t_L g1296 ( .A(n_247), .Y(n_1296) );
INVx1_ASAP7_75t_L g482 ( .A(n_248), .Y(n_482) );
INVx1_ASAP7_75t_L g877 ( .A(n_249), .Y(n_877) );
OAI211xp5_ASAP7_75t_L g926 ( .A1(n_249), .A2(n_574), .B(n_738), .C(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1233 ( .A(n_251), .Y(n_1233) );
INVx1_ASAP7_75t_L g969 ( .A(n_252), .Y(n_969) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_253), .Y(n_1012) );
INVx1_ASAP7_75t_L g901 ( .A(n_254), .Y(n_901) );
INVx1_ASAP7_75t_L g1295 ( .A(n_256), .Y(n_1295) );
INVx1_ASAP7_75t_L g1333 ( .A(n_257), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g1476 ( .A(n_259), .Y(n_1476) );
INVx1_ASAP7_75t_L g828 ( .A(n_261), .Y(n_828) );
INVx1_ASAP7_75t_L g1292 ( .A(n_262), .Y(n_1292) );
INVx1_ASAP7_75t_L g373 ( .A(n_263), .Y(n_373) );
INVx1_ASAP7_75t_L g435 ( .A(n_263), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_264), .A2(n_544), .B1(n_545), .B2(n_644), .Y(n_543) );
INVxp67_ASAP7_75t_L g644 ( .A(n_264), .Y(n_644) );
INVx1_ASAP7_75t_L g1299 ( .A(n_265), .Y(n_1299) );
INVx1_ASAP7_75t_L g1376 ( .A(n_266), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_268), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_269), .Y(n_551) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_269), .A2(n_317), .B1(n_630), .B2(n_631), .C(n_634), .Y(n_629) );
OAI211xp5_ASAP7_75t_L g1251 ( .A1(n_270), .A2(n_797), .B(n_874), .C(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1260 ( .A(n_270), .Y(n_1260) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_271), .Y(n_1006) );
INVx1_ASAP7_75t_L g841 ( .A(n_272), .Y(n_841) );
INVx1_ASAP7_75t_L g1336 ( .A(n_273), .Y(n_1336) );
INVx1_ASAP7_75t_L g498 ( .A(n_274), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_275), .Y(n_565) );
INVx1_ASAP7_75t_L g1425 ( .A(n_276), .Y(n_1425) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_277), .A2(n_870), .B1(n_871), .B2(n_932), .Y(n_869) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_277), .Y(n_932) );
CKINVDCx5p33_ASAP7_75t_R g1472 ( .A(n_278), .Y(n_1472) );
INVx1_ASAP7_75t_L g1515 ( .A(n_279), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_279), .B(n_1514), .Y(n_1520) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_280), .Y(n_1017) );
INVx1_ASAP7_75t_L g1463 ( .A(n_281), .Y(n_1463) );
OAI211xp5_ASAP7_75t_L g1443 ( .A1(n_282), .A2(n_688), .B(n_865), .C(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1454 ( .A(n_282), .Y(n_1454) );
INVx1_ASAP7_75t_L g964 ( .A(n_284), .Y(n_964) );
INVx1_ASAP7_75t_L g1158 ( .A(n_285), .Y(n_1158) );
INVx1_ASAP7_75t_L g725 ( .A(n_286), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_287), .A2(n_322), .B1(n_1511), .B2(n_1516), .Y(n_1552) );
INVx1_ASAP7_75t_L g661 ( .A(n_289), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_289), .A2(n_686), .B(n_688), .C(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g571 ( .A(n_290), .Y(n_571) );
INVx1_ASAP7_75t_L g1087 ( .A(n_291), .Y(n_1087) );
INVx1_ASAP7_75t_L g1045 ( .A(n_292), .Y(n_1045) );
OAI211xp5_ASAP7_75t_L g1051 ( .A1(n_292), .A2(n_688), .B(n_1052), .C(n_1054), .Y(n_1051) );
INVx1_ASAP7_75t_L g1227 ( .A(n_293), .Y(n_1227) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_294), .Y(n_596) );
INVx1_ASAP7_75t_L g1298 ( .A(n_295), .Y(n_1298) );
INVx1_ASAP7_75t_L g762 ( .A(n_297), .Y(n_762) );
AOI211xp5_ASAP7_75t_SL g1491 ( .A1(n_298), .A2(n_1492), .B(n_1493), .C(n_1495), .Y(n_1491) );
AOI21xp5_ASAP7_75t_SL g1082 ( .A1(n_300), .A2(n_488), .B(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1095 ( .A(n_300), .Y(n_1095) );
INVx1_ASAP7_75t_L g1196 ( .A(n_301), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_302), .A2(n_326), .B1(n_693), .B2(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g1157 ( .A(n_303), .Y(n_1157) );
XNOR2xp5_ASAP7_75t_L g1365 ( .A(n_304), .B(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1379 ( .A(n_305), .Y(n_1379) );
INVx1_ASAP7_75t_L g1322 ( .A(n_306), .Y(n_1322) );
XOR2x2_ASAP7_75t_L g1317 ( .A(n_307), .B(n_1318), .Y(n_1317) );
INVxp67_ASAP7_75t_L g1102 ( .A(n_308), .Y(n_1102) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_309), .Y(n_1000) );
INVxp67_ASAP7_75t_SL g1115 ( .A(n_310), .Y(n_1115) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
INVx1_ASAP7_75t_L g891 ( .A(n_312), .Y(n_891) );
INVx1_ASAP7_75t_L g907 ( .A(n_313), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g1762 ( .A(n_315), .Y(n_1762) );
INVx1_ASAP7_75t_L g509 ( .A(n_316), .Y(n_509) );
INVx1_ASAP7_75t_L g555 ( .A(n_317), .Y(n_555) );
INVx1_ASAP7_75t_L g980 ( .A(n_320), .Y(n_980) );
INVx1_ASAP7_75t_L g1293 ( .A(n_321), .Y(n_1293) );
INVx1_ASAP7_75t_L g382 ( .A(n_323), .Y(n_382) );
INVx1_ASAP7_75t_L g424 ( .A(n_323), .Y(n_424) );
INVx2_ASAP7_75t_L g504 ( .A(n_323), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g1763 ( .A(n_324), .Y(n_1763) );
INVx1_ASAP7_75t_L g823 ( .A(n_325), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g1464 ( .A(n_327), .Y(n_1464) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_354), .B(n_1504), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_339), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g1799 ( .A(n_333), .B(n_342), .Y(n_1799) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g1803 ( .A(n_335), .B(n_338), .Y(n_1803) );
INVx1_ASAP7_75t_L g1810 ( .A(n_335), .Y(n_1810) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g1812 ( .A(n_338), .B(n_1810), .Y(n_1812) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g679 ( .A(n_342), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g458 ( .A(n_343), .B(n_352), .Y(n_458) );
AND2x4_ASAP7_75t_L g490 ( .A(n_343), .B(n_353), .Y(n_490) );
INVx1_ASAP7_75t_L g879 ( .A(n_344), .Y(n_879) );
AND2x4_ASAP7_75t_SL g1798 ( .A(n_344), .B(n_1799), .Y(n_1798) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_346), .B(n_351), .Y(n_345) );
OR2x6_ASAP7_75t_L g668 ( .A(n_346), .B(n_669), .Y(n_668) );
BUFx4f_ASAP7_75t_L g979 ( .A(n_346), .Y(n_979) );
INVxp67_ASAP7_75t_L g1324 ( .A(n_346), .Y(n_1324) );
INVx1_ASAP7_75t_L g1390 ( .A(n_346), .Y(n_1390) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx4f_ASAP7_75t_L g705 ( .A(n_347), .Y(n_705) );
INVx3_ASAP7_75t_L g949 ( .A(n_347), .Y(n_949) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
AND2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g456 ( .A(n_349), .B(n_350), .Y(n_456) );
INVx2_ASAP7_75t_L g464 ( .A(n_349), .Y(n_464) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_349), .B(n_350), .Y(n_486) );
INVx1_ASAP7_75t_L g638 ( .A(n_349), .Y(n_638) );
INVx1_ASAP7_75t_L g394 ( .A(n_350), .Y(n_394) );
INVx2_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
AND2x2_ASAP7_75t_L g463 ( .A(n_350), .B(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g473 ( .A(n_350), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_350), .B(n_464), .Y(n_674) );
OR2x2_ASAP7_75t_L g716 ( .A(n_350), .B(n_393), .Y(n_716) );
OR2x6_ASAP7_75t_L g948 ( .A(n_351), .B(n_949), .Y(n_948) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g655 ( .A(n_352), .Y(n_655) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g660 ( .A(n_353), .Y(n_660) );
AND2x4_ASAP7_75t_L g664 ( .A(n_353), .B(n_637), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_1314), .B2(n_1503), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
XNOR2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_934), .Y(n_356) );
XOR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_810), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_645), .B2(n_809), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
XOR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_543), .Y(n_360) );
INVx1_ASAP7_75t_L g541 ( .A(n_362), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_383), .C(n_418), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_364), .A2(n_495), .B1(n_498), .B2(n_499), .Y(n_494) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx5_ASAP7_75t_L g1151 ( .A(n_366), .Y(n_1151) );
OR2x6_ASAP7_75t_L g366 ( .A(n_367), .B(n_379), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_368), .B(n_374), .Y(n_367) );
BUFx3_ASAP7_75t_L g518 ( .A(n_368), .Y(n_518) );
INVx8_ASAP7_75t_L g534 ( .A(n_368), .Y(n_534) );
BUFx3_ASAP7_75t_L g590 ( .A(n_368), .Y(n_590) );
HB1xp67_ASAP7_75t_L g1776 ( .A(n_368), .Y(n_1776) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
AND2x4_ASAP7_75t_L g410 ( .A(n_369), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g398 ( .A(n_370), .B(n_372), .Y(n_398) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_370), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_370), .B(n_435), .Y(n_442) );
AND2x4_ASAP7_75t_L g520 ( .A(n_370), .B(n_434), .Y(n_520) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
AND2x4_ASAP7_75t_L g422 ( .A(n_374), .B(n_423), .Y(n_422) );
AND2x6_ASAP7_75t_L g1767 ( .A(n_374), .B(n_425), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_374), .B(n_432), .Y(n_1769) );
INVx1_ASAP7_75t_L g1773 ( .A(n_374), .Y(n_1773) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
NAND3x1_ASAP7_75t_L g538 ( .A(n_375), .B(n_539), .C(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g550 ( .A(n_375), .Y(n_550) );
OR2x6_ASAP7_75t_L g553 ( .A(n_375), .B(n_513), .Y(n_553) );
OR2x4_ASAP7_75t_L g570 ( .A(n_375), .B(n_398), .Y(n_570) );
AND2x4_ASAP7_75t_L g575 ( .A(n_375), .B(n_520), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g992 ( .A(n_375), .B(n_540), .Y(n_992) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp33_ASAP7_75t_SL g523 ( .A(n_376), .B(n_378), .Y(n_523) );
BUFx3_ASAP7_75t_L g559 ( .A(n_376), .Y(n_559) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_378), .Y(n_578) );
AND3x4_ASAP7_75t_L g867 ( .A(n_378), .B(n_559), .C(n_643), .Y(n_867) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g388 ( .A(n_380), .Y(n_388) );
INVx1_ASAP7_75t_L g680 ( .A(n_380), .Y(n_680) );
OR2x2_ASAP7_75t_L g1760 ( .A(n_380), .B(n_636), .Y(n_1760) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g402 ( .A(n_381), .Y(n_402) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_404), .B2(n_405), .Y(n_383) );
INVxp67_ASAP7_75t_L g815 ( .A(n_385), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_395), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g1761 ( .A1(n_387), .A2(n_413), .B1(n_1762), .B2(n_1763), .Y(n_1761) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AND2x4_ASAP7_75t_L g413 ( .A(n_388), .B(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_389), .Y(n_609) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
AND2x2_ASAP7_75t_L g414 ( .A(n_390), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g495 ( .A(n_390), .B(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_SL g500 ( .A(n_390), .B(n_455), .Y(n_500) );
AND2x4_ASAP7_75t_L g613 ( .A(n_390), .B(n_415), .Y(n_613) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_390), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1735 ( .A(n_390), .B(n_424), .Y(n_1735) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_391), .Y(n_669) );
INVx3_ASAP7_75t_L g461 ( .A(n_392), .Y(n_461) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_392), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_392), .B(n_480), .Y(n_630) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_393), .Y(n_470) );
OR2x6_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_396), .A2(n_702), .B1(n_723), .B2(n_738), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g771 ( .A1(n_396), .A2(n_750), .B1(n_758), .B2(n_765), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_396), .A2(n_686), .B1(n_759), .B2(n_766), .Y(n_781) );
INVx2_ASAP7_75t_SL g890 ( .A(n_396), .Y(n_890) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g856 ( .A(n_397), .Y(n_856) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x4_ASAP7_75t_L g573 ( .A(n_398), .B(n_550), .Y(n_573) );
BUFx4f_ASAP7_75t_L g749 ( .A(n_398), .Y(n_749) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_398), .Y(n_1003) );
BUFx3_ASAP7_75t_L g1184 ( .A(n_398), .Y(n_1184) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g407 ( .A(n_400), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g439 ( .A(n_401), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g445 ( .A(n_401), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g1129 ( .A(n_401), .Y(n_1129) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
OR2x2_ASAP7_75t_L g522 ( .A(n_402), .B(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_402), .Y(n_580) );
INVx1_ASAP7_75t_L g730 ( .A(n_402), .Y(n_730) );
AND2x2_ASAP7_75t_SL g977 ( .A(n_402), .B(n_490), .Y(n_977) );
INVx1_ASAP7_75t_L g1784 ( .A(n_403), .Y(n_1784) );
INVx1_ASAP7_75t_L g816 ( .A(n_405), .Y(n_816) );
NAND2x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_412), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g1101 ( .A(n_408), .Y(n_1101) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g529 ( .A(n_409), .Y(n_529) );
BUFx2_ASAP7_75t_L g595 ( .A(n_409), .Y(n_595) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_410), .Y(n_508) );
BUFx8_ASAP7_75t_L g743 ( .A(n_410), .Y(n_743) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_410), .Y(n_774) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
INVx2_ASAP7_75t_L g1163 ( .A(n_415), .Y(n_1163) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g619 ( .A(n_416), .Y(n_619) );
AND2x4_ASAP7_75t_L g677 ( .A(n_416), .B(n_669), .Y(n_677) );
BUFx3_ASAP7_75t_L g838 ( .A(n_416), .Y(n_838) );
NOR3xp33_ASAP7_75t_SL g418 ( .A(n_419), .B(n_449), .C(n_505), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_421), .A2(n_429), .B1(n_525), .B2(n_1147), .C(n_1148), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g1474 ( .A1(n_421), .A2(n_429), .B1(n_525), .B2(n_1475), .C(n_1476), .Y(n_1474) );
AND2x4_ASAP7_75t_SL g421 ( .A(n_422), .B(n_425), .Y(n_421) );
AND2x4_ASAP7_75t_SL g429 ( .A(n_422), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g525 ( .A(n_422), .B(n_526), .Y(n_525) );
NAND2x1_ASAP7_75t_L g820 ( .A(n_422), .B(n_425), .Y(n_820) );
AND2x4_ASAP7_75t_L g822 ( .A(n_422), .B(n_430), .Y(n_822) );
OR2x2_ASAP7_75t_L g1731 ( .A(n_423), .B(n_630), .Y(n_1731) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g539 ( .A(n_424), .Y(n_539) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_427), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g531 ( .A(n_427), .B(n_433), .Y(n_531) );
BUFx2_ASAP7_75t_L g560 ( .A(n_427), .Y(n_560) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g448 ( .A(n_435), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_443), .B2(n_444), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_437), .B(n_467), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g1130 ( .A1(n_438), .A2(n_444), .B1(n_1131), .B2(n_1132), .C1(n_1134), .C2(n_1135), .Y(n_1130) );
AOI222xp33_ASAP7_75t_L g1461 ( .A1(n_438), .A2(n_444), .B1(n_1132), .B2(n_1462), .C1(n_1463), .C2(n_1464), .Y(n_1461) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_441), .Y(n_586) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g513 ( .A(n_442), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_443), .A2(n_469), .B1(n_471), .B2(n_474), .C(n_475), .Y(n_468) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g687 ( .A(n_446), .Y(n_687) );
INVx4_ASAP7_75t_L g858 ( .A(n_446), .Y(n_858) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_446), .Y(n_894) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g740 ( .A(n_447), .Y(n_740) );
BUFx2_ASAP7_75t_L g789 ( .A(n_447), .Y(n_789) );
BUFx2_ASAP7_75t_L g564 ( .A(n_448), .Y(n_564) );
AOI31xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_481), .A3(n_494), .B(n_501), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_459), .B(n_465), .Y(n_450) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_454), .A2(n_1127), .B1(n_1148), .B2(n_1162), .C(n_1164), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1486 ( .A1(n_454), .A2(n_1162), .B1(n_1472), .B2(n_1476), .C(n_1487), .Y(n_1486) );
BUFx2_ASAP7_75t_L g1741 ( .A(n_454), .Y(n_1741) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x6_ASAP7_75t_L g639 ( .A(n_455), .B(n_480), .Y(n_639) );
AND2x2_ASAP7_75t_L g654 ( .A(n_455), .B(n_655), .Y(n_654) );
BUFx3_ASAP7_75t_L g1492 ( .A(n_455), .Y(n_1492) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g477 ( .A(n_456), .Y(n_477) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g626 ( .A(n_458), .Y(n_626) );
INVx1_ASAP7_75t_L g1083 ( .A(n_458), .Y(n_1083) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_458), .A2(n_842), .B1(n_917), .B2(n_1157), .C(n_1158), .Y(n_1156) );
OAI221xp5_ASAP7_75t_L g1481 ( .A1(n_458), .A2(n_842), .B1(n_1482), .B2(n_1483), .C(n_1484), .Y(n_1481) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g467 ( .A(n_461), .Y(n_467) );
INVx1_ASAP7_75t_L g492 ( .A(n_461), .Y(n_492) );
INVx2_ASAP7_75t_L g1751 ( .A(n_461), .Y(n_1751) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g493 ( .A(n_463), .Y(n_493) );
INVx2_ASAP7_75t_L g497 ( .A(n_463), .Y(n_497) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_463), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_468), .B(n_478), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_469), .A2(n_821), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g1090 ( .A(n_469), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_469), .A2(n_833), .B1(n_1131), .B2(n_1147), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_469), .A2(n_473), .B1(n_1462), .B2(n_1475), .Y(n_1490) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g1089 ( .A(n_471), .Y(n_1089) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_472), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g659 ( .A(n_473), .B(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g833 ( .A(n_473), .Y(n_833) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_473), .B(n_660), .Y(n_1041) );
INVx1_ASAP7_75t_L g1759 ( .A(n_473), .Y(n_1759) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g1359 ( .A(n_477), .Y(n_1359) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g827 ( .A1(n_479), .A2(n_828), .B(n_829), .C(n_830), .Y(n_827) );
A2O1A1Ixp33_ASAP7_75t_SL g1086 ( .A1(n_479), .A2(n_829), .B(n_1087), .C(n_1088), .Y(n_1086) );
A2O1A1Ixp33_ASAP7_75t_L g1488 ( .A1(n_479), .A2(n_621), .B(n_1464), .C(n_1489), .Y(n_1488) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g633 ( .A(n_480), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_480), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_480), .B(n_504), .Y(n_1755) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_487), .C(n_491), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_483), .A2(n_720), .B1(n_765), .B2(n_766), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_483), .A2(n_1029), .B1(n_1188), .B2(n_1191), .Y(n_1200) );
OAI22xp5_ASAP7_75t_L g1244 ( .A1(n_483), .A2(n_1029), .B1(n_1230), .B2(n_1233), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_483), .A2(n_917), .B1(n_1295), .B2(n_1296), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_483), .A2(n_1026), .B1(n_1332), .B2(n_1333), .Y(n_1331) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_483), .A2(n_713), .B1(n_1371), .B2(n_1380), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_483), .A2(n_973), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
INVx5_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g616 ( .A(n_485), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_485), .B(n_1168), .Y(n_1167) );
BUFx2_ASAP7_75t_SL g1202 ( .A(n_485), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_485), .B(n_1490), .Y(n_1489) );
OR2x2_ASAP7_75t_L g1736 ( .A(n_485), .B(n_1735), .Y(n_1736) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_486), .Y(n_652) );
INVx4_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_490), .B(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_490), .B(n_729), .Y(n_1032) );
OAI221xp5_ASAP7_75t_L g1171 ( .A1(n_490), .A2(n_652), .B1(n_722), .B2(n_1172), .C(n_1173), .Y(n_1171) );
OAI21xp33_ASAP7_75t_L g1493 ( .A1(n_490), .A2(n_722), .B(n_1494), .Y(n_1493) );
INVx2_ASAP7_75t_L g610 ( .A(n_495), .Y(n_610) );
AND2x4_ASAP7_75t_L g1733 ( .A(n_496), .B(n_1734), .Y(n_1733) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g1085 ( .A(n_497), .Y(n_1085) );
AOI211xp5_ASAP7_75t_SL g628 ( .A1(n_499), .A2(n_561), .B(n_629), .C(n_639), .Y(n_628) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g848 ( .A(n_500), .Y(n_848) );
OAI31xp67_ASAP7_75t_L g1764 ( .A1(n_501), .A2(n_1765), .A3(n_1774), .B(n_1785), .Y(n_1764) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g699 ( .A(n_503), .B(n_700), .Y(n_699) );
OR2x6_ASAP7_75t_L g991 ( .A(n_503), .B(n_992), .Y(n_991) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g643 ( .A(n_504), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_521), .B(n_524), .C(n_527), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_509), .B1(n_510), .B2(n_514), .C(n_515), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g1437 ( .A1(n_507), .A2(n_585), .B1(n_1422), .B2(n_1429), .Y(n_1437) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g549 ( .A(n_508), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g1007 ( .A(n_508), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g1094 ( .A(n_508), .Y(n_1094) );
BUFx6f_ASAP7_75t_L g1343 ( .A(n_508), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_510), .A2(n_1006), .B1(n_1007), .B2(n_1008), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_510), .A2(n_1329), .B1(n_1336), .B2(n_1342), .Y(n_1341) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g779 ( .A(n_512), .Y(n_779) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g744 ( .A(n_513), .Y(n_744) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g1779 ( .A1(n_519), .A2(n_852), .B1(n_1780), .B2(n_1781), .Y(n_1779) );
BUFx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g526 ( .A(n_520), .Y(n_526) );
INVx2_ASAP7_75t_L g536 ( .A(n_520), .Y(n_536) );
BUFx2_ASAP7_75t_L g566 ( .A(n_520), .Y(n_566) );
BUFx2_ASAP7_75t_L g1104 ( .A(n_520), .Y(n_1104) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_520), .Y(n_1109) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_520), .Y(n_1143) );
OAI33xp33_ASAP7_75t_L g736 ( .A1(n_521), .A2(n_604), .A3(n_737), .B1(n_741), .B2(n_745), .B3(n_747), .Y(n_736) );
OAI33xp33_ASAP7_75t_L g770 ( .A1(n_521), .A2(n_771), .A3(n_772), .B1(n_775), .B2(n_780), .B3(n_781), .Y(n_770) );
OAI33xp33_ASAP7_75t_L g1181 ( .A1(n_521), .A2(n_1013), .A3(n_1182), .B1(n_1187), .B2(n_1190), .B3(n_1194), .Y(n_1181) );
OAI33xp33_ASAP7_75t_L g1300 ( .A1(n_521), .A2(n_604), .A3(n_1301), .B1(n_1304), .B2(n_1305), .B3(n_1308), .Y(n_1300) );
OAI33xp33_ASAP7_75t_L g1368 ( .A1(n_521), .A2(n_604), .A3(n_1369), .B1(n_1372), .B2(n_1375), .B3(n_1378), .Y(n_1368) );
BUFx4f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx4f_ASAP7_75t_L g593 ( .A(n_522), .Y(n_593) );
BUFx2_ASAP7_75t_L g985 ( .A(n_522), .Y(n_985) );
BUFx8_ASAP7_75t_L g998 ( .A(n_522), .Y(n_998) );
BUFx2_ASAP7_75t_L g1794 ( .A(n_523), .Y(n_1794) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_525), .A2(n_537), .B1(n_851), .B2(n_859), .C(n_866), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .C(n_537), .Y(n_527) );
INVx1_ASAP7_75t_L g583 ( .A(n_529), .Y(n_583) );
INVx1_ASAP7_75t_L g1234 ( .A(n_529), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_530), .A2(n_1087), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
BUFx12f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g852 ( .A(n_531), .Y(n_852) );
BUFx3_ASAP7_75t_L g1124 ( .A(n_531), .Y(n_1124) );
INVx5_ASAP7_75t_L g1141 ( .A(n_531), .Y(n_1141) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g1098 ( .A(n_534), .Y(n_1098) );
INVx8_ASAP7_75t_L g1112 ( .A(n_534), .Y(n_1112) );
INVx2_ASAP7_75t_L g1133 ( .A(n_534), .Y(n_1133) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g591 ( .A(n_536), .Y(n_591) );
INVx2_ASAP7_75t_L g1099 ( .A(n_536), .Y(n_1099) );
INVx1_ASAP7_75t_L g1470 ( .A(n_536), .Y(n_1470) );
INVx2_ASAP7_75t_L g604 ( .A(n_537), .Y(n_604) );
INVx2_ASAP7_75t_L g780 ( .A(n_537), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_537), .Y(n_1013) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g904 ( .A(n_538), .Y(n_904) );
OAI33xp33_ASAP7_75t_L g1337 ( .A1(n_538), .A2(n_998), .A3(n_1338), .B1(n_1340), .B2(n_1341), .B3(n_1344), .Y(n_1337) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI211xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_576), .B(n_581), .C(n_605), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_554), .C(n_567), .D(n_574), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_551), .B2(n_552), .Y(n_547) );
INVx1_ASAP7_75t_L g693 ( .A(n_549), .Y(n_693) );
INVx2_ASAP7_75t_L g794 ( .A(n_549), .Y(n_794) );
INVx2_ASAP7_75t_L g925 ( .A(n_549), .Y(n_925) );
INVx1_ASAP7_75t_L g959 ( .A(n_549), .Y(n_959) );
INVx1_ASAP7_75t_L g1215 ( .A(n_549), .Y(n_1215) );
INVxp67_ASAP7_75t_L g1442 ( .A(n_549), .Y(n_1442) );
INVx2_ASAP7_75t_L g952 ( .A(n_552), .Y(n_952) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx3_ASAP7_75t_L g694 ( .A(n_553), .Y(n_694) );
INVx1_ASAP7_75t_L g1058 ( .A(n_553), .Y(n_1058) );
INVx1_ASAP7_75t_L g1263 ( .A(n_553), .Y(n_1263) );
AOI222xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_561), .B2(n_562), .C1(n_565), .C2(n_566), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_556), .A2(n_562), .B1(n_1253), .B2(n_1260), .Y(n_1259) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx3_ASAP7_75t_L g928 ( .A(n_557), .Y(n_928) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x4_ASAP7_75t_L g563 ( .A(n_558), .B(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g690 ( .A(n_558), .B(n_560), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g1106 ( .A1(n_558), .A2(n_1107), .B(n_1110), .C(n_1114), .Y(n_1106) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_562), .A2(n_876), .B1(n_928), .B2(n_929), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_562), .A2(n_928), .B1(n_1209), .B2(n_1218), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_562), .A2(n_928), .B1(n_1274), .B2(n_1281), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_562), .A2(n_928), .B1(n_1394), .B2(n_1395), .Y(n_1393) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_563), .A2(n_657), .B1(n_690), .B2(n_691), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_563), .A2(n_690), .B1(n_791), .B2(n_792), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_563), .A2(n_690), .B1(n_943), .B2(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_563), .A2(n_690), .B1(n_1042), .B2(n_1055), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_563), .A2(n_690), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_563), .A2(n_690), .B1(n_1349), .B2(n_1350), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_563), .A2(n_690), .B1(n_1445), .B2(n_1446), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_565), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g603 ( .A(n_566), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_571), .B2(n_572), .Y(n_567) );
INVx2_ASAP7_75t_L g683 ( .A(n_569), .Y(n_683) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g924 ( .A(n_570), .Y(n_924) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_570), .Y(n_1214) );
INVx1_ASAP7_75t_L g1441 ( .A(n_570), .Y(n_1441) );
INVx2_ASAP7_75t_L g784 ( .A(n_572), .Y(n_784) );
INVx1_ASAP7_75t_L g931 ( .A(n_572), .Y(n_931) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g684 ( .A(n_573), .Y(n_684) );
BUFx2_ASAP7_75t_L g1220 ( .A(n_573), .Y(n_1220) );
BUFx3_ASAP7_75t_L g1352 ( .A(n_573), .Y(n_1352) );
CKINVDCx8_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
CKINVDCx8_ASAP7_75t_R g688 ( .A(n_575), .Y(n_688) );
OAI31xp33_ASAP7_75t_L g1105 ( .A1(n_575), .A2(n_1106), .A3(n_1117), .B(n_1118), .Y(n_1105) );
OAI31xp33_ASAP7_75t_L g782 ( .A1(n_576), .A2(n_783), .A3(n_785), .B(n_793), .Y(n_782) );
OAI31xp33_ASAP7_75t_L g1049 ( .A1(n_576), .A2(n_1050), .A3(n_1051), .B(n_1056), .Y(n_1049) );
CKINVDCx14_ASAP7_75t_R g1283 ( .A(n_576), .Y(n_1283) );
OAI31xp33_ASAP7_75t_L g1391 ( .A1(n_576), .A2(n_1392), .A3(n_1396), .B(n_1397), .Y(n_1391) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
AND2x2_ASAP7_75t_SL g695 ( .A(n_577), .B(n_579), .Y(n_695) );
AND2x2_ASAP7_75t_L g960 ( .A(n_577), .B(n_579), .Y(n_960) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_577), .B(n_579), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_577), .B(n_579), .Y(n_1353) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_592), .B1(n_594), .B2(n_604), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_585), .B2(n_587), .C(n_588), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g1304 ( .A1(n_583), .A2(n_898), .B1(n_1292), .B2(n_1298), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_585), .A2(n_1010), .B1(n_1011), .B2(n_1012), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_585), .A2(n_1093), .B1(n_1095), .B2(n_1096), .C(n_1097), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_585), .A2(n_1081), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_585), .A2(n_773), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_585), .A2(n_1011), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_585), .A2(n_1101), .B1(n_1327), .B2(n_1335), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1788 ( .A1(n_585), .A2(n_1789), .B1(n_1790), .B2(n_1791), .Y(n_1788) );
CKINVDCx8_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g597 ( .A(n_586), .Y(n_597) );
INVx3_ASAP7_75t_L g898 ( .A(n_586), .Y(n_898) );
INVx1_ASAP7_75t_L g988 ( .A(n_586), .Y(n_988) );
INVx3_ASAP7_75t_L g1193 ( .A(n_586), .Y(n_1193) );
BUFx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g601 ( .A(n_590), .Y(n_601) );
OAI33xp33_ASAP7_75t_L g886 ( .A1(n_592), .A2(n_887), .A3(n_895), .B1(n_899), .B2(n_902), .B3(n_905), .Y(n_886) );
OAI22xp33_ASAP7_75t_L g1091 ( .A1(n_592), .A2(n_780), .B1(n_1092), .B2(n_1100), .Y(n_1091) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_598), .C(n_599), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_595), .A2(n_969), .B1(n_980), .B2(n_988), .Y(n_987) );
OAI211xp5_ASAP7_75t_SL g623 ( .A1(n_596), .A2(n_616), .B(n_624), .C(n_627), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_597), .A2(n_717), .B1(n_735), .B2(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_597), .A2(n_971), .B1(n_983), .B2(n_990), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_597), .A2(n_1293), .B1(n_1299), .B2(n_1306), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_597), .A2(n_1421), .B1(n_1427), .B2(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_628), .B(n_640), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B(n_617), .C(n_620), .Y(n_614) );
BUFx2_ASAP7_75t_L g797 ( .A(n_616), .Y(n_797) );
INVx1_ASAP7_75t_L g1039 ( .A(n_616), .Y(n_1039) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g625 ( .A(n_619), .Y(n_625) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_621), .Y(n_829) );
A2O1A1Ixp33_ASAP7_75t_L g1166 ( .A1(n_621), .A2(n_1135), .B(n_1167), .C(n_1169), .Y(n_1166) );
INVx3_ASAP7_75t_L g1480 ( .A(n_621), .Y(n_1480) );
INVx1_ASAP7_75t_L g1155 ( .A(n_622), .Y(n_1155) );
INVx2_ASAP7_75t_L g1740 ( .A(n_625), .Y(n_1740) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g1169 ( .A(n_633), .Y(n_1169) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_641), .Y(n_849) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_642), .Y(n_1066) );
OAI31xp33_ASAP7_75t_L g1152 ( .A1(n_642), .A2(n_1153), .A3(n_1159), .B(n_1170), .Y(n_1152) );
OAI31xp33_ASAP7_75t_L g1477 ( .A1(n_642), .A2(n_1478), .A3(n_1485), .B(n_1491), .Y(n_1477) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g809 ( .A(n_645), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_751), .B1(n_752), .B2(n_808), .Y(n_645) );
INVx1_ASAP7_75t_L g808 ( .A(n_646), .Y(n_808) );
NAND3xp33_ASAP7_75t_SL g647 ( .A(n_648), .B(n_681), .C(n_696), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_665), .A3(n_675), .B(n_678), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g835 ( .A1(n_650), .A2(n_836), .B(n_837), .C(n_839), .Y(n_835) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g724 ( .A(n_651), .Y(n_724) );
INVx1_ASAP7_75t_L g831 ( .A(n_651), .Y(n_831) );
INVx2_ASAP7_75t_L g842 ( .A(n_651), .Y(n_842) );
INVx4_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx4f_ASAP7_75t_L g718 ( .A(n_652), .Y(n_718) );
BUFx4f_ASAP7_75t_L g763 ( .A(n_652), .Y(n_763) );
BUFx6f_ASAP7_75t_L g941 ( .A(n_652), .Y(n_941) );
BUFx4f_ASAP7_75t_L g1074 ( .A(n_652), .Y(n_1074) );
BUFx4f_ASAP7_75t_L g1330 ( .A(n_652), .Y(n_1330) );
OR2x6_ASAP7_75t_L g1752 ( .A(n_652), .B(n_1753), .Y(n_1752) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g874 ( .A(n_654), .Y(n_874) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_655), .B(n_1359), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_661), .B2(n_662), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_658), .A2(n_791), .B1(n_799), .B2(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_658), .A2(n_800), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_658), .A2(n_800), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_658), .A2(n_1043), .B1(n_1394), .B2(n_1407), .Y(n_1406) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_659), .A2(n_664), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_659), .A2(n_664), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_659), .A2(n_664), .B1(n_1445), .B2(n_1454), .Y(n_1453) );
OR2x2_ASAP7_75t_L g672 ( .A(n_660), .B(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_662), .A2(n_1041), .B1(n_1349), .B2(n_1361), .Y(n_1360) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g800 ( .A(n_664), .Y(n_800) );
INVx2_ASAP7_75t_L g1044 ( .A(n_664), .Y(n_1044) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_668), .Y(n_802) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_668), .Y(n_882) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_668), .Y(n_1047) );
INVx2_ASAP7_75t_L g1270 ( .A(n_670), .Y(n_1270) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g804 ( .A(n_672), .Y(n_804) );
INVx2_ASAP7_75t_L g884 ( .A(n_672), .Y(n_884) );
INVx8_ASAP7_75t_L g710 ( .A(n_673), .Y(n_710) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx4_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
CKINVDCx16_ASAP7_75t_R g806 ( .A(n_677), .Y(n_806) );
INVx3_ASAP7_75t_SL g880 ( .A(n_677), .Y(n_880) );
OAI31xp33_ASAP7_75t_L g1035 ( .A1(n_678), .A2(n_1036), .A3(n_1037), .B(n_1046), .Y(n_1035) );
OAI31xp33_ASAP7_75t_L g1205 ( .A1(n_678), .A2(n_1206), .A3(n_1207), .B(n_1211), .Y(n_1205) );
OAI31xp33_ASAP7_75t_L g1354 ( .A1(n_678), .A2(n_1355), .A3(n_1356), .B(n_1362), .Y(n_1354) );
BUFx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_SL g807 ( .A(n_679), .Y(n_807) );
OAI31xp33_ASAP7_75t_L g872 ( .A1(n_679), .A2(n_873), .A3(n_878), .B(n_881), .Y(n_872) );
INVx1_ASAP7_75t_L g1266 ( .A(n_679), .Y(n_1266) );
BUFx2_ASAP7_75t_L g1456 ( .A(n_679), .Y(n_1456) );
OAI31xp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_685), .A3(n_692), .B(n_695), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_686), .A2(n_855), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g865 ( .A(n_687), .Y(n_865) );
OAI31xp33_ASAP7_75t_L g921 ( .A1(n_695), .A2(n_922), .A3(n_926), .B(n_930), .Y(n_921) );
OAI31xp33_ASAP7_75t_L g1212 ( .A1(n_695), .A2(n_1213), .A3(n_1216), .B(n_1219), .Y(n_1212) );
OAI31xp33_ASAP7_75t_L g1256 ( .A1(n_695), .A2(n_1257), .A3(n_1258), .B(n_1261), .Y(n_1256) );
NOR2xp33_ASAP7_75t_SL g696 ( .A(n_697), .B(n_736), .Y(n_696) );
OAI33xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .A3(n_711), .B1(n_719), .B2(n_726), .B3(n_731), .Y(n_697) );
OAI33xp33_ASAP7_75t_L g908 ( .A1(n_698), .A2(n_726), .A3(n_909), .B1(n_916), .B2(n_919), .B3(n_920), .Y(n_908) );
INVx1_ASAP7_75t_L g1745 ( .A(n_698), .Y(n_1745) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx4_ASAP7_75t_L g756 ( .A(n_699), .Y(n_756) );
INVx2_ASAP7_75t_L g967 ( .A(n_699), .Y(n_967) );
INVx2_ASAP7_75t_L g1021 ( .A(n_699), .Y(n_1021) );
INVx1_ASAP7_75t_L g1383 ( .A(n_699), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_706), .B2(n_707), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_703), .A2(n_732), .B1(n_733), .B2(n_735), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_703), .A2(n_707), .B1(n_758), .B2(n_759), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_703), .A2(n_733), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g1242 ( .A(n_704), .Y(n_1242) );
INVx2_ASAP7_75t_L g1248 ( .A(n_704), .Y(n_1248) );
INVx3_ASAP7_75t_L g1428 ( .A(n_704), .Y(n_1428) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g912 ( .A(n_705), .Y(n_912) );
INVx4_ASAP7_75t_L g1497 ( .A(n_705), .Y(n_1497) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_706), .A2(n_725), .B1(n_748), .B2(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g1321 ( .A1(n_709), .A2(n_1322), .B1(n_1323), .B2(n_1325), .Y(n_1321) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g734 ( .A(n_710), .Y(n_734) );
INVx4_ASAP7_75t_L g915 ( .A(n_710), .Y(n_915) );
BUFx6f_ASAP7_75t_L g982 ( .A(n_710), .Y(n_982) );
INVx2_ASAP7_75t_L g1034 ( .A(n_710), .Y(n_1034) );
INVx2_ASAP7_75t_L g1072 ( .A(n_710), .Y(n_1072) );
INVx2_ASAP7_75t_L g1165 ( .A(n_710), .Y(n_1165) );
INVx1_ASAP7_75t_L g1243 ( .A(n_710), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_717), .B2(n_718), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_712), .A2(n_732), .B1(n_742), .B2(n_744), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_713), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx4_ASAP7_75t_L g973 ( .A(n_714), .Y(n_973) );
INVx2_ASAP7_75t_L g1246 ( .A(n_714), .Y(n_1246) );
INVx2_ASAP7_75t_L g1328 ( .A(n_714), .Y(n_1328) );
INVx4_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g722 ( .A(n_716), .Y(n_722) );
INVx2_ASAP7_75t_L g918 ( .A(n_716), .Y(n_918) );
BUFx2_ASAP7_75t_L g970 ( .A(n_716), .Y(n_970) );
INVx1_ASAP7_75t_L g1027 ( .A(n_716), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_718), .A2(n_896), .B1(n_900), .B2(n_917), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_718), .A2(n_891), .B1(n_907), .B2(n_917), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g1291 ( .A1(n_718), .A2(n_917), .B1(n_1292), .B2(n_1293), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_722), .A2(n_763), .B1(n_1373), .B2(n_1376), .Y(n_1384) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_724), .A2(n_973), .B1(n_974), .B2(n_975), .Y(n_972) );
OAI33xp33_ASAP7_75t_L g1285 ( .A1(n_726), .A2(n_967), .A3(n_1286), .B1(n_1291), .B2(n_1294), .B3(n_1297), .Y(n_1285) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI33xp33_ASAP7_75t_L g755 ( .A1(n_728), .A2(n_756), .A3(n_757), .B1(n_760), .B2(n_764), .B3(n_767), .Y(n_755) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_738), .A2(n_889), .B1(n_906), .B2(n_907), .Y(n_905) );
OAI22xp33_ASAP7_75t_L g999 ( .A1(n_738), .A2(n_1000), .B1(n_1001), .B2(n_1004), .Y(n_999) );
OAI22xp33_ASAP7_75t_L g1301 ( .A1(n_738), .A2(n_1287), .B1(n_1295), .B2(n_1302), .Y(n_1301) );
OAI22xp33_ASAP7_75t_L g1378 ( .A1(n_738), .A2(n_1015), .B1(n_1379), .B2(n_1380), .Y(n_1378) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_740), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_740), .A2(n_856), .B1(n_966), .B2(n_975), .Y(n_993) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_740), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_740), .Y(n_1239) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_742), .A2(n_1193), .B1(n_1376), .B2(n_1377), .Y(n_1375) );
INVx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx3_ASAP7_75t_L g746 ( .A(n_743), .Y(n_746) );
INVx2_ASAP7_75t_SL g861 ( .A(n_743), .Y(n_861) );
INVx2_ASAP7_75t_SL g990 ( .A(n_743), .Y(n_990) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_743), .B(n_1129), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_744), .A2(n_761), .B1(n_768), .B2(n_773), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_744), .A2(n_1233), .B1(n_1234), .B2(n_1235), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_744), .A2(n_776), .B1(n_1373), .B2(n_1374), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_746), .A2(n_898), .B1(n_900), .B2(n_901), .Y(n_899) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_749), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
INVx1_ASAP7_75t_L g1303 ( .A(n_749), .Y(n_1303) );
OAI22xp33_ASAP7_75t_L g1308 ( .A1(n_750), .A2(n_1290), .B1(n_1296), .B2(n_1309), .Y(n_1308) );
OAI22xp33_ASAP7_75t_L g1369 ( .A1(n_750), .A2(n_1015), .B1(n_1370), .B2(n_1371), .Y(n_1369) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_782), .C(n_795), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_770), .Y(n_754) );
INVx2_ASAP7_75t_SL g1416 ( .A(n_756), .Y(n_1416) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_762), .A2(n_769), .B1(n_776), .B2(n_779), .Y(n_775) );
INVx2_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx5_ASAP7_75t_L g778 ( .A(n_774), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_774), .A2(n_1111), .B1(n_1112), .B2(n_1113), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1139 ( .A(n_774), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1307 ( .A(n_774), .Y(n_1307) );
INVx3_ASAP7_75t_L g1778 ( .A(n_774), .Y(n_1778) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_776), .A2(n_896), .B1(n_897), .B2(n_898), .Y(n_895) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx8_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx3_ASAP7_75t_L g1011 ( .A(n_778), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_787), .A2(n_1015), .B1(n_1017), .B2(n_1018), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g1339 ( .A(n_788), .Y(n_1339) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g1436 ( .A(n_789), .Y(n_1436) );
OAI31xp33_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_801), .A3(n_805), .B(n_807), .Y(n_795) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_SL g1402 ( .A(n_804), .Y(n_1402) );
OAI31xp33_ASAP7_75t_L g939 ( .A1(n_807), .A2(n_940), .A3(n_945), .B(n_947), .Y(n_939) );
OAI31xp33_ASAP7_75t_L g1249 ( .A1(n_807), .A2(n_1250), .A3(n_1251), .B(n_1255), .Y(n_1249) );
OAI31xp33_ASAP7_75t_L g1398 ( .A1(n_807), .A2(n_1399), .A3(n_1400), .B(n_1403), .Y(n_1398) );
AO22x2_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_868), .B1(n_869), .B2(n_933), .Y(n_810) );
INVx1_ASAP7_75t_SL g933 ( .A(n_811), .Y(n_933) );
XNOR2x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NOR2x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_817), .Y(n_813) );
NAND3xp33_ASAP7_75t_SL g817 ( .A(n_818), .B(n_825), .C(n_850), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_821), .B1(n_822), .B2(n_823), .C(n_824), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_845), .B(n_849), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_835), .C(n_840), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_831), .B(n_832), .Y(n_830) );
OAI22xp5_ASAP7_75t_SL g968 ( .A1(n_831), .A2(n_969), .B1(n_970), .B2(n_971), .Y(n_968) );
OAI211xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B(n_843), .C(n_844), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_841), .A2(n_854), .B1(n_855), .B2(n_857), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_842), .A2(n_1004), .B1(n_1018), .B2(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx4_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx4f_ASAP7_75t_SL g855 ( .A(n_856), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g986 ( .A1(n_856), .A2(n_865), .B1(n_964), .B2(n_974), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_856), .A2(n_1053), .B1(n_1418), .B2(n_1424), .Y(n_1431) );
OAI22xp33_ASAP7_75t_L g1434 ( .A1(n_856), .A2(n_1419), .B1(n_1425), .B2(n_1435), .Y(n_1434) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g955 ( .A(n_858), .Y(n_955) );
INVx1_ASAP7_75t_L g1053 ( .A(n_858), .Y(n_1053) );
INVx1_ASAP7_75t_L g1279 ( .A(n_858), .Y(n_1279) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g1792 ( .A1(n_865), .A2(n_1748), .B(n_1793), .C(n_1795), .Y(n_1792) );
BUFx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g1122 ( .A(n_867), .B(n_1123), .C(n_1125), .Y(n_1122) );
AOI33xp33_ASAP7_75t_L g1465 ( .A1(n_867), .A2(n_1144), .A3(n_1466), .B1(n_1467), .B2(n_1468), .B3(n_1469), .Y(n_1465) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_885), .C(n_921), .Y(n_871) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g946 ( .A(n_884), .Y(n_946) );
INVx1_ASAP7_75t_L g1048 ( .A(n_884), .Y(n_1048) );
NOR2xp33_ASAP7_75t_SL g885 ( .A(n_886), .B(n_908), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_891), .B2(n_892), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_888), .A2(n_906), .B1(n_910), .B2(n_913), .Y(n_909) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g1309 ( .A(n_890), .Y(n_1309) );
INVx2_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_894), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_897), .A2(n_901), .B1(n_910), .B2(n_913), .Y(n_920) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_910), .A2(n_1183), .B1(n_1195), .B2(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_SL g911 ( .A(n_912), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_912), .A2(n_1189), .B1(n_1192), .B2(n_1199), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_913), .A2(n_1287), .B1(n_1288), .B2(n_1290), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_913), .A2(n_1288), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_915), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_915), .A2(n_1496), .B1(n_1497), .B2(n_1498), .Y(n_1495) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_918), .Y(n_1030) );
INVx2_ASAP7_75t_L g1484 ( .A(n_918), .Y(n_1484) );
INVx2_ASAP7_75t_SL g923 ( .A(n_924), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_1176), .B1(n_1312), .B2(n_1313), .Y(n_934) );
INVx1_ASAP7_75t_L g1312 ( .A(n_935), .Y(n_1312) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_1059), .B1(n_1060), .B2(n_1175), .Y(n_935) );
INVx1_ASAP7_75t_L g1175 ( .A(n_936), .Y(n_1175) );
XNOR2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_994), .Y(n_936) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_950), .C(n_961), .Y(n_938) );
OAI22xp5_ASAP7_75t_SL g1025 ( .A1(n_941), .A2(n_1006), .B1(n_1010), .B2(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1451 ( .A(n_948), .Y(n_1451) );
BUFx6f_ASAP7_75t_L g965 ( .A(n_949), .Y(n_965) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_949), .Y(n_1024) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_949), .Y(n_1070) );
OAI31xp33_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_953), .A3(n_958), .B(n_960), .Y(n_950) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g1786 ( .A1(n_955), .A2(n_1184), .B1(n_1744), .B2(n_1749), .C(n_1787), .Y(n_1786) );
OAI31xp33_ASAP7_75t_L g1438 ( .A1(n_960), .A2(n_1439), .A3(n_1443), .B(n_1447), .Y(n_1438) );
NOR2xp33_ASAP7_75t_SL g961 ( .A(n_962), .B(n_984), .Y(n_961) );
OAI33xp33_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_967), .A3(n_968), .B1(n_972), .B2(n_976), .B3(n_978), .Y(n_962) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_980), .B1(n_981), .B2(n_983), .Y(n_978) );
OAI22xp33_ASAP7_75t_L g1417 ( .A1(n_979), .A2(n_1071), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_981), .A2(n_1000), .B1(n_1017), .B2(n_1023), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_981), .A2(n_1023), .B1(n_1335), .B2(n_1336), .Y(n_1334) );
OAI22xp33_ASAP7_75t_L g1386 ( .A1(n_981), .A2(n_1374), .B1(n_1377), .B2(n_1387), .Y(n_1386) );
INVx5_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx6_ASAP7_75t_L g1199 ( .A(n_982), .Y(n_1199) );
OAI33xp33_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .A3(n_987), .B1(n_989), .B2(n_991), .B3(n_993), .Y(n_984) );
INVx1_ASAP7_75t_L g1144 ( .A(n_991), .Y(n_1144) );
OAI33xp33_ASAP7_75t_L g1430 ( .A1(n_991), .A2(n_998), .A3(n_1431), .B1(n_1432), .B2(n_1434), .B3(n_1437), .Y(n_1430) );
INVx3_ASAP7_75t_L g1787 ( .A(n_992), .Y(n_1787) );
NAND3xp33_ASAP7_75t_L g995 ( .A(n_996), .B(n_1035), .C(n_1049), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_1019), .Y(n_996) );
OAI33xp33_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .A3(n_1005), .B1(n_1009), .B2(n_1013), .B3(n_1014), .Y(n_997) );
OAI33xp33_ASAP7_75t_L g1224 ( .A1(n_998), .A2(n_1013), .A3(n_1225), .B1(n_1229), .B2(n_1232), .B3(n_1236), .Y(n_1224) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_1001), .A2(n_1322), .B1(n_1332), .B2(n_1339), .Y(n_1338) );
OAI22xp33_ASAP7_75t_L g1344 ( .A1(n_1001), .A2(n_1279), .B1(n_1325), .B2(n_1333), .Y(n_1344) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1003), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1007), .A2(n_1191), .B1(n_1192), .B2(n_1193), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_1008), .A2(n_1012), .B1(n_1023), .B2(n_1034), .Y(n_1033) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
OAI33xp33_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1022), .A3(n_1025), .B1(n_1028), .B2(n_1031), .B3(n_1033), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g1197 ( .A1(n_1020), .A2(n_1198), .A3(n_1200), .B1(n_1201), .B2(n_1203), .B3(n_1204), .Y(n_1197) );
OAI33xp33_ASAP7_75t_L g1240 ( .A1(n_1020), .A2(n_1203), .A3(n_1241), .B1(n_1244), .B2(n_1245), .B3(n_1247), .Y(n_1240) );
OAI33xp33_ASAP7_75t_L g1320 ( .A1(n_1020), .A2(n_1031), .A3(n_1321), .B1(n_1326), .B2(n_1331), .B3(n_1334), .Y(n_1320) );
BUFx6f_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g1747 ( .A1(n_1026), .A2(n_1074), .B1(n_1748), .B2(n_1749), .C(n_1750), .Y(n_1747) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_1029), .A2(n_1185), .B1(n_1196), .B2(n_1202), .Y(n_1201) );
INVx4_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
OAI33xp33_ASAP7_75t_L g1414 ( .A1(n_1031), .A2(n_1415), .A3(n_1417), .B1(n_1420), .B2(n_1423), .B3(n_1426), .Y(n_1414) );
OAI21xp5_ASAP7_75t_L g1746 ( .A1(n_1031), .A2(n_1747), .B(n_1752), .Y(n_1746) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1032), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_1034), .A2(n_1427), .B1(n_1428), .B2(n_1429), .Y(n_1426) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .B1(n_1043), .B2(n_1045), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1041), .A2(n_1043), .B1(n_1209), .B2(n_1210), .Y(n_1208) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
XOR2xp5_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1119), .Y(n_1061) );
XNOR2x1_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1105), .Y(n_1064) );
AOI21xp5_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1067), .B(n_1091), .Y(n_1065) );
NAND4xp25_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1076), .C(n_1080), .D(n_1086), .Y(n_1067) );
OAI21xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1073), .B(n_1075), .Y(n_1068) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1070), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1742 ( .A1(n_1070), .A2(n_1071), .B1(n_1743), .B2(n_1744), .Y(n_1742) );
BUFx6f_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
OAI211xp5_ASAP7_75t_SL g1076 ( .A1(n_1074), .A2(n_1077), .B(n_1078), .C(n_1079), .Y(n_1076) );
OAI211xp5_ASAP7_75t_SL g1080 ( .A1(n_1074), .A2(n_1081), .B(n_1082), .C(n_1084), .Y(n_1080) );
INVxp67_ASAP7_75t_L g1160 ( .A(n_1075), .Y(n_1160) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1789 ( .A(n_1094), .Y(n_1789) );
A2O1A1Ixp33_ASAP7_75t_L g1770 ( .A1(n_1098), .A2(n_1109), .B(n_1771), .C(n_1772), .Y(n_1770) );
XNOR2x1_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1174), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1145), .Y(n_1120) );
NAND4xp25_ASAP7_75t_SL g1121 ( .A(n_1122), .B(n_1126), .C(n_1130), .D(n_1136), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1128), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1128), .B(n_1472), .Y(n_1471) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_1129), .B(n_1133), .Y(n_1132) );
NAND3xp33_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1142), .C(n_1144), .Y(n_1136) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NAND3xp33_ASAP7_75t_SL g1145 ( .A(n_1146), .B(n_1149), .C(n_1152), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1151), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1151), .B(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
OAI21xp5_ASAP7_75t_SL g1159 ( .A1(n_1160), .A2(n_1161), .B(n_1166), .Y(n_1159) );
OAI21xp33_ASAP7_75t_L g1485 ( .A1(n_1160), .A2(n_1486), .B(n_1488), .Y(n_1485) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1176), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1264), .B1(n_1310), .B2(n_1311), .Y(n_1176) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1177), .Y(n_1310) );
XOR2x2_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1221), .Y(n_1177) );
AND3x1_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1205), .C(n_1212), .Y(n_1179) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1197), .Y(n_1180) );
OAI22xp33_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1184), .B1(n_1185), .B2(n_1186), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g1225 ( .A1(n_1184), .A2(n_1226), .B1(n_1227), .B2(n_1228), .Y(n_1225) );
OAI22xp33_ASAP7_75t_L g1236 ( .A1(n_1184), .A2(n_1237), .B1(n_1238), .B2(n_1239), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_1199), .A2(n_1231), .B1(n_1235), .B2(n_1248), .Y(n_1247) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_1199), .A2(n_1248), .B1(n_1370), .B2(n_1379), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_1202), .A2(n_1227), .B1(n_1238), .B2(n_1246), .Y(n_1245) );
OAI33xp33_ASAP7_75t_L g1381 ( .A1(n_1203), .A2(n_1382), .A3(n_1383), .B1(n_1384), .B2(n_1385), .B3(n_1386), .Y(n_1381) );
AND3x1_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1249), .C(n_1256), .Y(n_1222) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1240), .Y(n_1223) );
OAI22xp33_ASAP7_75t_L g1241 ( .A1(n_1226), .A2(n_1237), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1264), .Y(n_1311) );
OAI221xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1267), .B1(n_1276), .B2(n_1283), .C(n_1284), .Y(n_1265) );
NOR3xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1271), .C(n_1272), .Y(n_1267) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NOR3xp33_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .C(n_1282), .Y(n_1276) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1300), .Y(n_1284) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1314), .Y(n_1503) );
XOR2xp5_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1408), .Y(n_1314) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_1316), .A2(n_1317), .B1(n_1363), .B2(n_1364), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
NAND3xp33_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1345), .C(n_1354), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1337), .Y(n_1319) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1328), .B1(n_1329), .B2(n_1330), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1423 ( .A1(n_1328), .A2(n_1330), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1330), .Y(n_1405) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1343), .Y(n_1433) );
OAI31xp33_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1347), .A3(n_1351), .B(n_1353), .Y(n_1345) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
AND3x1_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1391), .C(n_1398), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1381), .Y(n_1367) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
AOI22xp5_ASAP7_75t_L g1409 ( .A1(n_1410), .A2(n_1411), .B1(n_1457), .B2(n_1502), .Y(n_1409) );
INVx2_ASAP7_75t_SL g1410 ( .A(n_1411), .Y(n_1410) );
NAND3xp33_ASAP7_75t_L g1412 ( .A(n_1413), .B(n_1438), .C(n_1448), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1430), .Y(n_1413) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
OAI31xp33_ASAP7_75t_SL g1448 ( .A1(n_1449), .A2(n_1452), .A3(n_1455), .B(n_1456), .Y(n_1448) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1458), .Y(n_1502) );
XNOR2x1_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1501), .Y(n_1458) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1473), .Y(n_1459) );
NAND3xp33_ASAP7_75t_L g1460 ( .A(n_1461), .B(n_1465), .C(n_1471), .Y(n_1460) );
NAND3xp33_ASAP7_75t_SL g1473 ( .A(n_1474), .B(n_1477), .C(n_1499), .Y(n_1473) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
OAI221xp5_ASAP7_75t_L g1504 ( .A1(n_1505), .A2(n_1719), .B1(n_1723), .B2(n_1796), .C(n_1800), .Y(n_1504) );
AOI211xp5_ASAP7_75t_L g1505 ( .A1(n_1506), .A2(n_1631), .B(n_1635), .C(n_1694), .Y(n_1505) );
NAND5xp2_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1566), .C(n_1582), .D(n_1601), .E(n_1623), .Y(n_1506) );
AOI211xp5_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1538), .B(n_1547), .C(n_1559), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1523), .Y(n_1508) );
INVx2_ASAP7_75t_L g1557 ( .A(n_1509), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1509), .B(n_1525), .Y(n_1576) );
AOI311xp33_ASAP7_75t_L g1601 ( .A1(n_1509), .A2(n_1602), .A3(n_1607), .B(n_1611), .C(n_1619), .Y(n_1601) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_1509), .B(n_1560), .Y(n_1627) );
OR2x2_ASAP7_75t_L g1653 ( .A(n_1509), .B(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1509), .B(n_1534), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_1509), .B(n_1530), .Y(n_1692) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1509), .B(n_1530), .Y(n_1709) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1518), .Y(n_1509) );
AND2x4_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1513), .Y(n_1511) );
AND2x6_ASAP7_75t_L g1516 ( .A(n_1512), .B(n_1517), .Y(n_1516) );
AND2x6_ASAP7_75t_L g1519 ( .A(n_1512), .B(n_1520), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1512), .B(n_1522), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1512), .B(n_1522), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1512), .B(n_1522), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1515), .Y(n_1513) );
OAI21xp5_ASAP7_75t_L g1809 ( .A1(n_1522), .A2(n_1810), .B(n_1811), .Y(n_1809) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1528), .Y(n_1523) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1524), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1524), .B(n_1609), .Y(n_1608) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1524), .B(n_1564), .Y(n_1620) );
OAI21xp33_ASAP7_75t_L g1641 ( .A1(n_1524), .A2(n_1642), .B(n_1643), .Y(n_1641) );
OAI332xp33_ASAP7_75t_L g1686 ( .A1(n_1524), .A2(n_1627), .A3(n_1687), .B1(n_1689), .B2(n_1690), .B3(n_1691), .C1(n_1692), .C2(n_1693), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1687 ( .A(n_1524), .B(n_1688), .Y(n_1687) );
CKINVDCx5p33_ASAP7_75t_R g1524 ( .A(n_1525), .Y(n_1524) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_1525), .B(n_1586), .Y(n_1585) );
INVx3_ASAP7_75t_L g1590 ( .A(n_1525), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1525), .B(n_1618), .Y(n_1624) );
NOR2xp33_ASAP7_75t_L g1650 ( .A(n_1525), .B(n_1593), .Y(n_1650) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1525), .B(n_1528), .Y(n_1654) );
OR2x2_ASAP7_75t_L g1708 ( .A(n_1525), .B(n_1709), .Y(n_1708) );
AND2x4_ASAP7_75t_SL g1525 ( .A(n_1526), .B(n_1527), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1528), .B(n_1576), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1534), .Y(n_1528) );
OR2x2_ASAP7_75t_L g1560 ( .A(n_1529), .B(n_1535), .Y(n_1560) );
AOI322xp5_ASAP7_75t_L g1623 ( .A1(n_1529), .A2(n_1609), .A3(n_1624), .B1(n_1625), .B2(n_1626), .C1(n_1628), .C2(n_1630), .Y(n_1623) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1530), .B(n_1535), .Y(n_1558) );
NOR2xp33_ASAP7_75t_L g1574 ( .A(n_1530), .B(n_1575), .Y(n_1574) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1530), .B(n_1594), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1530), .B(n_1557), .Y(n_1645) );
NOR3xp33_ASAP7_75t_SL g1679 ( .A(n_1530), .B(n_1555), .C(n_1631), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1532), .Y(n_1530) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1535), .Y(n_1588) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1535), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1535), .B(n_1557), .Y(n_1688) );
NAND2x1_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1537), .Y(n_1535) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1538), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1543), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1540), .Y(n_1562) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1540), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1540), .B(n_1543), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1540), .B(n_1544), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1542), .Y(n_1540) );
OR2x2_ASAP7_75t_L g1597 ( .A(n_1543), .B(n_1549), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1543), .B(n_1550), .Y(n_1610) );
HB1xp67_ASAP7_75t_SL g1659 ( .A(n_1543), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_1543), .B(n_1648), .Y(n_1691) );
CKINVDCx5p33_ASAP7_75t_R g1543 ( .A(n_1544), .Y(n_1543) );
NAND2xp5_ASAP7_75t_L g1564 ( .A(n_1544), .B(n_1565), .Y(n_1564) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1544), .B(n_1550), .Y(n_1569) );
HB1xp67_ASAP7_75t_SL g1595 ( .A(n_1544), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1544), .B(n_1562), .Y(n_1630) );
AND2x4_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1546), .Y(n_1544) );
NOR2xp33_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1553), .Y(n_1547) );
OAI32xp33_ASAP7_75t_L g1683 ( .A1(n_1548), .A2(n_1549), .A3(n_1613), .B1(n_1643), .B2(n_1684), .Y(n_1683) );
NAND2xp5_ASAP7_75t_L g1693 ( .A(n_1548), .B(n_1579), .Y(n_1693) );
INVx2_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1549), .B(n_1629), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1699 ( .A(n_1549), .B(n_1666), .Y(n_1699) );
INVx2_ASAP7_75t_SL g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1550), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1550), .B(n_1590), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1552), .Y(n_1550) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
O2A1O1Ixp33_ASAP7_75t_L g1649 ( .A1(n_1554), .A2(n_1650), .B(n_1651), .C(n_1652), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1556), .Y(n_1554) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_1555), .B(n_1581), .Y(n_1580) );
AOI221xp5_ASAP7_75t_L g1566 ( .A1(n_1556), .A2(n_1567), .B1(n_1570), .B2(n_1574), .C(n_1577), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
OR2x2_ASAP7_75t_L g1581 ( .A(n_1557), .B(n_1560), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1557), .B(n_1588), .Y(n_1587) );
OR2x2_ASAP7_75t_L g1592 ( .A(n_1557), .B(n_1593), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1557), .B(n_1590), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1638 ( .A(n_1557), .B(n_1639), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1557), .B(n_1606), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1702 ( .A(n_1557), .B(n_1599), .Y(n_1702) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1558), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1558), .B(n_1576), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1558), .B(n_1590), .Y(n_1639) );
NOR2xp33_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1561), .Y(n_1559) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1560), .Y(n_1605) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1561), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1563), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1567 ( .A(n_1562), .B(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1562), .Y(n_1618) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1562), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1562), .B(n_1617), .Y(n_1715) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1564), .Y(n_1642) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1564), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1565), .B(n_1584), .Y(n_1583) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1565), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1568), .B(n_1572), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1568), .B(n_1590), .Y(n_1682) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
NOR2xp33_ASAP7_75t_L g1717 ( .A(n_1569), .B(n_1590), .Y(n_1717) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
OAI332xp33_ASAP7_75t_L g1668 ( .A1(n_1573), .A2(n_1608), .A3(n_1654), .B1(n_1669), .B2(n_1670), .B3(n_1671), .C1(n_1672), .C2(n_1675), .Y(n_1668) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1576), .B(n_1606), .Y(n_1613) );
NOR2xp33_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1580), .Y(n_1577) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
AOI21xp33_ASAP7_75t_L g1619 ( .A1(n_1581), .A2(n_1620), .B(n_1621), .Y(n_1619) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1581), .Y(n_1664) );
AOI221xp5_ASAP7_75t_L g1582 ( .A1(n_1583), .A2(n_1585), .B1(n_1589), .B2(n_1595), .C(n_1596), .Y(n_1582) );
OAI31xp33_ASAP7_75t_L g1695 ( .A1(n_1584), .A2(n_1637), .A3(n_1696), .B(n_1698), .Y(n_1695) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
A2O1A1Ixp33_ASAP7_75t_L g1716 ( .A1(n_1588), .A2(n_1676), .B(n_1717), .C(n_1718), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1591), .Y(n_1589) );
NOR2xp33_ASAP7_75t_L g1646 ( .A(n_1590), .B(n_1597), .Y(n_1646) );
CKINVDCx14_ASAP7_75t_R g1663 ( .A(n_1590), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1697 ( .A(n_1591), .B(n_1617), .Y(n_1697) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1593), .Y(n_1606) );
A2O1A1Ixp33_ASAP7_75t_L g1636 ( .A1(n_1595), .A2(n_1637), .B(n_1640), .C(n_1648), .Y(n_1636) );
NOR2xp33_ASAP7_75t_L g1596 ( .A(n_1597), .B(n_1598), .Y(n_1596) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1597), .Y(n_1625) );
OAI22xp33_ASAP7_75t_L g1705 ( .A1(n_1597), .A2(n_1614), .B1(n_1621), .B2(n_1706), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1600), .Y(n_1598) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1600), .Y(n_1615) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1605), .B(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1609), .Y(n_1667) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
OR2x2_ASAP7_75t_L g1656 ( .A(n_1610), .B(n_1657), .Y(n_1656) );
AOI21xp5_ASAP7_75t_L g1611 ( .A1(n_1612), .A2(n_1614), .B(n_1616), .Y(n_1611) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
OAI22xp5_ASAP7_75t_L g1652 ( .A1(n_1616), .A2(n_1653), .B1(n_1655), .B2(n_1656), .Y(n_1652) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1616), .Y(n_1703) );
OR2x2_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1618), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1617), .B(n_1618), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1617), .B(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1617), .Y(n_1690) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1625), .B(n_1626), .Y(n_1647) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
NOR2xp33_ASAP7_75t_SL g1675 ( .A(n_1630), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1630), .Y(n_1710) );
INVx3_ASAP7_75t_L g1648 ( .A(n_1631), .Y(n_1648) );
NOR2xp33_ASAP7_75t_L g1676 ( .A(n_1631), .B(n_1657), .Y(n_1676) );
NOR3xp33_ASAP7_75t_L g1707 ( .A(n_1631), .B(n_1708), .C(n_1710), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1634), .Y(n_1631) );
HB1xp67_ASAP7_75t_L g1722 ( .A(n_1633), .Y(n_1722) );
NAND4xp25_ASAP7_75t_L g1635 ( .A(n_1636), .B(n_1649), .C(n_1658), .D(n_1677), .Y(n_1635) );
AOI22xp5_ASAP7_75t_L g1711 ( .A1(n_1637), .A2(n_1666), .B1(n_1712), .B2(n_1715), .Y(n_1711) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1639), .Y(n_1684) );
NAND3xp33_ASAP7_75t_SL g1640 ( .A(n_1641), .B(n_1644), .C(n_1647), .Y(n_1640) );
INVx2_ASAP7_75t_L g1655 ( .A(n_1643), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1643), .B(n_1663), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1645), .B(n_1646), .Y(n_1644) );
CKINVDCx14_ASAP7_75t_R g1669 ( .A(n_1645), .Y(n_1669) );
CKINVDCx14_ASAP7_75t_R g1670 ( .A(n_1648), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1648), .B(n_1657), .Y(n_1685) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1656), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1656), .B(n_1713), .Y(n_1712) );
AOI211xp5_ASAP7_75t_L g1658 ( .A1(n_1659), .A2(n_1660), .B(n_1661), .C(n_1668), .Y(n_1658) );
AOI21xp33_ASAP7_75t_L g1661 ( .A1(n_1662), .A2(n_1665), .B(n_1667), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1662 ( .A(n_1663), .B(n_1664), .Y(n_1662) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
CKINVDCx14_ASAP7_75t_R g1704 ( .A(n_1670), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1674), .Y(n_1672) );
OAI21xp5_ASAP7_75t_L g1680 ( .A1(n_1673), .A2(n_1681), .B(n_1683), .Y(n_1680) );
INVxp67_ASAP7_75t_SL g1689 ( .A(n_1676), .Y(n_1689) );
AOI221xp5_ASAP7_75t_L g1677 ( .A1(n_1678), .A2(n_1679), .B1(n_1680), .B2(n_1685), .C(n_1686), .Y(n_1677) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
NAND4xp25_ASAP7_75t_L g1694 ( .A(n_1695), .B(n_1700), .C(n_1711), .D(n_1716), .Y(n_1694) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
AOI311xp33_ASAP7_75t_L g1700 ( .A1(n_1701), .A2(n_1703), .A3(n_1704), .B(n_1705), .C(n_1707), .Y(n_1700) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1706), .Y(n_1718) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
CKINVDCx20_ASAP7_75t_R g1719 ( .A(n_1720), .Y(n_1719) );
CKINVDCx20_ASAP7_75t_R g1720 ( .A(n_1721), .Y(n_1720) );
INVx4_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
XNOR2x1_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1727), .Y(n_1725) );
HB1xp67_ASAP7_75t_L g1806 ( .A(n_1727), .Y(n_1806) );
NAND4xp75_ASAP7_75t_L g1727 ( .A(n_1728), .B(n_1737), .C(n_1761), .D(n_1764), .Y(n_1727) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
AOI211x1_ASAP7_75t_L g1737 ( .A1(n_1738), .A2(n_1745), .B(n_1746), .C(n_1756), .Y(n_1737) );
INVx2_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
NAND2x2_ASAP7_75t_L g1757 ( .A(n_1754), .B(n_1758), .Y(n_1757) );
INVx2_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
INVx2_ASAP7_75t_SL g1758 ( .A(n_1759), .Y(n_1758) );
AOI22xp33_ASAP7_75t_L g1775 ( .A1(n_1762), .A2(n_1763), .B1(n_1776), .B2(n_1777), .Y(n_1775) );
INVx4_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
INVx2_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
AOI21xp33_ASAP7_75t_L g1774 ( .A1(n_1775), .A2(n_1779), .B(n_1782), .Y(n_1774) );
INVx2_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
HB1xp67_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
OAI21xp5_ASAP7_75t_SL g1785 ( .A1(n_1786), .A2(n_1788), .B(n_1792), .Y(n_1785) );
INVx2_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
BUFx3_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
BUFx2_ASAP7_75t_SL g1801 ( .A(n_1802), .Y(n_1801) );
BUFx3_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
INVxp33_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
endmodule