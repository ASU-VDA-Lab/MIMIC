module fake_netlist_1_11324_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_9), .B(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
OAI22xp5_ASAP7_75t_SL g14 ( .A1(n_3), .A2(n_1), .B1(n_7), .B2(n_0), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
OR2x2_ASAP7_75t_L g17 ( .A(n_15), .B(n_2), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_16), .B(n_13), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_17), .A2(n_11), .B1(n_10), .B2(n_12), .Y(n_22) );
INVx5_ASAP7_75t_SL g23 ( .A(n_22), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
NAND2x1p5_ASAP7_75t_L g26 ( .A(n_24), .B(n_17), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_24), .B1(n_23), .B2(n_21), .Y(n_27) );
XOR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_14), .Y(n_28) );
OAI211xp5_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_19), .B(n_10), .C(n_11), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_23), .B1(n_20), .B2(n_18), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_23), .B1(n_18), .B2(n_19), .Y(n_31) );
INVxp67_ASAP7_75t_SL g32 ( .A(n_30), .Y(n_32) );
INVx2_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
OAI221xp5_ASAP7_75t_L g34 ( .A1(n_29), .A2(n_19), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_34) );
OR3x1_ASAP7_75t_L g35 ( .A(n_33), .B(n_2), .C(n_5), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI21xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_32), .B(n_34), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_36), .B1(n_35), .B2(n_8), .Y(n_38) );
endmodule