module fake_aes_2472_n_670 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_670);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_670;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_195;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g79 ( .A(n_27), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_57), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_8), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_73), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_31), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_24), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_21), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_45), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_53), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_14), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_77), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_26), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_76), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_17), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_8), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_18), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_7), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_64), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_22), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_62), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_56), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_19), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_54), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_5), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_32), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_36), .Y(n_112) );
XNOR2xp5_ASAP7_75t_L g113 ( .A(n_49), .B(n_66), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_20), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_75), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_14), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_65), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_68), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_39), .B(n_34), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_70), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_10), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_25), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_41), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_96), .B(n_108), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_95), .A2(n_33), .B(n_69), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_79), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_89), .B(n_0), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_82), .B(n_0), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_82), .B(n_1), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_111), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_111), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_79), .Y(n_146) );
BUFx8_ASAP7_75t_L g147 ( .A(n_79), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
NAND2xp33_ASAP7_75t_L g150 ( .A(n_84), .B(n_74), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_80), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_88), .B(n_1), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_88), .B(n_2), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_102), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_103), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_81), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_92), .B(n_3), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_90), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_83), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_83), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_125), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_104), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_92), .B(n_3), .Y(n_171) );
AO22x2_ASAP7_75t_L g172 ( .A1(n_143), .A2(n_126), .B1(n_98), .B2(n_114), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_134), .A2(n_110), .B1(n_101), .B2(n_123), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_128), .A2(n_126), .B1(n_114), .B2(n_98), .Y(n_174) );
INVx1_ASAP7_75t_SL g175 ( .A(n_162), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_134), .B(n_99), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_134), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_162), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_143), .A2(n_99), .B1(n_100), .B2(n_117), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_170), .B(n_119), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_170), .B(n_84), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
NOR3xp33_ASAP7_75t_L g186 ( .A(n_140), .B(n_100), .C(n_117), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_164), .B(n_93), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVxp33_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_160), .Y(n_193) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_139), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_140), .B(n_93), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_140), .B(n_94), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_163), .B(n_85), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_159), .B(n_94), .Y(n_200) );
AO22x2_ASAP7_75t_L g201 ( .A1(n_163), .A2(n_144), .B1(n_148), .B2(n_128), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_163), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_147), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_159), .B(n_124), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_136), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_165), .B(n_85), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_129), .B(n_116), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
NAND2xp33_ASAP7_75t_SL g213 ( .A(n_141), .B(n_122), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_165), .B(n_4), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_129), .B(n_116), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_147), .B(n_113), .C(n_112), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_136), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_130), .B(n_109), .Y(n_221) );
AND2x6_ASAP7_75t_L g222 ( .A(n_130), .B(n_121), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_167), .B(n_107), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_167), .B(n_118), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_169), .B(n_106), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_131), .B(n_113), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_169), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_139), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
BUFx10_ASAP7_75t_L g232 ( .A(n_131), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_147), .Y(n_233) );
INVx4_ASAP7_75t_SL g234 ( .A(n_132), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_139), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_132), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_194), .A2(n_171), .B1(n_141), .B2(n_156), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_201), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_232), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_201), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_193), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_232), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_227), .B(n_149), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_175), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_180), .Y(n_245) );
AND3x1_ASAP7_75t_L g246 ( .A(n_186), .B(n_171), .C(n_156), .Y(n_246) );
INVx5_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
INVx4_ASAP7_75t_SL g248 ( .A(n_198), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
NOR2x1p5_ASAP7_75t_L g250 ( .A(n_193), .B(n_157), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_172), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_221), .B(n_148), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_205), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_221), .B(n_149), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_221), .B(n_145), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_172), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_189), .B(n_153), .Y(n_260) );
INVxp33_ASAP7_75t_SL g261 ( .A(n_196), .Y(n_261) );
OR2x6_ASAP7_75t_L g262 ( .A(n_226), .B(n_157), .Y(n_262) );
NOR3xp33_ASAP7_75t_L g263 ( .A(n_179), .B(n_150), .C(n_137), .Y(n_263) );
BUFx2_ASAP7_75t_SL g264 ( .A(n_233), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_223), .B(n_137), .Y(n_265) );
CKINVDCx6p67_ASAP7_75t_R g266 ( .A(n_207), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_206), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_215), .B(n_144), .Y(n_268) );
OR2x2_ASAP7_75t_SL g269 ( .A(n_219), .B(n_138), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_223), .B(n_145), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_208), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_225), .B(n_152), .Y(n_274) );
AOI22xp5_ASAP7_75t_SL g275 ( .A1(n_226), .A2(n_192), .B1(n_197), .B2(n_233), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_225), .B(n_152), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_181), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_181), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_200), .B(n_153), .Y(n_279) );
BUFx8_ASAP7_75t_L g280 ( .A(n_176), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_181), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_177), .A2(n_178), .B1(n_188), .B2(n_194), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_224), .B(n_133), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_216), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_192), .A2(n_133), .B1(n_154), .B2(n_151), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_182), .B(n_133), .Y(n_287) );
OAI21xp33_ASAP7_75t_SL g288 ( .A1(n_183), .A2(n_151), .B(n_155), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_182), .B(n_154), .Y(n_291) );
AOI22xp5_ASAP7_75t_SL g292 ( .A1(n_184), .A2(n_138), .B1(n_161), .B2(n_155), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_202), .B(n_154), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_236), .B(n_154), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_210), .A2(n_151), .B1(n_161), .B2(n_155), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_213), .A2(n_154), .B1(n_161), .B2(n_168), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_210), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_183), .B(n_168), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_218), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_213), .A2(n_168), .B1(n_161), .B2(n_147), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_199), .B(n_168), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_211), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_209), .B(n_166), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_209), .A2(n_166), .B1(n_138), .B2(n_142), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_173), .B(n_166), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_302), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_289), .B(n_234), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_244), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_247), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_259), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_251), .A2(n_222), .B1(n_220), .B2(n_174), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_244), .B(n_174), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_267), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_245), .B(n_234), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_247), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_294), .A2(n_217), .B(n_214), .Y(n_317) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_239), .B(n_214), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_267), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_272), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_260), .B(n_222), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_280), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_272), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_242), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_238), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_240), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_268), .B(n_234), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_268), .A2(n_214), .B1(n_217), .B2(n_166), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_260), .B(n_222), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_247), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_247), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_242), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_242), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_266), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_249), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_264), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_258), .A2(n_222), .B1(n_217), .B2(n_166), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_279), .B(n_166), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_237), .A2(n_231), .B(n_135), .C(n_142), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_239), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_261), .B(n_222), .Y(n_345) );
NAND2xp33_ASAP7_75t_L g346 ( .A(n_284), .B(n_166), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_252), .B(n_166), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_273), .A2(n_138), .B1(n_135), .B2(n_142), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_284), .B(n_138), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_254), .B(n_231), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_265), .A2(n_185), .B(n_230), .C(n_229), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_289), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_261), .B(n_4), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_243), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_256), .B(n_5), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
INVx4_ASAP7_75t_L g358 ( .A(n_248), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_355), .A2(n_345), .B1(n_313), .B2(n_312), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_355), .B(n_262), .Y(n_362) );
OAI222xp33_ASAP7_75t_L g363 ( .A1(n_309), .A2(n_275), .B1(n_262), .B2(n_241), .C1(n_300), .C2(n_296), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_313), .B(n_262), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_339), .B(n_241), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_331), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_331), .A2(n_255), .B1(n_270), .B2(n_299), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_307), .Y(n_369) );
OAI22xp5_ASAP7_75t_SL g370 ( .A1(n_322), .A2(n_246), .B1(n_299), .B2(n_281), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_354), .A2(n_277), .B1(n_278), .B2(n_263), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_322), .A2(n_270), .B1(n_255), .B2(n_257), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_314), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_319), .Y(n_377) );
CKINVDCx6p67_ASAP7_75t_R g378 ( .A(n_337), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_319), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_320), .Y(n_380) );
OR2x6_ASAP7_75t_L g381 ( .A(n_332), .B(n_290), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_321), .A2(n_263), .B1(n_250), .B2(n_301), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_332), .B(n_248), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_323), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_332), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_320), .Y(n_386) );
CKINVDCx11_ASAP7_75t_R g387 ( .A(n_316), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_329), .A2(n_305), .B1(n_301), .B2(n_282), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_330), .B(n_274), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_383), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_365), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_382), .A2(n_271), .B1(n_276), .B2(n_282), .C(n_356), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_362), .A2(n_306), .B1(n_297), .B2(n_342), .Y(n_395) );
OAI222xp33_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_349), .B1(n_292), .B2(n_306), .C1(n_358), .C2(n_326), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_385), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_360), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_362), .A2(n_342), .B1(n_352), .B2(n_333), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_360), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_359), .A2(n_344), .B1(n_295), .B2(n_328), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_364), .B(n_325), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_288), .B1(n_295), .B2(n_291), .C(n_287), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_369), .B(n_325), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_370), .A2(n_352), .B1(n_333), .B2(n_330), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_361), .A2(n_326), .B1(n_338), .B2(n_253), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_363), .A2(n_366), .B1(n_375), .B2(n_390), .C(n_389), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_286), .B(n_304), .C(n_343), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_369), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_371), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_387), .A2(n_338), .B1(n_253), .B2(n_344), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_334), .B1(n_316), .B2(n_310), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_391), .B(n_327), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_304), .B(n_341), .C(n_283), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_334), .B1(n_336), .B2(n_340), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_367), .A2(n_346), .B1(n_293), .B2(n_347), .C(n_285), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_371), .B(n_340), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_376), .A2(n_315), .B1(n_293), .B2(n_327), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_394), .A2(n_317), .B(n_351), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_399), .B(n_376), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_399), .B(n_377), .Y(n_423) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_413), .B(n_381), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_408), .A2(n_381), .B1(n_379), .B2(n_384), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_401), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_401), .B(n_388), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_406), .B(n_388), .C(n_377), .D(n_384), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_418), .A2(n_379), .A3(n_385), .B(n_315), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_410), .B(n_374), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_410), .B(n_374), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_393), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_395), .A2(n_381), .B1(n_386), .B2(n_380), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_402), .A2(n_378), .B1(n_383), .B2(n_349), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_412), .A2(n_367), .B1(n_348), .B2(n_303), .C(n_386), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_414), .A2(n_380), .B1(n_383), .B2(n_308), .C(n_310), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_411), .B(n_349), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_397), .Y(n_438) );
AOI31xp33_ASAP7_75t_SL g439 ( .A1(n_403), .A2(n_6), .A3(n_7), .B(n_9), .Y(n_439) );
OAI21x1_ASAP7_75t_L g440 ( .A1(n_396), .A2(n_324), .B(n_335), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g441 ( .A1(n_409), .A2(n_383), .A3(n_308), .B(n_340), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_403), .B(n_308), .Y(n_442) );
OAI21x1_ASAP7_75t_L g443 ( .A1(n_393), .A2(n_324), .B(n_335), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_411), .B(n_308), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_407), .B(n_139), .C(n_146), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_400), .A2(n_349), .B1(n_269), .B2(n_336), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_419), .A2(n_349), .B1(n_358), .B2(n_357), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_405), .B(n_324), .Y(n_449) );
INVx6_ASAP7_75t_SL g450 ( .A(n_419), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_392), .A2(n_358), .B1(n_372), .B2(n_336), .Y(n_451) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_392), .B(n_358), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g454 ( .A1(n_420), .A2(n_318), .B(n_350), .C(n_146), .Y(n_454) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_417), .A2(n_191), .B(n_185), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_415), .A2(n_335), .B1(n_336), .B2(n_357), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_447), .B(n_417), .Y(n_457) );
AOI211xp5_ASAP7_75t_L g458 ( .A1(n_439), .A2(n_416), .B(n_419), .C(n_404), .Y(n_458) );
AOI33xp33_ASAP7_75t_L g459 ( .A1(n_425), .A2(n_398), .A3(n_230), .B1(n_229), .B2(n_203), .B3(n_191), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_424), .A2(n_392), .B1(n_398), .B2(n_372), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_428), .A2(n_357), .B1(n_372), .B2(n_397), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g462 ( .A(n_434), .B(n_372), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_437), .B(n_397), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_424), .A2(n_397), .B1(n_357), .B2(n_318), .Y(n_464) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_446), .A2(n_203), .B(n_190), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_447), .B(n_397), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_437), .B(n_9), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
OA332x1_ASAP7_75t_L g469 ( .A1(n_433), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_15), .C1(n_16), .C2(n_17), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_426), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_429), .A2(n_12), .A3(n_13), .B(n_15), .Y(n_472) );
INVx3_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_432), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_431), .B(n_16), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_454), .A2(n_357), .B(n_146), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_442), .B(n_19), .C(n_190), .D(n_187), .Y(n_477) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_421), .A2(n_187), .B(n_139), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_248), .B1(n_146), .B2(n_139), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_435), .A2(n_146), .B1(n_228), .B2(n_212), .C(n_195), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_449), .B(n_146), .C(n_28), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_438), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_432), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_455), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_453), .B(n_146), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_422), .B(n_23), .Y(n_488) );
OAI31xp33_ASAP7_75t_L g489 ( .A1(n_441), .A2(n_30), .A3(n_35), .B(n_37), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_455), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_453), .B(n_38), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_427), .B(n_40), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_450), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_443), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_453), .B(n_444), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_443), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_445), .B(n_235), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_448), .B(n_42), .Y(n_498) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_456), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_440), .B(n_44), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_455), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_456), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_455), .B(n_47), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_450), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_493), .Y(n_506) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_477), .A2(n_452), .A3(n_450), .B(n_451), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_463), .B(n_471), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_468), .B(n_452), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_463), .B(n_484), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_483), .B(n_50), .Y(n_511) );
NAND2xp67_ASAP7_75t_L g512 ( .A(n_475), .B(n_51), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_486), .B(n_52), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_486), .B(n_55), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_470), .B(n_58), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_485), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_474), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_485), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_474), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_474), .B(n_59), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_483), .B(n_60), .Y(n_523) );
OAI31xp33_ASAP7_75t_L g524 ( .A1(n_477), .A2(n_61), .A3(n_63), .B(n_67), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_484), .B(n_195), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_484), .Y(n_526) );
OAI21xp33_ASAP7_75t_L g527 ( .A1(n_460), .A2(n_195), .B(n_212), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_472), .B(n_212), .C(n_228), .D(n_235), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_473), .B(n_228), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_473), .B(n_228), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_473), .B(n_235), .Y(n_531) );
BUFx2_ASAP7_75t_L g532 ( .A(n_482), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_482), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_466), .B(n_235), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_467), .B(n_505), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_466), .B(n_490), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_475), .B(n_467), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_457), .B(n_502), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_500), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_490), .B(n_460), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_494), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_494), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_472), .A2(n_495), .B1(n_498), .B2(n_489), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_500), .B(n_487), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_496), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_459), .B(n_458), .C(n_488), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_487), .B(n_496), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_461), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_493), .A2(n_498), .B1(n_469), .B2(n_505), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_465), .B(n_501), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_461), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_478), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_465), .B(n_501), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_465), .B(n_503), .Y(n_556) );
OAI211xp5_ASAP7_75t_L g557 ( .A1(n_458), .A2(n_489), .B(n_462), .C(n_505), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_499), .B(n_465), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_504), .B(n_478), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_488), .B(n_492), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_508), .B(n_464), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_548), .A2(n_491), .B1(n_481), .B2(n_492), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_538), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_538), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_507), .B(n_491), .C(n_476), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_532), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_508), .B(n_504), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_510), .B(n_478), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_532), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_510), .B(n_497), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_513), .B(n_497), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_539), .B(n_476), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g573 ( .A(n_507), .B(n_479), .C(n_480), .D(n_551), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_557), .B(n_560), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_539), .B(n_537), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_533), .B(n_536), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_506), .B(n_535), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g578 ( .A1(n_528), .A2(n_524), .B(n_523), .C(n_516), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_533), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_544), .A2(n_509), .B1(n_523), .B2(n_527), .C(n_555), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_517), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_510), .B(n_509), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_517), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_513), .B(n_527), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_510), .B(n_549), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_516), .A2(n_552), .B(n_555), .C(n_511), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_546), .A2(n_554), .B(n_519), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_526), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_518), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_520), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_521), .B(n_526), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_549), .B(n_545), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_513), .B(n_514), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_540), .Y(n_594) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_552), .A2(n_541), .B(n_556), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_512), .B(n_558), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_514), .B(n_515), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_542), .Y(n_598) );
OA21x2_ASAP7_75t_L g599 ( .A1(n_558), .A2(n_554), .B(n_547), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_563), .B(n_558), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_574), .A2(n_558), .B1(n_543), .B2(n_547), .C(n_559), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_564), .B(n_543), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_574), .B(n_512), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_575), .B(n_553), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_571), .B(n_546), .Y(n_605) );
NOR2x1_ASAP7_75t_L g606 ( .A(n_565), .B(n_515), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_594), .B(n_550), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_585), .B(n_546), .Y(n_608) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_578), .A2(n_522), .B(n_546), .Y(n_609) );
XNOR2xp5_ASAP7_75t_L g610 ( .A(n_582), .B(n_529), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_579), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_576), .B(n_534), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_568), .B(n_529), .Y(n_613) );
AO22x2_ASAP7_75t_L g614 ( .A1(n_566), .A2(n_534), .B1(n_530), .B2(n_531), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_598), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_595), .B(n_530), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_598), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_599), .B(n_531), .Y(n_618) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_590), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_599), .B(n_525), .Y(n_620) );
NAND3x1_ASAP7_75t_L g621 ( .A(n_593), .B(n_525), .C(n_597), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_580), .A2(n_573), .B(n_596), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_591), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_577), .B(n_566), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_569), .B(n_579), .Y(n_625) );
NOR2xp33_ASAP7_75t_SL g626 ( .A(n_578), .B(n_580), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_589), .B(n_569), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_561), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_583), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_562), .A2(n_596), .B1(n_586), .B2(n_570), .Y(n_630) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_584), .B(n_567), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_588), .Y(n_632) );
NAND2x1_ASAP7_75t_L g633 ( .A(n_571), .B(n_581), .Y(n_633) );
AOI322xp5_ASAP7_75t_L g634 ( .A1(n_583), .A2(n_574), .A3(n_592), .B1(n_597), .B2(n_577), .C1(n_544), .C2(n_551), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_587), .A2(n_584), .B(n_578), .Y(n_635) );
XOR2xp5_ASAP7_75t_L g636 ( .A(n_572), .B(n_587), .Y(n_636) );
NOR2x1_ASAP7_75t_L g637 ( .A(n_565), .B(n_528), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_574), .A2(n_595), .B(n_580), .Y(n_638) );
INVxp67_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
OAI322xp33_ASAP7_75t_L g640 ( .A1(n_626), .A2(n_636), .A3(n_635), .B1(n_628), .B2(n_630), .C1(n_639), .C2(n_609), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_627), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g642 ( .A1(n_622), .A2(n_638), .B(n_603), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_603), .A2(n_637), .B1(n_606), .B2(n_631), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_616), .A2(n_601), .B1(n_624), .B2(n_635), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_616), .A2(n_604), .B1(n_614), .B2(n_621), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_608), .A2(n_614), .B1(n_605), .B2(n_613), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_614), .A2(n_623), .B1(n_617), .B2(n_615), .C(n_629), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_627), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_611), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_605), .B(n_629), .C(n_625), .Y(n_650) );
XOR2xp5_ASAP7_75t_L g651 ( .A(n_610), .B(n_612), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g652 ( .A(n_642), .B(n_634), .C(n_633), .Y(n_652) );
NOR4xp25_ASAP7_75t_L g653 ( .A(n_640), .B(n_621), .C(n_632), .D(n_619), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_641), .B(n_602), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_648), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_643), .A2(n_618), .B(n_620), .C(n_600), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_649), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_650), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_652), .B(n_645), .C(n_644), .D(n_646), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_655), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_652), .A2(n_647), .B1(n_651), .B2(n_607), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_660), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_659), .B(n_658), .C(n_656), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_661), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_663), .B(n_657), .Y(n_665) );
XOR2xp5_ASAP7_75t_L g666 ( .A(n_664), .B(n_654), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_665), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_667), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_668), .Y(n_669) );
O2A1O1Ixp5_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_662), .B(n_666), .C(n_653), .Y(n_670) );
endmodule