module fake_netlist_6_1897_n_1734 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1734);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1734;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_73),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_20),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_114),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_25),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_90),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_46),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_84),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_38),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_67),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_12),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_31),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_76),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_120),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_66),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_68),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_57),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_39),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_5),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_58),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_126),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_59),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_51),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_20),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_29),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_55),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_49),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_119),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_117),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_121),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_52),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_24),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_142),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_93),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_50),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_24),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_69),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_38),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_133),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_18),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_138),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_111),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_100),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_8),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_131),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_116),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_125),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_78),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_56),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_21),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_16),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_139),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_130),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_115),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_153),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_18),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_87),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_23),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_135),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_64),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_31),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_46),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_30),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_122),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_102),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_82),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_6),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_39),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_83),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_33),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_28),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_108),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_19),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_85),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_63),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_89),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_71),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_140),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_48),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_77),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_27),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_25),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_149),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_3),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_3),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_21),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_65),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_146),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_99),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_33),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_49),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_61),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_62),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_60),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_11),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_5),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_129),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_14),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_92),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_42),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_53),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_159),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_41),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_26),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_54),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_136),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_48),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_35),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_35),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_15),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_37),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_27),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_55),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_26),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_79),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_163),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_184),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_184),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_0),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_198),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_165),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_202),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_205),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_167),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_175),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_205),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_168),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_316),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_169),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_172),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_264),
.B(n_0),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_192),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_199),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_194),
.B(n_2),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_174),
.B(n_4),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_219),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_234),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_234),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_196),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_197),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_203),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_204),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_331),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_207),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_291),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_268),
.B(n_7),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_212),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_245),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_214),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_225),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_214),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_231),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_235),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_291),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_291),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_174),
.B(n_7),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_247),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_191),
.B(n_213),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_191),
.B(n_213),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_247),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_285),
.B(n_9),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_199),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_187),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_264),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_235),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_239),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_210),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_217),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_241),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_219),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_220),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_263),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_248),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_251),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_263),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_199),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_200),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_240),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_285),
.B(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_242),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_257),
.Y(n_416)
);

BUFx6f_ASAP7_75t_SL g417 ( 
.A(n_171),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_162),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_254),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_335),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_195),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_345),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_245),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_334),
.B(n_170),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_359),
.B(n_268),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_334),
.B(n_173),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_350),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_380),
.B(n_215),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_337),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_367),
.B(n_229),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_338),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_R g451 ( 
.A(n_355),
.B(n_258),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_366),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_339),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_340),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_392),
.B(n_180),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_344),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_374),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_346),
.B(n_185),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_351),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_343),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_351),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_392),
.B(n_193),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_398),
.B(n_201),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_377),
.B(n_176),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_357),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_358),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_347),
.A2(n_166),
.B1(n_261),
.B2(n_302),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_391),
.B(n_211),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_360),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_397),
.Y(n_482)
);

CKINVDCx11_ASAP7_75t_R g483 ( 
.A(n_348),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_361),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_342),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_369),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_401),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_394),
.B(n_414),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_378),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_365),
.A2(n_266),
.B(n_255),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_370),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_482),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_494),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_482),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_437),
.B(n_372),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_219),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_420),
.B(n_166),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_435),
.B(n_378),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_373),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_435),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_219),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_437),
.B(n_376),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_492),
.B(n_379),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_382),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_426),
.Y(n_517)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

AND3x2_ASAP7_75t_L g519 ( 
.A(n_442),
.B(n_363),
.C(n_467),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_288),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_424),
.B(n_384),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_480),
.A2(n_388),
.B1(n_356),
.B2(n_375),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_461),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_398),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_439),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_451),
.B(n_400),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_435),
.B(n_441),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_435),
.B(n_403),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_497),
.B(n_408),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_496),
.B(n_288),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_443),
.B(n_409),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_448),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_436),
.B(n_416),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_423),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_423),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_440),
.B(n_418),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_453),
.B(n_362),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_448),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_448),
.B(n_216),
.Y(n_549)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_496),
.B(n_259),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_475),
.A2(n_417),
.B1(n_396),
.B2(n_411),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_442),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_458),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_475),
.B(n_419),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_472),
.B(n_171),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_458),
.B(n_228),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_486),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_483),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_440),
.B(n_186),
.C(n_164),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_473),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_458),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_430),
.A2(n_261),
.B1(n_302),
.B2(n_321),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_444),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_462),
.B(n_230),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_480),
.A2(n_319),
.B1(n_278),
.B2(n_282),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_429),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_462),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_480),
.A2(n_292),
.B1(n_267),
.B2(n_284),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_481),
.B(n_171),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_463),
.B(n_236),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_433),
.B(n_419),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_243),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_486),
.B(n_288),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_484),
.B(n_487),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_461),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_433),
.B(n_405),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_463),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_486),
.B(n_288),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_486),
.B(n_296),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_470),
.B(n_417),
.Y(n_585)
);

INVxp33_ASAP7_75t_L g586 ( 
.A(n_476),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_470),
.B(n_190),
.C(n_189),
.Y(n_587)
);

CKINVDCx6p67_ASAP7_75t_R g588 ( 
.A(n_483),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_465),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_480),
.B(n_206),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_465),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_480),
.B(n_222),
.C(n_218),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_427),
.B(n_405),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_496),
.Y(n_594)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_427),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_433),
.B(n_349),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_496),
.A2(n_181),
.B1(n_176),
.B2(n_183),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_469),
.B(n_206),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_469),
.B(n_413),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_453),
.B(n_298),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_469),
.B(n_354),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_465),
.B(n_244),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_457),
.B(n_206),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_488),
.Y(n_604)
);

INVxp33_ASAP7_75t_SL g605 ( 
.A(n_476),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_488),
.A2(n_321),
.B1(n_277),
.B2(n_330),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_444),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_496),
.B(n_246),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_468),
.B(n_296),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_468),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_460),
.B(n_249),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_468),
.B(n_221),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_461),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_489),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_489),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_460),
.A2(n_490),
.B1(n_491),
.B2(n_332),
.Y(n_616)
);

OAI22x1_ASAP7_75t_L g617 ( 
.A1(n_490),
.A2(n_312),
.B1(n_223),
.B2(n_301),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_491),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_421),
.B(n_413),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_421),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_428),
.Y(n_621)
);

NAND3x1_ASAP7_75t_L g622 ( 
.A(n_485),
.B(n_300),
.C(n_327),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_444),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_422),
.B(n_250),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_446),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_422),
.B(n_252),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_425),
.B(n_296),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_444),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_422),
.B(n_253),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_425),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_432),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_428),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_485),
.B(n_415),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_445),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_445),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_447),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_447),
.B(n_381),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_449),
.B(n_383),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_449),
.B(n_311),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_614),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_508),
.A2(n_269),
.B1(n_280),
.B2(n_324),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_558),
.B(n_415),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_515),
.B(n_177),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_524),
.B(n_493),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_594),
.A2(n_260),
.B1(n_317),
.B2(n_274),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_615),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_518),
.A2(n_385),
.B1(n_399),
.B2(n_406),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_618),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_596),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_620),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_594),
.A2(n_273),
.B1(n_493),
.B2(n_320),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_557),
.B(n_311),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_506),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_630),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_631),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_558),
.B(n_224),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_518),
.Y(n_657)
);

AOI221xp5_ASAP7_75t_L g658 ( 
.A1(n_606),
.A2(n_313),
.B1(n_322),
.B2(n_325),
.C(n_238),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_557),
.B(n_311),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_546),
.B(n_177),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_518),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_570),
.B(n_493),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_554),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_499),
.B(n_178),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_517),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_545),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_610),
.B(n_540),
.Y(n_667)
);

NOR2x1p5_ASAP7_75t_L g668 ( 
.A(n_588),
.B(n_226),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_565),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_601),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_540),
.B(n_450),
.Y(n_671)
);

BUFx4_ASAP7_75t_L g672 ( 
.A(n_625),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_507),
.B(n_454),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_498),
.B(n_459),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_502),
.B(n_459),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_593),
.B(n_471),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_539),
.B(n_320),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_509),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_499),
.B(n_178),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_593),
.B(n_471),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_608),
.A2(n_320),
.B1(n_478),
.B2(n_477),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_530),
.B(n_474),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_634),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_530),
.B(n_477),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_578),
.B(n_265),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_539),
.B(n_479),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_636),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_536),
.B(n_479),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_635),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_536),
.B(n_495),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_516),
.B(n_495),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_503),
.B(n_179),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_595),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_595),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_525),
.B(n_179),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_595),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_575),
.B(n_410),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_534),
.B(n_276),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_552),
.B(n_227),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_619),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_500),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_SL g702 ( 
.A(n_511),
.B(n_444),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_510),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_500),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_513),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_619),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_580),
.B(n_208),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_599),
.A2(n_299),
.B1(n_293),
.B2(n_221),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_514),
.B(n_181),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_560),
.B(n_182),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_547),
.B(n_600),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_599),
.B(n_495),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_600),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_534),
.B(n_283),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_600),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_585),
.B(n_431),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_592),
.B(n_182),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_526),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_550),
.B(n_286),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_500),
.B(n_431),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_550),
.B(n_289),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_590),
.B(n_183),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_633),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_597),
.B(n_294),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_562),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_527),
.B(n_431),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_587),
.B(n_333),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_569),
.A2(n_333),
.B1(n_309),
.B2(n_304),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_529),
.B(n_531),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_637),
.B(n_233),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_638),
.B(n_237),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_598),
.A2(n_305),
.B1(n_306),
.B2(n_310),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_549),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_532),
.B(n_535),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_537),
.B(n_434),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_505),
.B(n_208),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_549),
.A2(n_395),
.B(n_393),
.C(n_434),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_541),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_528),
.B(n_314),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_548),
.B(n_553),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_538),
.B(n_256),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_563),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_547),
.B(n_208),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_566),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_556),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_542),
.B(n_262),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_571),
.B(n_434),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_547),
.B(n_209),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_582),
.Y(n_749)
);

INVxp33_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_556),
.A2(n_395),
.B(n_456),
.C(n_455),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_589),
.B(n_444),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_511),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_591),
.B(n_444),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_569),
.A2(n_295),
.B(n_271),
.C(n_329),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_561),
.B(n_221),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_613),
.B(n_452),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_579),
.B(n_293),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_616),
.B(n_452),
.Y(n_759)
);

AO221x1_ASAP7_75t_L g760 ( 
.A1(n_606),
.A2(n_293),
.B1(n_299),
.B2(n_209),
.C(n_232),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_555),
.B(n_573),
.Y(n_761)
);

BUFx8_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_605),
.A2(n_299),
.B1(n_464),
.B2(n_209),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_568),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_604),
.A2(n_464),
.B1(n_232),
.B2(n_323),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_603),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_581),
.B(n_452),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_501),
.B(n_452),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_533),
.B(n_287),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_501),
.B(n_452),
.Y(n_770)
);

NOR3x1_ASAP7_75t_L g771 ( 
.A(n_612),
.B(n_232),
.C(n_270),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_519),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_632),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_568),
.A2(n_272),
.B(n_275),
.C(n_279),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_521),
.B(n_452),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_504),
.B(n_281),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_572),
.A2(n_326),
.B1(n_318),
.B2(n_308),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_521),
.B(n_428),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_574),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_519),
.B(n_290),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_522),
.B(n_428),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_564),
.B(n_297),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_504),
.B(n_307),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_522),
.B(n_428),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_504),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_543),
.B(n_161),
.Y(n_786)
);

NAND2x1_ASAP7_75t_L g787 ( 
.A(n_621),
.B(n_156),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_564),
.B(n_10),
.C(n_11),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_543),
.B(n_154),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_572),
.A2(n_602),
.B(n_576),
.C(n_611),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_551),
.B(n_13),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_586),
.B(n_13),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_576),
.B(n_132),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_504),
.Y(n_794)
);

OAI321xp33_ASAP7_75t_L g795 ( 
.A1(n_658),
.A2(n_611),
.A3(n_602),
.B1(n_629),
.B2(n_624),
.C(n_626),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_657),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_641),
.A2(n_583),
.B(n_626),
.C(n_629),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_646),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_686),
.A2(n_624),
.B(n_577),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_712),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_730),
.A2(n_609),
.B(n_628),
.C(n_567),
.Y(n_801)
);

AOI21x1_ASAP7_75t_L g802 ( 
.A1(n_677),
.A2(n_767),
.B(n_757),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_790),
.A2(n_577),
.B(n_584),
.Y(n_803)
);

AO21x1_ASAP7_75t_L g804 ( 
.A1(n_721),
.A2(n_512),
.B(n_523),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_670),
.B(n_559),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_665),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_691),
.B(n_584),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_649),
.B(n_544),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_648),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_792),
.A2(n_622),
.B1(n_628),
.B2(n_544),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_730),
.A2(n_577),
.B1(n_512),
.B2(n_523),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_677),
.A2(n_577),
.B(n_512),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_767),
.A2(n_584),
.B(n_523),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_697),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_733),
.B(n_584),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_707),
.B(n_663),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_699),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_745),
.B(n_512),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_704),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_764),
.A2(n_523),
.B(n_577),
.Y(n_820)
);

BUFx12f_ASAP7_75t_L g821 ( 
.A(n_762),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_644),
.A2(n_623),
.B(n_520),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_660),
.B(n_22),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_731),
.B(n_660),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_650),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_650),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_779),
.A2(n_639),
.B(n_627),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_654),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_654),
.Y(n_829)
);

CKINVDCx10_ASAP7_75t_R g830 ( 
.A(n_672),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_688),
.A2(n_639),
.B(n_627),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_721),
.A2(n_639),
.B(n_627),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_792),
.A2(n_607),
.B1(n_29),
.B2(n_30),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_655),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_655),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_731),
.A2(n_22),
.B(n_32),
.C(n_34),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_662),
.A2(n_639),
.B(n_627),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_671),
.B(n_36),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_SL g839 ( 
.A(n_761),
.B(n_725),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_690),
.B(n_683),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_36),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_768),
.A2(n_775),
.B(n_770),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_643),
.B(n_128),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_687),
.B(n_673),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_704),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_643),
.A2(n_40),
.B(n_43),
.C(n_44),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_666),
.A2(n_105),
.B1(n_103),
.B2(n_96),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_719),
.A2(n_81),
.B(n_80),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_SL g849 ( 
.A(n_703),
.B(n_705),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_682),
.A2(n_40),
.B(n_43),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_687),
.B(n_44),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_684),
.A2(n_45),
.B(n_47),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_723),
.B(n_47),
.Y(n_853)
);

BUFx4f_ASAP7_75t_L g854 ( 
.A(n_711),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_703),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_664),
.B(n_50),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_720),
.A2(n_52),
.B(n_53),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_653),
.B(n_54),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_651),
.A2(n_645),
.B(n_681),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_693),
.A2(n_696),
.B(n_694),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_759),
.A2(n_676),
.B(n_680),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_717),
.A2(n_692),
.B(n_709),
.C(n_722),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_718),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_674),
.B(n_675),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_685),
.B(n_741),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_778),
.A2(n_784),
.B(n_781),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_716),
.A2(n_753),
.B(n_661),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_664),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_669),
.B(n_692),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_709),
.B(n_678),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_718),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_679),
.B(n_717),
.C(n_710),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_753),
.A2(n_729),
.B(n_734),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_700),
.B(n_706),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_753),
.A2(n_740),
.B(n_714),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_679),
.B(n_769),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_724),
.A2(n_698),
.B(n_714),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_701),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_698),
.A2(n_755),
.B(n_744),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_769),
.B(n_722),
.Y(n_880)
);

BUFx4f_ASAP7_75t_L g881 ( 
.A(n_711),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_738),
.A2(n_749),
.B(n_744),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_742),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_741),
.B(n_746),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_727),
.A2(n_710),
.B(n_746),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_753),
.A2(n_652),
.B(n_659),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_652),
.A2(n_659),
.B(n_754),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_766),
.B(n_736),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_701),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_752),
.A2(n_739),
.B(n_786),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_727),
.A2(n_739),
.B1(n_689),
.B2(n_640),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_695),
.A2(n_774),
.B(n_793),
.C(n_751),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_789),
.A2(n_773),
.B(n_735),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_773),
.A2(n_747),
.B(n_726),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_713),
.B(n_715),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_642),
.B(n_647),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_772),
.A2(n_780),
.B1(n_750),
.B2(n_758),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_656),
.B(n_782),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_793),
.A2(n_787),
.B(n_783),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_728),
.B(n_758),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_756),
.B(n_708),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_785),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_785),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_756),
.B(n_732),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_794),
.B(n_702),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_780),
.B(n_748),
.Y(n_906)
);

CKINVDCx10_ASAP7_75t_R g907 ( 
.A(n_711),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_791),
.Y(n_908)
);

BUFx4f_ASAP7_75t_L g909 ( 
.A(n_743),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_771),
.Y(n_910)
);

BUFx8_ASAP7_75t_L g911 ( 
.A(n_762),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_763),
.A2(n_777),
.B1(n_788),
.B2(n_765),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_776),
.B(n_737),
.C(n_760),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_668),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_762),
.A2(n_492),
.B(n_641),
.C(n_667),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_667),
.B(n_508),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_686),
.A2(n_790),
.B(n_594),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_667),
.B(n_508),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_646),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_712),
.Y(n_920)
);

CKINVDCx8_ASAP7_75t_R g921 ( 
.A(n_665),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_667),
.B(n_508),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_670),
.B(n_508),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_SL g924 ( 
.A(n_730),
.B(n_505),
.C(n_731),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_704),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_670),
.B(n_649),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_646),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_667),
.A2(n_492),
.B1(n_572),
.B2(n_569),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_667),
.B(n_508),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_712),
.Y(n_930)
);

BUFx4f_ASAP7_75t_L g931 ( 
.A(n_711),
.Y(n_931)
);

AOI21x1_ASAP7_75t_L g932 ( 
.A1(n_677),
.A2(n_686),
.B(n_767),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_641),
.A2(n_492),
.B(n_667),
.C(n_724),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_721),
.A2(n_677),
.B(n_659),
.C(n_652),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_704),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_700),
.B(n_706),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_641),
.A2(n_492),
.B(n_667),
.C(n_724),
.Y(n_937)
);

AO21x1_ASAP7_75t_L g938 ( 
.A1(n_721),
.A2(n_677),
.B(n_719),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_733),
.B(n_745),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_712),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_670),
.B(n_649),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_733),
.B(n_745),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_700),
.B(n_706),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_733),
.A2(n_508),
.B1(n_764),
.B2(n_745),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_657),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_667),
.A2(n_492),
.B1(n_572),
.B2(n_569),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_733),
.B(n_745),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_712),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_670),
.B(n_649),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_733),
.B(n_745),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_824),
.B(n_884),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_921),
.Y(n_952)
);

OAI22xp33_ASAP7_75t_L g953 ( 
.A1(n_876),
.A2(n_880),
.B1(n_922),
.B2(n_918),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_796),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_923),
.B(n_926),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_842),
.A2(n_866),
.B(n_893),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_916),
.B(n_929),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_917),
.A2(n_861),
.B(n_885),
.Y(n_958)
);

AO31x2_ASAP7_75t_L g959 ( 
.A1(n_938),
.A2(n_804),
.A3(n_801),
.B(n_875),
.Y(n_959)
);

AND3x4_ASAP7_75t_L g960 ( 
.A(n_910),
.B(n_895),
.C(n_914),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_819),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_944),
.B(n_939),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_908),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_822),
.A2(n_894),
.B(n_867),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_796),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_855),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_939),
.B(n_942),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_885),
.A2(n_872),
.B(n_933),
.C(n_937),
.Y(n_968)
);

AOI211x1_ASAP7_75t_L g969 ( 
.A1(n_942),
.A2(n_950),
.B(n_947),
.C(n_912),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_871),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_941),
.B(n_949),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_863),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_947),
.A2(n_950),
.B1(n_946),
.B2(n_928),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_864),
.B(n_800),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_814),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_928),
.A2(n_946),
.B1(n_859),
.B2(n_844),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_868),
.B(n_888),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_936),
.B(n_943),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_859),
.A2(n_900),
.B1(n_912),
.B2(n_823),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_806),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_920),
.B(n_930),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_934),
.A2(n_803),
.B(n_799),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_908),
.Y(n_983)
);

AO21x1_ASAP7_75t_L g984 ( 
.A1(n_877),
.A2(n_892),
.B(n_843),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_819),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_816),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_830),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_840),
.A2(n_899),
.B(n_873),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_945),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_SL g990 ( 
.A1(n_906),
.A2(n_898),
.B(n_896),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_890),
.A2(n_799),
.B(n_865),
.Y(n_991)
);

OAI21x1_ASAP7_75t_SL g992 ( 
.A1(n_879),
.A2(n_877),
.B(n_848),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_908),
.B(n_869),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_839),
.B(n_870),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_940),
.B(n_948),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_839),
.B(n_901),
.Y(n_996)
);

AOI21xp33_ASAP7_75t_L g997 ( 
.A1(n_795),
.A2(n_856),
.B(n_838),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_932),
.A2(n_802),
.B(n_807),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_817),
.B(n_909),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_819),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_902),
.B(n_903),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_845),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_821),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_845),
.B(n_925),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_883),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_887),
.A2(n_886),
.B(n_815),
.Y(n_1006)
);

O2A1O1Ixp5_ASAP7_75t_L g1007 ( 
.A1(n_879),
.A2(n_820),
.B(n_904),
.C(n_812),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_882),
.A2(n_813),
.B(n_860),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_795),
.A2(n_882),
.B(n_818),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_820),
.A2(n_797),
.B(n_812),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_895),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_845),
.B(n_925),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_925),
.B(n_935),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_909),
.B(n_805),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_924),
.A2(n_897),
.B1(n_891),
.B2(n_936),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_811),
.A2(n_905),
.B(n_831),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_810),
.A2(n_831),
.B(n_837),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_825),
.B(n_829),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_878),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_874),
.B(n_853),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_808),
.B(n_834),
.Y(n_1021)
);

BUFx4f_ASAP7_75t_SL g1022 ( 
.A(n_911),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_915),
.A2(n_833),
.B(n_841),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_835),
.Y(n_1024)
);

AND2x6_ASAP7_75t_L g1025 ( 
.A(n_798),
.B(n_809),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_833),
.A2(n_851),
.B(n_858),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_826),
.A2(n_927),
.B(n_919),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_828),
.A2(n_889),
.B(n_905),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_935),
.B(n_810),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_827),
.A2(n_913),
.B(n_836),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_849),
.B(n_850),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_827),
.A2(n_852),
.B(n_846),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_854),
.B(n_881),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_854),
.B(n_881),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_857),
.A2(n_847),
.B(n_832),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_931),
.A2(n_832),
.B(n_907),
.C(n_911),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_931),
.A2(n_842),
.B(n_866),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_855),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_819),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_842),
.A2(n_866),
.B(n_893),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_824),
.A2(n_862),
.B(n_885),
.C(n_872),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_842),
.A2(n_866),
.B(n_893),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_916),
.B(n_918),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_R g1044 ( 
.A(n_821),
.B(n_483),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_936),
.B(n_943),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_L g1046 ( 
.A1(n_932),
.A2(n_721),
.B(n_802),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_824),
.B(n_884),
.Y(n_1047)
);

AND3x2_ASAP7_75t_L g1048 ( 
.A(n_824),
.B(n_505),
.C(n_658),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_916),
.B(n_918),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_842),
.A2(n_866),
.B(n_893),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_824),
.A2(n_862),
.B(n_885),
.C(n_872),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_916),
.B(n_918),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_842),
.A2(n_866),
.B(n_893),
.Y(n_1053)
);

OAI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_824),
.A2(n_731),
.B(n_730),
.Y(n_1054)
);

AOI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_824),
.A2(n_884),
.B(n_872),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_923),
.B(n_697),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_923),
.B(n_697),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_819),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_916),
.B(n_918),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_819),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_923),
.B(n_697),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_916),
.B(n_918),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_819),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_842),
.A2(n_866),
.B(n_893),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_819),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_938),
.A2(n_804),
.A3(n_862),
.B(n_801),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_819),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_814),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_814),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_917),
.A2(n_862),
.B(n_824),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_824),
.B(n_916),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_L g1072 ( 
.A1(n_824),
.A2(n_885),
.B(n_884),
.C(n_862),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_819),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_916),
.B(n_918),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_916),
.B(n_918),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_806),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_824),
.A2(n_862),
.B(n_885),
.C(n_872),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_824),
.A2(n_731),
.B(n_730),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_SL g1079 ( 
.A1(n_939),
.A2(n_950),
.B(n_947),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_917),
.A2(n_862),
.B(n_824),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_824),
.B(n_884),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_938),
.A2(n_804),
.A3(n_862),
.B(n_801),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_980),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_1001),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1068),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_961),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_978),
.B(n_1045),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1056),
.B(n_1057),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_978),
.B(n_1045),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_1011),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_1001),
.Y(n_1091)
);

INVx5_ASAP7_75t_L g1092 ( 
.A(n_1004),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_963),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_967),
.B(n_1071),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_1068),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_967),
.B(n_1071),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_SL g1097 ( 
.A1(n_968),
.A2(n_1080),
.B(n_1070),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1061),
.B(n_955),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1004),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1076),
.Y(n_1100)
);

AO21x2_ASAP7_75t_L g1101 ( 
.A1(n_992),
.A2(n_958),
.B(n_1070),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_961),
.Y(n_1102)
);

AND2x6_ASAP7_75t_L g1103 ( 
.A(n_1015),
.B(n_1029),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_972),
.Y(n_1104)
);

OR2x6_ASAP7_75t_L g1105 ( 
.A(n_1004),
.B(n_983),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_957),
.B(n_1043),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1002),
.B(n_1058),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_993),
.B(n_1002),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_974),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1024),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_971),
.B(n_1014),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1038),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_958),
.A2(n_1080),
.B(n_982),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1049),
.B(n_1059),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_975),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_970),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_952),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1054),
.B(n_1078),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1052),
.B(n_1062),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1005),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_979),
.A2(n_1055),
.B1(n_951),
.B2(n_1047),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_953),
.B(n_1081),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_1051),
.B1(n_1077),
.B2(n_979),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_961),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_987),
.B(n_1022),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1003),
.Y(n_1127)
);

BUFx8_ASAP7_75t_L g1128 ( 
.A(n_999),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1058),
.B(n_1060),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_1069),
.B(n_986),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1079),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_985),
.Y(n_1132)
);

CKINVDCx11_ASAP7_75t_R g1133 ( 
.A(n_1069),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_986),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_962),
.B(n_1055),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1060),
.B(n_1063),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1063),
.B(n_1067),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1018),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_985),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_1013),
.B(n_1033),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_981),
.A2(n_995),
.B1(n_969),
.B2(n_973),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_973),
.B(n_1020),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_996),
.B(n_976),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_985),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1021),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_994),
.A2(n_960),
.B1(n_977),
.B2(n_1034),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_954),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_990),
.B(n_1048),
.Y(n_1148)
);

CKINVDCx16_ASAP7_75t_R g1149 ( 
.A(n_1000),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1072),
.B(n_1013),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_997),
.A2(n_1030),
.B(n_982),
.C(n_976),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1000),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_997),
.B(n_989),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1026),
.A2(n_1023),
.B1(n_984),
.B2(n_1030),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1026),
.A2(n_1023),
.B1(n_1032),
.B2(n_1010),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1039),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_1039),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1039),
.B(n_1073),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_965),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1065),
.B(n_1073),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1019),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1065),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1032),
.A2(n_1010),
.B1(n_1036),
.B2(n_1009),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1009),
.A2(n_1016),
.B1(n_1017),
.B2(n_1031),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1073),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_989),
.B(n_1012),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1017),
.A2(n_1019),
.B1(n_1028),
.B2(n_1027),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1025),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1025),
.B(n_1082),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1025),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1066),
.B(n_1082),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1037),
.A2(n_1035),
.B1(n_1008),
.B2(n_964),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1044),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_959),
.Y(n_1174)
);

AO21x1_ASAP7_75t_L g1175 ( 
.A1(n_1046),
.A2(n_1006),
.B(n_998),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_959),
.B(n_1064),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1007),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_956),
.A2(n_1040),
.B1(n_1042),
.B2(n_1050),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1053),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_980),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1054),
.A2(n_824),
.B1(n_1078),
.B2(n_885),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_980),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_SL g1183 ( 
.A(n_980),
.B(n_665),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_980),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_966),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_971),
.B(n_824),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1070),
.A2(n_824),
.B(n_1080),
.C(n_1054),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1071),
.A2(n_967),
.B1(n_1043),
.B2(n_957),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1056),
.B(n_1057),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_978),
.B(n_1045),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1054),
.A2(n_824),
.B1(n_1078),
.B2(n_885),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1052),
.B(n_1074),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1056),
.B(n_1057),
.Y(n_1193)
);

CKINVDCx16_ASAP7_75t_R g1194 ( 
.A(n_1003),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_980),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1052),
.B(n_1074),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_978),
.B(n_1045),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_961),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_963),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_SL g1201 ( 
.A(n_967),
.B(n_996),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1003),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_988),
.A2(n_884),
.B(n_991),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1071),
.A2(n_967),
.B1(n_1043),
.B2(n_957),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1056),
.B(n_1057),
.Y(n_1205)
);

AOI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1054),
.A2(n_824),
.B(n_1078),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1011),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_961),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_967),
.B(n_1071),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_966),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1068),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_967),
.B(n_1071),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_967),
.B(n_1071),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_980),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_966),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_978),
.B(n_1045),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1004),
.B(n_963),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_978),
.B(n_1045),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1150),
.B(n_1131),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1092),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1186),
.A2(n_1103),
.B1(n_1118),
.B2(n_1206),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1092),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1110),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1186),
.A2(n_1103),
.B1(n_1118),
.B2(n_1206),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1157),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1211),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1148),
.A2(n_1124),
.B1(n_1103),
.B2(n_1111),
.Y(n_1227)
);

BUFx2_ASAP7_75t_R g1228 ( 
.A(n_1083),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1210),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1109),
.B(n_1122),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1215),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1211),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_SL g1233 ( 
.A(n_1180),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1146),
.A2(n_1096),
.B1(n_1209),
.B2(n_1094),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1104),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1112),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1106),
.B(n_1114),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1202),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1185),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1134),
.Y(n_1240)
);

BUFx8_ASAP7_75t_L g1241 ( 
.A(n_1093),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1085),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1128),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1103),
.A2(n_1191),
.B1(n_1181),
.B2(n_1148),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1106),
.B(n_1114),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1095),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1116),
.Y(n_1247)
);

CKINVDCx11_ASAP7_75t_R g1248 ( 
.A(n_1195),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1108),
.B(n_1140),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1128),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1103),
.A2(n_1181),
.B1(n_1191),
.B2(n_1124),
.Y(n_1251)
);

BUFx2_ASAP7_75t_SL g1252 ( 
.A(n_1092),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1130),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1122),
.B(n_1094),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1098),
.A2(n_1142),
.B1(n_1163),
.B2(n_1155),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1187),
.A2(n_1154),
.B(n_1155),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1120),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1133),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1096),
.B(n_1209),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1125),
.Y(n_1261)
);

BUFx2_ASAP7_75t_R g1262 ( 
.A(n_1182),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1115),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1121),
.B(n_1119),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1138),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1125),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1194),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1125),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1105),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1188),
.A2(n_1204),
.B1(n_1187),
.B2(n_1142),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1135),
.B(n_1123),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1177),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1145),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1125),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1147),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1088),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1135),
.B(n_1123),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1163),
.A2(n_1154),
.B1(n_1143),
.B2(n_1205),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1201),
.B(n_1171),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1143),
.A2(n_1189),
.B1(n_1193),
.B2(n_1113),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1203),
.A2(n_1151),
.B(n_1178),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1183),
.A2(n_1164),
.B1(n_1196),
.B2(n_1192),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1153),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1159),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1113),
.A2(n_1141),
.B1(n_1164),
.B2(n_1101),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1127),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1176),
.B(n_1174),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1167),
.A2(n_1179),
.B(n_1175),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1140),
.A2(n_1090),
.B1(n_1207),
.B2(n_1105),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1141),
.A2(n_1100),
.B1(n_1184),
.B2(n_1214),
.Y(n_1291)
);

BUFx4f_ASAP7_75t_SL g1292 ( 
.A(n_1117),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1161),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1153),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1165),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1101),
.A2(n_1108),
.B1(n_1097),
.B2(n_1099),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1166),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1158),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1105),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1217),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1217),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1167),
.A2(n_1172),
.B(n_1169),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1140),
.B(n_1084),
.Y(n_1303)
);

BUFx2_ASAP7_75t_R g1304 ( 
.A(n_1162),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1151),
.B(n_1084),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1091),
.B(n_1198),
.Y(n_1306)
);

INVx6_ASAP7_75t_L g1307 ( 
.A(n_1149),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1091),
.B(n_1198),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1170),
.A2(n_1144),
.B(n_1156),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1099),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1168),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1160),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1086),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1200),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1087),
.A2(n_1218),
.B1(n_1089),
.B2(n_1197),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1107),
.A2(n_1217),
.B(n_1152),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1086),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1218),
.A2(n_1216),
.B1(n_1087),
.B2(n_1089),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_1107),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1086),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1102),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1102),
.Y(n_1322)
);

AO21x2_ASAP7_75t_L g1323 ( 
.A1(n_1160),
.A2(n_1129),
.B(n_1136),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1102),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1132),
.Y(n_1325)
);

BUFx2_ASAP7_75t_SL g1326 ( 
.A(n_1136),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1132),
.Y(n_1327)
);

BUFx2_ASAP7_75t_R g1328 ( 
.A(n_1139),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1152),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1199),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1190),
.A2(n_1197),
.B1(n_1216),
.B2(n_1126),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1137),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1208),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1137),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1190),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1173),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1211),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1337),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1337),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1237),
.B(n_1245),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1242),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1232),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1221),
.A2(n_1224),
.B(n_1271),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1272),
.B(n_1278),
.Y(n_1344)
);

INVxp33_ASAP7_75t_L g1345 ( 
.A(n_1240),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1272),
.B(n_1278),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1273),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1264),
.B(n_1260),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1289),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1253),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1283),
.A2(n_1251),
.B(n_1244),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1260),
.B(n_1268),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1282),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1282),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1234),
.B(n_1227),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1302),
.A2(n_1254),
.B(n_1286),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1253),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1255),
.B(n_1268),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1284),
.B(n_1294),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1257),
.A2(n_1302),
.B(n_1230),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1230),
.A2(n_1255),
.B(n_1305),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1288),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1288),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1226),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1256),
.A2(n_1279),
.B(n_1291),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1219),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1219),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1281),
.A2(n_1305),
.B(n_1280),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1297),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1280),
.A2(n_1265),
.B(n_1276),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1270),
.B(n_1299),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1235),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1309),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1236),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1239),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1277),
.A2(n_1274),
.B(n_1296),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1309),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1285),
.A2(n_1290),
.B(n_1300),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1263),
.B(n_1247),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1316),
.A2(n_1220),
.B(n_1222),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1303),
.B(n_1301),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1249),
.B(n_1220),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1246),
.Y(n_1383)
);

AO21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1223),
.A2(n_1231),
.B(n_1229),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1249),
.B(n_1220),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1249),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1298),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1314),
.B(n_1258),
.Y(n_1388)
);

CKINVDCx8_ASAP7_75t_R g1389 ( 
.A(n_1326),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1293),
.A2(n_1306),
.B(n_1308),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1252),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1323),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1319),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1331),
.A2(n_1336),
.B1(n_1335),
.B2(n_1315),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1241),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1311),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1310),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1310),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1334),
.B(n_1312),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1332),
.B(n_1312),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1355),
.B(n_1376),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1370),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1361),
.B(n_1320),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1320),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1370),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1361),
.B(n_1325),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1361),
.B(n_1325),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1360),
.B(n_1336),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1380),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1356),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1358),
.B(n_1330),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1358),
.B(n_1330),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1392),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1360),
.B(n_1322),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1373),
.B(n_1225),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1370),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1368),
.B(n_1370),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1368),
.B(n_1329),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1368),
.B(n_1327),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1368),
.B(n_1390),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1390),
.B(n_1324),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1390),
.B(n_1321),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1344),
.B(n_1333),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1390),
.B(n_1317),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1384),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1377),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1346),
.B(n_1313),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1346),
.B(n_1313),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1353),
.B(n_1225),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1377),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1354),
.B(n_1295),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1349),
.B(n_1295),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1395),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1356),
.B(n_1295),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1394),
.B(n_1307),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1401),
.A2(n_1343),
.B1(n_1351),
.B2(n_1365),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1415),
.B(n_1350),
.Y(n_1437)
);

OAI21xp33_ASAP7_75t_L g1438 ( 
.A1(n_1401),
.A2(n_1365),
.B(n_1343),
.Y(n_1438)
);

NOR3xp33_ASAP7_75t_L g1439 ( 
.A(n_1435),
.B(n_1340),
.C(n_1398),
.Y(n_1439)
);

AND2x2_ASAP7_75t_SL g1440 ( 
.A(n_1417),
.B(n_1386),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1415),
.B(n_1357),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1435),
.B(n_1394),
.C(n_1341),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1429),
.A2(n_1381),
.B1(n_1386),
.B2(n_1385),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1403),
.B(n_1362),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1434),
.A2(n_1259),
.B(n_1345),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1415),
.B(n_1342),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1429),
.B(n_1338),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1403),
.B(n_1362),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1429),
.A2(n_1381),
.B1(n_1385),
.B2(n_1382),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1408),
.B(n_1383),
.C(n_1369),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1408),
.B(n_1388),
.C(n_1371),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1411),
.B(n_1348),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1411),
.B(n_1352),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1408),
.A2(n_1318),
.B1(n_1371),
.B2(n_1379),
.C(n_1388),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1433),
.A2(n_1238),
.B1(n_1389),
.B2(n_1287),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1412),
.B(n_1339),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1420),
.A2(n_1364),
.B(n_1387),
.Y(n_1457)
);

AND4x1_ASAP7_75t_L g1458 ( 
.A(n_1434),
.B(n_1398),
.C(n_1397),
.D(n_1391),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1433),
.A2(n_1389),
.B1(n_1328),
.B2(n_1307),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1404),
.B(n_1363),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1412),
.B(n_1339),
.Y(n_1461)
);

OA211x2_ASAP7_75t_L g1462 ( 
.A1(n_1425),
.A2(n_1359),
.B(n_1399),
.C(n_1267),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_L g1463 ( 
.A(n_1431),
.B(n_1396),
.C(n_1372),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1431),
.B(n_1372),
.C(n_1347),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1423),
.B(n_1374),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1434),
.A2(n_1380),
.B(n_1400),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1406),
.B(n_1363),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1425),
.A2(n_1307),
.B1(n_1393),
.B2(n_1381),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1423),
.B(n_1427),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1406),
.B(n_1366),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1427),
.B(n_1374),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1409),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1428),
.B(n_1374),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1407),
.B(n_1366),
.Y(n_1474)
);

AND2x2_ASAP7_75t_SL g1475 ( 
.A(n_1417),
.B(n_1367),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1402),
.A2(n_1416),
.B(n_1405),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1420),
.A2(n_1382),
.B(n_1385),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1418),
.B(n_1419),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1428),
.B(n_1375),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1476),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1479),
.B(n_1417),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1476),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1438),
.B(n_1431),
.C(n_1414),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1476),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1479),
.B(n_1420),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1478),
.B(n_1421),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1478),
.B(n_1421),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1476),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1451),
.B(n_1421),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1444),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1451),
.B(n_1465),
.Y(n_1492)
);

NAND4xp25_ASAP7_75t_L g1493 ( 
.A(n_1436),
.B(n_1243),
.C(n_1250),
.D(n_1414),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1472),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1475),
.B(n_1418),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1475),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1475),
.B(n_1418),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1469),
.B(n_1422),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1440),
.B(n_1419),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1471),
.B(n_1422),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1444),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1448),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1440),
.B(n_1419),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1448),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1440),
.B(n_1426),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1437),
.B(n_1413),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1464),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1466),
.B(n_1430),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1472),
.B(n_1430),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1441),
.B(n_1413),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1473),
.B(n_1422),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1472),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1460),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1460),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1467),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1502),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1492),
.B(n_1453),
.Y(n_1517)
);

AND2x4_ASAP7_75t_SL g1518 ( 
.A(n_1505),
.B(n_1439),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1507),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1502),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1523)
);

AND2x4_ASAP7_75t_SL g1524 ( 
.A(n_1505),
.B(n_1432),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1507),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1495),
.B(n_1477),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1491),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1501),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1498),
.B(n_1452),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1495),
.B(n_1477),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1501),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1533)
);

CKINVDCx16_ASAP7_75t_R g1534 ( 
.A(n_1505),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1490),
.B(n_1480),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1504),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1500),
.B(n_1457),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1506),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1504),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1513),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1513),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1514),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1487),
.B(n_1456),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1496),
.B(n_1458),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1506),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1485),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1514),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1515),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_L g1550 ( 
.A1(n_1484),
.A2(n_1438),
.B(n_1457),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1484),
.A2(n_1445),
.B(n_1442),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1508),
.Y(n_1553)
);

NAND4xp25_ASAP7_75t_L g1554 ( 
.A(n_1493),
.B(n_1442),
.C(n_1462),
.D(n_1454),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1518),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1528),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1487),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1529),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1525),
.B(n_1488),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1534),
.B(n_1497),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1553),
.B(n_1508),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1524),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1520),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1535),
.B(n_1488),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1522),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1510),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1526),
.B(n_1531),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1536),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1547),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1547),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1533),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1540),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1552),
.A2(n_1493),
.B(n_1459),
.C(n_1445),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1541),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1543),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1517),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1546),
.B(n_1527),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

AOI32xp33_ASAP7_75t_L g1586 ( 
.A1(n_1550),
.A2(n_1518),
.A3(n_1531),
.B1(n_1496),
.B2(n_1553),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1524),
.B(n_1499),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1527),
.B(n_1510),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1530),
.B(n_1499),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1516),
.Y(n_1590)
);

AOI21xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1545),
.A2(n_1455),
.B(n_1508),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1533),
.B(n_1503),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1542),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1554),
.B(n_1228),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1542),
.B(n_1503),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1538),
.A2(n_1462),
.B1(n_1455),
.B2(n_1508),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1537),
.B(n_1503),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1559),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1572),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1563),
.B(n_1545),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

INVx3_ASAP7_75t_SL g1602 ( 
.A(n_1556),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1584),
.B(n_1544),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1557),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1566),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1560),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1584),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1570),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1564),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1594),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1564),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1563),
.B(n_1545),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

CKINVDCx16_ASAP7_75t_R g1616 ( 
.A(n_1596),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1544),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1561),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1568),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1573),
.B(n_1551),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1597),
.B(n_1523),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1486),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1571),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1588),
.B(n_1511),
.Y(n_1625)
);

CKINVDCx16_ASAP7_75t_R g1626 ( 
.A(n_1587),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1589),
.B(n_1569),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1591),
.B(n_1458),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1586),
.A2(n_1508),
.B(n_1238),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1558),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1569),
.B(n_1511),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1574),
.Y(n_1633)
);

NOR4xp25_ASAP7_75t_L g1634 ( 
.A(n_1609),
.B(n_1558),
.C(n_1562),
.D(n_1583),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1616),
.A2(n_1565),
.B1(n_1450),
.B2(n_1562),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1592),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1599),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1615),
.C(n_1630),
.Y(n_1640)
);

AO22x1_ASAP7_75t_L g1641 ( 
.A1(n_1612),
.A2(n_1564),
.B1(n_1565),
.B2(n_1595),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1610),
.Y(n_1642)
);

OAI21xp33_ASAP7_75t_L g1643 ( 
.A1(n_1623),
.A2(n_1629),
.B(n_1606),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1600),
.A2(n_1614),
.B1(n_1626),
.B2(n_1627),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1601),
.Y(n_1645)
);

OAI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1631),
.A2(n_1600),
.B1(n_1614),
.B2(n_1608),
.C(n_1603),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1620),
.B(n_1595),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1611),
.A2(n_1580),
.B(n_1578),
.Y(n_1648)
);

NAND4xp25_ASAP7_75t_SL g1649 ( 
.A(n_1620),
.B(n_1577),
.C(n_1593),
.D(n_1567),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1621),
.B(n_1577),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1604),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1621),
.B(n_1619),
.Y(n_1652)
);

OAI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1628),
.A2(n_1567),
.B(n_1593),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1611),
.A2(n_1585),
.B(n_1581),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1624),
.B(n_1486),
.Y(n_1655)
);

AO22x1_ASAP7_75t_L g1656 ( 
.A1(n_1611),
.A2(n_1576),
.B1(n_1575),
.B2(n_1243),
.Y(n_1656)
);

OAI32xp33_ASAP7_75t_L g1657 ( 
.A1(n_1613),
.A2(n_1481),
.A3(n_1576),
.B1(n_1575),
.B2(n_1485),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1613),
.A2(n_1287),
.B(n_1450),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1605),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1637),
.B(n_1617),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1642),
.B(n_1633),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1638),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1639),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1642),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1640),
.B(n_1613),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1643),
.B(n_1644),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1607),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1645),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1651),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1652),
.B(n_1617),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1627),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1641),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1635),
.B(n_1622),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1649),
.A2(n_1653),
.B1(n_1635),
.B2(n_1658),
.Y(n_1675)
);

AND2x4_ASAP7_75t_SL g1676 ( 
.A(n_1647),
.B(n_1659),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1618),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1655),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1665),
.A2(n_1654),
.B(n_1657),
.Y(n_1681)
);

NAND4xp25_ASAP7_75t_L g1682 ( 
.A(n_1666),
.B(n_1250),
.C(n_1632),
.D(n_1625),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1674),
.A2(n_1656),
.B(n_1632),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1664),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1673),
.B(n_1625),
.Y(n_1685)
);

NOR4xp25_ASAP7_75t_L g1686 ( 
.A(n_1672),
.B(n_1485),
.C(n_1267),
.D(n_1483),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1667),
.B(n_1241),
.C(n_1248),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1675),
.A2(n_1432),
.B1(n_1424),
.B2(n_1468),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_L g1689 ( 
.A(n_1663),
.B(n_1432),
.C(n_1449),
.D(n_1443),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_SL g1690 ( 
.A1(n_1667),
.A2(n_1307),
.B1(n_1410),
.B2(n_1241),
.Y(n_1690)
);

AOI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1680),
.A2(n_1481),
.B(n_1494),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1685),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1681),
.B(n_1687),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1660),
.Y(n_1694)
);

AOI211x1_ASAP7_75t_L g1695 ( 
.A1(n_1683),
.A2(n_1682),
.B(n_1671),
.C(n_1661),
.Y(n_1695)
);

NOR3xp33_ASAP7_75t_L g1696 ( 
.A(n_1690),
.B(n_1661),
.C(n_1678),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1691),
.Y(n_1697)
);

NOR3xp33_ASAP7_75t_L g1698 ( 
.A(n_1688),
.B(n_1677),
.C(n_1669),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1686),
.B(n_1670),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1689),
.Y(n_1700)
);

NAND4xp75_ASAP7_75t_L g1701 ( 
.A(n_1681),
.B(n_1677),
.C(n_1668),
.D(n_1662),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1699),
.A2(n_1676),
.B(n_1679),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1693),
.A2(n_1262),
.B(n_1233),
.Y(n_1703)
);

NAND2xp33_ASAP7_75t_R g1704 ( 
.A(n_1694),
.B(n_1248),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1692),
.B(n_1486),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1701),
.B(n_1292),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1698),
.A2(n_1463),
.B(n_1397),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1705),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1706),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1704),
.A2(n_1696),
.B1(n_1700),
.B2(n_1697),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1702),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1707),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1703),
.A2(n_1695),
.B1(n_1424),
.B2(n_1509),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1706),
.Y(n_1714)
);

AND3x4_ASAP7_75t_L g1715 ( 
.A(n_1714),
.B(n_1304),
.C(n_1509),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1709),
.B(n_1482),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1711),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1708),
.B(n_1482),
.Y(n_1718)
);

NOR3xp33_ASAP7_75t_SL g1719 ( 
.A(n_1712),
.B(n_1463),
.C(n_1461),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1717),
.B(n_1710),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_L g1721 ( 
.A(n_1719),
.B(n_1713),
.C(n_1275),
.Y(n_1721)
);

AND3x4_ASAP7_75t_L g1722 ( 
.A(n_1716),
.B(n_1718),
.C(n_1715),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1720),
.Y(n_1723)
);

O2A1O1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1721),
.B(n_1722),
.C(n_1485),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1724),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1724),
.B(n_1266),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1512),
.B1(n_1509),
.B2(n_1494),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1726),
.A2(n_1261),
.B1(n_1269),
.B2(n_1266),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1728),
.Y(n_1729)
);

AOI21xp33_ASAP7_75t_L g1730 ( 
.A1(n_1727),
.A2(n_1269),
.B(n_1261),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1729),
.B(n_1482),
.Y(n_1731)
);

AOI322xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1730),
.A3(n_1512),
.B1(n_1494),
.B2(n_1483),
.C1(n_1489),
.C2(n_1509),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1489),
.B1(n_1512),
.B2(n_1275),
.C(n_1266),
.Y(n_1733)
);

AOI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1266),
.B(n_1275),
.C(n_1391),
.Y(n_1734)
);


endmodule