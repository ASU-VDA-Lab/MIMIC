module fake_jpeg_21830_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_7),
.A2(n_9),
.B1(n_10),
.B2(n_6),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_17),
.B1(n_9),
.B2(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_10),
.C(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_21),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_13),
.C(n_17),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_25),
.B(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_6),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_19),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_19),
.C(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_11),
.Y(n_34)
);

OAI211xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B(n_12),
.C(n_4),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_30),
.C(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NAND4xp25_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_14),
.C(n_20),
.D(n_36),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_20),
.Y(n_39)
);


endmodule