module fake_netlist_6_1933_n_1779 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1779);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1779;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_71),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_63),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_1),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_18),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

BUFx2_ASAP7_75t_SL g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_55),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_34),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_34),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_120),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_51),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_42),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_62),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_10),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_79),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_132),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_32),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_22),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_27),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_98),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_17),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_22),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_3),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_70),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_119),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_58),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_20),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_18),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_21),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_45),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_52),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_1),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_116),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_96),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_64),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_83),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_9),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_117),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_140),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_23),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_16),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_61),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_3),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_48),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_146),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_102),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_35),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_47),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_109),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_26),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_59),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_57),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_41),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_138),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_33),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_95),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_137),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_7),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_39),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_106),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_133),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_80),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_43),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_65),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_13),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_20),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_91),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_5),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_8),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_39),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_121),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_136),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_130),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_41),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_60),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_50),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_53),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_93),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_100),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_105),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_21),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_69),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_87),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_86),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_77),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_42),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_124),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_6),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_25),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_30),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_50),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_49),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_6),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_13),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_104),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_54),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_56),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_38),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_46),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_12),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_40),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_67),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_44),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_188),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_212),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_213),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_188),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_188),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_188),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_201),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_188),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_160),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_224),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_155),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_202),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_155),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_160),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_203),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_209),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_215),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_217),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_186),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_186),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_0),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_206),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_252),
.B(n_0),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_162),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_221),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_175),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_175),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_229),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_2),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_233),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_195),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_239),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_178),
.B(n_4),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_161),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_196),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_181),
.B(n_5),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_244),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_222),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_190),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_207),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_223),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_208),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_162),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_161),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_208),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_245),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_191),
.B(n_7),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_231),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_248),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_161),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_253),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_255),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_181),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_256),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_238),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_261),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_262),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_241),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_219),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_259),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_219),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_194),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_341),
.B(n_156),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_191),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_156),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_198),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_314),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_314),
.B(n_198),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_214),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_159),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_316),
.B(n_214),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_320),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_265),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_360),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_333),
.B(n_190),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_333),
.B(n_337),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_331),
.B(n_265),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

OR2x6_ASAP7_75t_L g432 ( 
.A(n_337),
.B(n_164),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_350),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g434 ( 
.A(n_368),
.B(n_298),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_355),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_331),
.B(n_159),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_319),
.B(n_200),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_332),
.B(n_168),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_361),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_348),
.B(n_298),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_317),
.B(n_272),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_369),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_448),
.A2(n_352),
.B1(n_327),
.B2(n_345),
.Y(n_453)
);

NOR2x1p5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_318),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_321),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_442),
.B(n_360),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_416),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_392),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_328),
.C(n_325),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_433),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_392),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_417),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_436),
.B(n_329),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_436),
.B(n_330),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_392),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

BUFx8_ASAP7_75t_SL g478 ( 
.A(n_439),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_397),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_222),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_434),
.A2(n_336),
.B1(n_353),
.B2(n_324),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_433),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_399),
.B(n_339),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_408),
.B(n_376),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_392),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_417),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_379),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_440),
.B(n_358),
.C(n_349),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_434),
.A2(n_338),
.B1(n_300),
.B2(n_293),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_399),
.B(n_370),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_439),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_439),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_443),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_384),
.B(n_372),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_388),
.B(n_399),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_443),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_384),
.B(n_373),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_399),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_447),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_434),
.A2(n_304),
.B1(n_263),
.B2(n_264),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_391),
.B(n_375),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_391),
.B(n_377),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_399),
.B(n_378),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_409),
.B(n_315),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_400),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_409),
.B(n_367),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_400),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_410),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_447),
.Y(n_524)
);

BUFx6f_ASAP7_75t_SL g525 ( 
.A(n_446),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_428),
.B(n_363),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_449),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_388),
.B(n_234),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_404),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_390),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_404),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_425),
.B(n_366),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_444),
.B(n_379),
.C(n_334),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_404),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_428),
.B(n_351),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_388),
.B(n_157),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_444),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_414),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_425),
.B(n_190),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_408),
.B(n_222),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_408),
.B(n_421),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_390),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_449),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_421),
.B(n_351),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_414),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_407),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_410),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_446),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_424),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_386),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_410),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_386),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_421),
.B(n_332),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_446),
.B(n_222),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_386),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_446),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_410),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_429),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_446),
.B(n_158),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_424),
.B(n_334),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_387),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_424),
.B(n_335),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_414),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_424),
.B(n_335),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_405),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_432),
.B(n_340),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_405),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_434),
.A2(n_290),
.B1(n_296),
.B2(n_271),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_407),
.Y(n_577)
);

INVx8_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_387),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_446),
.B(n_168),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_414),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_387),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_434),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_431),
.B(n_171),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_394),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_452),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_431),
.B(n_171),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_434),
.B(n_163),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_394),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_429),
.B(n_309),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_434),
.A2(n_310),
.B1(n_312),
.B2(n_270),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_432),
.B(n_340),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_434),
.B(n_165),
.Y(n_594)
);

BUFx6f_ASAP7_75t_SL g595 ( 
.A(n_432),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_401),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_401),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_407),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_434),
.B(n_166),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_429),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_452),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_549),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_466),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_542),
.B(n_432),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_499),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_SL g607 ( 
.A(n_555),
.B(n_564),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_455),
.B(n_526),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_515),
.B(n_434),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_555),
.B(n_432),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_564),
.A2(n_432),
.B1(n_179),
.B2(n_176),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_488),
.B(n_343),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_499),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_566),
.B(n_600),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_466),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_470),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_504),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_583),
.B(n_222),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_504),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_343),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_458),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_517),
.A2(n_432),
.B1(n_270),
.B2(n_189),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_470),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_462),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_552),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_493),
.B(n_187),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_552),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_546),
.B(n_407),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_601),
.B(n_407),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_472),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_411),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_501),
.Y(n_633)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_560),
.A2(n_205),
.B(n_211),
.C(n_273),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_553),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_583),
.B(n_267),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_501),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_459),
.A2(n_413),
.B(n_405),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_568),
.B(n_411),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_484),
.B(n_381),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_577),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_463),
.B(n_346),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_570),
.B(n_411),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_572),
.B(n_573),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_501),
.B(n_411),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_549),
.B(n_346),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_501),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_556),
.B(n_267),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_598),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_598),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_469),
.B(n_288),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_501),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_541),
.A2(n_430),
.B(n_450),
.C(n_445),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_472),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_467),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_519),
.B(n_172),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_556),
.B(n_267),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_479),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_467),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_599),
.B(n_267),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_475),
.A2(n_413),
.B(n_405),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_476),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_523),
.A2(n_492),
.B(n_483),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_484),
.B(n_533),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_479),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_501),
.B(n_464),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_476),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_547),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_456),
.B(n_172),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_589),
.B(n_267),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_594),
.B(n_161),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_453),
.B(n_422),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_484),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_465),
.B(n_411),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_486),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_460),
.B(n_381),
.C(n_220),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_547),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_491),
.A2(n_411),
.B1(n_282),
.B2(n_161),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_463),
.B(n_208),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_516),
.B(n_174),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_525),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_482),
.B(n_431),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_469),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_574),
.B(n_161),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_578),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_495),
.B(n_431),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_490),
.B(n_422),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_486),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_575),
.B(n_161),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_497),
.B(n_502),
.Y(n_691)
);

INVx8_ASAP7_75t_L g692 ( 
.A(n_489),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_514),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_496),
.B(n_174),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_514),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_557),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_503),
.B(n_177),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_591),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_481),
.B(n_537),
.C(n_531),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_560),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_513),
.B(n_177),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_511),
.A2(n_161),
.B1(n_218),
.B2(n_277),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_575),
.B(n_431),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_575),
.B(n_431),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_591),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_471),
.B(n_182),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_557),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_506),
.B(n_431),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_498),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_527),
.B(n_431),
.Y(n_710)
);

AND2x4_ASAP7_75t_SL g711 ( 
.A(n_489),
.B(n_257),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_585),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_507),
.B(n_431),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_559),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_473),
.B(n_182),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_524),
.B(n_451),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_525),
.A2(n_301),
.B1(n_185),
.B2(n_184),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_530),
.B(n_451),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_494),
.Y(n_719)
);

AND2x4_ASAP7_75t_SL g720 ( 
.A(n_489),
.B(n_257),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_489),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_563),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_480),
.A2(n_435),
.B(n_450),
.C(n_445),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_498),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_527),
.B(n_562),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_505),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_578),
.A2(n_167),
.B1(n_173),
.B2(n_193),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_527),
.B(n_451),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_540),
.B(n_548),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_550),
.B(n_451),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_587),
.B(n_451),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_536),
.B(n_184),
.Y(n_732)
);

AO22x2_ASAP7_75t_L g733 ( 
.A1(n_544),
.A2(n_197),
.B1(n_210),
.B2(n_216),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_505),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_562),
.B(n_451),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_593),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_508),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_563),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_569),
.B(n_451),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_508),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_569),
.B(n_451),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_579),
.B(n_451),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_562),
.B(n_385),
.Y(n_743)
);

OR2x2_ASAP7_75t_SL g744 ( 
.A(n_592),
.B(n_240),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_567),
.B(n_385),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_494),
.B(n_257),
.Y(n_746)
);

BUFx6f_ASAP7_75t_SL g747 ( 
.A(n_478),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_579),
.B(n_405),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_580),
.B(n_185),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_582),
.B(n_405),
.Y(n_750)
);

AND3x1_ASAP7_75t_L g751 ( 
.A(n_576),
.B(n_249),
.C(n_286),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_478),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_512),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_480),
.A2(n_258),
.B1(n_268),
.B2(n_283),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_582),
.B(n_413),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_468),
.B(n_385),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_454),
.B(n_169),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_586),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_593),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_586),
.B(n_413),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_593),
.B(n_584),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_512),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_545),
.B(n_413),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_590),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_593),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_518),
.Y(n_766)
);

BUFx8_ASAP7_75t_L g767 ( 
.A(n_595),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_590),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_588),
.B(n_525),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_596),
.B(n_189),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_518),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_596),
.B(n_269),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_608),
.B(n_578),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_608),
.B(n_597),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_696),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_614),
.B(n_597),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_712),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_614),
.B(n_578),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_725),
.A2(n_487),
.B(n_485),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_725),
.A2(n_487),
.B(n_485),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_665),
.B(n_280),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_712),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_669),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_604),
.B(n_674),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_686),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_657),
.B(n_545),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_604),
.B(n_269),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_657),
.B(n_645),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_699),
.A2(n_285),
.B(n_289),
.C(n_509),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_640),
.A2(n_487),
.B(n_485),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_674),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_644),
.A2(n_554),
.B(n_529),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_670),
.A2(n_509),
.B(n_457),
.C(n_500),
.Y(n_793)
);

AO21x1_ASAP7_75t_L g794 ( 
.A1(n_685),
.A2(n_554),
.B(n_529),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_700),
.B(n_275),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_605),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_643),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_664),
.A2(n_554),
.B(n_529),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_646),
.A2(n_468),
.B(n_477),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_670),
.A2(n_509),
.B(n_457),
.C(n_500),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_710),
.A2(n_468),
.B(n_477),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_653),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_681),
.B(n_545),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_609),
.A2(n_457),
.B(n_474),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_752),
.B(n_595),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_681),
.B(n_545),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_710),
.A2(n_558),
.B(n_468),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_634),
.A2(n_445),
.B(n_438),
.C(n_441),
.Y(n_809)
);

O2A1O1Ixp5_ASAP7_75t_L g810 ( 
.A1(n_685),
.A2(n_500),
.B(n_474),
.C(n_571),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_629),
.B(n_545),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_686),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_728),
.A2(n_477),
.B(n_468),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_678),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_749),
.A2(n_474),
.B(n_581),
.C(n_571),
.Y(n_815)
);

OAI21xp33_ASAP7_75t_L g816 ( 
.A1(n_706),
.A2(n_292),
.B(n_291),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_656),
.B(n_545),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_660),
.B(n_477),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_714),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_761),
.A2(n_595),
.B1(n_561),
.B2(n_558),
.Y(n_820)
);

BUFx8_ASAP7_75t_L g821 ( 
.A(n_747),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_700),
.B(n_275),
.Y(n_822)
);

O2A1O1Ixp5_ASAP7_75t_L g823 ( 
.A1(n_649),
.A2(n_528),
.B(n_521),
.C(n_522),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_728),
.A2(n_477),
.B(n_558),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_735),
.A2(n_558),
.B(n_565),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_686),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_722),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_761),
.A2(n_561),
.B1(n_558),
.B2(n_278),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_643),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_632),
.A2(n_653),
.B1(n_633),
.B2(n_648),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_634),
.A2(n_437),
.B(n_445),
.C(n_441),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_738),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_653),
.B(n_276),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_663),
.B(n_521),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_602),
.B(n_280),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_668),
.B(n_522),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_653),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_641),
.B(n_276),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_641),
.B(n_278),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_758),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_606),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_759),
.B(n_279),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_684),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_613),
.Y(n_845)
);

CKINVDCx10_ASAP7_75t_R g846 ( 
.A(n_747),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_279),
.C(n_281),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_689),
.B(n_528),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_618),
.A2(n_637),
.B(n_628),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_618),
.A2(n_581),
.B(n_532),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_617),
.Y(n_851)
);

NOR2x2_ASAP7_75t_L g852 ( 
.A(n_643),
.B(n_280),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_719),
.B(n_281),
.Y(n_853)
);

AO21x2_ASAP7_75t_L g854 ( 
.A1(n_610),
.A2(n_403),
.B(n_406),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_735),
.A2(n_565),
.B(n_461),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_743),
.A2(n_565),
.B(n_461),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_693),
.B(n_532),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_637),
.A2(n_430),
.B(n_435),
.C(n_437),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_619),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_695),
.B(n_534),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_686),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_621),
.B(n_624),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_SL g863 ( 
.A1(n_667),
.A2(n_534),
.B(n_535),
.C(n_538),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_652),
.B(n_169),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_694),
.B(n_697),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_649),
.A2(n_441),
.B(n_430),
.C(n_435),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_633),
.A2(n_306),
.B1(n_299),
.B2(n_287),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_658),
.A2(n_441),
.B(n_430),
.C(n_435),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_743),
.A2(n_565),
.B(n_461),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_764),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_697),
.B(n_199),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_638),
.A2(n_287),
.B1(n_301),
.B2(n_299),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_745),
.A2(n_565),
.B(n_461),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_692),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_SL g875 ( 
.A(n_701),
.B(n_306),
.C(n_170),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_647),
.B(n_620),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_745),
.A2(n_535),
.B(n_551),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_701),
.B(n_437),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_673),
.B(n_437),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_768),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_638),
.B(n_438),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_691),
.B(n_538),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_706),
.B(n_225),
.Y(n_883)
);

INVx3_ASAP7_75t_SL g884 ( 
.A(n_744),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_729),
.B(n_543),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_770),
.B(n_543),
.Y(n_886)
);

NOR2x2_ASAP7_75t_L g887 ( 
.A(n_612),
.B(n_297),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_770),
.B(n_551),
.Y(n_888)
);

BUFx8_ASAP7_75t_SL g889 ( 
.A(n_612),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_612),
.B(n_226),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_736),
.B(n_422),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_679),
.B(n_438),
.Y(n_892)
);

AO21x1_ASAP7_75t_L g893 ( 
.A1(n_658),
.A2(n_401),
.B(n_403),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_705),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_772),
.B(n_561),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_749),
.A2(n_385),
.B(n_389),
.C(n_426),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_625),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_715),
.A2(n_170),
.B(n_183),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_680),
.B(n_228),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_603),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_627),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_715),
.B(n_426),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_L g903 ( 
.A(n_692),
.B(n_561),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_702),
.A2(n_561),
.B1(n_297),
.B2(n_303),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_692),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_626),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_631),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_675),
.A2(n_520),
.B(n_510),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_639),
.A2(n_561),
.B(n_520),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_662),
.A2(n_520),
.B(n_510),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_615),
.Y(n_911)
);

AOI22x1_ASAP7_75t_L g912 ( 
.A1(n_635),
.A2(n_385),
.B1(n_389),
.B2(n_180),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_682),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_746),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_763),
.A2(n_520),
.B(n_510),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_756),
.A2(n_520),
.B(n_510),
.Y(n_916)
);

AOI21x1_ASAP7_75t_L g917 ( 
.A1(n_607),
.A2(n_406),
.B(n_403),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_732),
.B(n_230),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_732),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_772),
.B(n_438),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_736),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_756),
.A2(n_406),
.B(n_396),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_748),
.A2(n_510),
.B(n_461),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_688),
.B(n_450),
.Y(n_924)
);

BUFx4f_ASAP7_75t_L g925 ( 
.A(n_711),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_765),
.B(n_426),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_648),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_682),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_711),
.B(n_297),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_672),
.A2(n_450),
.B(n_427),
.C(n_420),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_616),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_622),
.B(n_415),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_767),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_767),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_636),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_750),
.A2(n_413),
.B(n_395),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_717),
.B(n_73),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_755),
.A2(n_395),
.B(n_385),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_698),
.B(n_243),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_642),
.B(n_389),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_765),
.B(n_415),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_760),
.A2(n_395),
.B(n_389),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_650),
.B(n_651),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_720),
.B(n_623),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_720),
.B(n_180),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_769),
.A2(n_389),
.B(n_415),
.C(n_420),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_769),
.A2(n_654),
.B(n_679),
.C(n_718),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_630),
.B(n_655),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_677),
.B(n_427),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_659),
.B(n_389),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_703),
.A2(n_395),
.B(n_396),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_666),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_703),
.A2(n_395),
.B(n_396),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_739),
.A2(n_396),
.B(n_415),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_683),
.A2(n_427),
.B(n_419),
.C(n_420),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_721),
.B(n_260),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_704),
.A2(n_427),
.B(n_420),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_721),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_704),
.A2(n_395),
.B(n_419),
.Y(n_959)
);

NOR2x1_ASAP7_75t_R g960 ( 
.A(n_690),
.B(n_291),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_796),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_865),
.B(n_733),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_SL g963 ( 
.A1(n_865),
.A2(n_733),
.B1(n_727),
.B2(n_611),
.Y(n_963)
);

O2A1O1Ixp5_ASAP7_75t_L g964 ( 
.A1(n_883),
.A2(n_671),
.B(n_661),
.C(n_716),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_894),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_810),
.A2(n_742),
.B(n_741),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_783),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_874),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_774),
.B(n_709),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_871),
.A2(n_723),
.B(n_730),
.C(n_731),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_781),
.B(n_757),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_871),
.A2(n_687),
.B(n_713),
.C(n_708),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_844),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_773),
.A2(n_672),
.B(n_690),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_775),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_899),
.B(n_876),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_874),
.B(n_733),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_919),
.B(n_751),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_918),
.A2(n_754),
.B(n_702),
.C(n_671),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_774),
.B(n_724),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_788),
.B(n_726),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_918),
.A2(n_754),
.B(n_661),
.C(n_762),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_830),
.A2(n_771),
.B(n_766),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_819),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_875),
.A2(n_753),
.B(n_740),
.C(n_737),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_875),
.A2(n_734),
.B1(n_423),
.B2(n_418),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_826),
.B(n_419),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_826),
.B(n_419),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_843),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_814),
.Y(n_990)
);

INVx6_ASAP7_75t_L g991 ( 
.A(n_821),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_892),
.A2(n_266),
.B1(n_227),
.B2(n_303),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_919),
.B(n_254),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_L g994 ( 
.A(n_913),
.B(n_88),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_913),
.B(n_423),
.Y(n_995)
);

AO32x1_ASAP7_75t_L g996 ( 
.A1(n_880),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_776),
.B(n_246),
.Y(n_997)
);

OR2x6_ASAP7_75t_SL g998 ( 
.A(n_864),
.B(n_183),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_827),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_821),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_776),
.B(n_247),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_SL g1002 ( 
.A(n_939),
.B(n_227),
.C(n_266),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_847),
.A2(n_423),
.B1(n_418),
.B2(n_251),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_874),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_832),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_840),
.B(n_423),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_892),
.B(n_418),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_914),
.B(n_292),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_790),
.A2(n_395),
.B(n_423),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_914),
.B(n_294),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_792),
.A2(n_395),
.B(n_423),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_905),
.B(n_84),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_SL g1013 ( 
.A1(n_947),
.A2(n_78),
.B(n_147),
.C(n_143),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_799),
.A2(n_395),
.B(n_423),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_847),
.A2(n_787),
.B(n_898),
.C(n_816),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_829),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_798),
.B(n_423),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_862),
.B(n_423),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_810),
.A2(n_302),
.B(n_294),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_904),
.A2(n_925),
.B1(n_820),
.B2(n_849),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_843),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_785),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_899),
.B(n_418),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_902),
.B(n_418),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_800),
.A2(n_418),
.B(n_110),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_779),
.A2(n_418),
.B(n_108),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_777),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_874),
.B(n_418),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_803),
.B(n_418),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_925),
.B(n_906),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_803),
.B(n_302),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_921),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_791),
.B(n_11),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_785),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_782),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_791),
.B(n_15),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_921),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_897),
.B(n_15),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_784),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_901),
.B(n_19),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_780),
.A2(n_141),
.B(n_134),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_837),
.B(n_122),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_907),
.B(n_24),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_943),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_841),
.B(n_25),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_870),
.Y(n_1046)
);

AO21x1_ASAP7_75t_L g1047 ( 
.A1(n_786),
.A2(n_26),
.B(n_28),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_933),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_906),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_904),
.A2(n_920),
.B1(n_937),
.B2(n_797),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_785),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_890),
.A2(n_29),
.B(n_31),
.C(n_35),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_797),
.B(n_115),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_834),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_845),
.B(n_29),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_805),
.A2(n_114),
.B(n_99),
.C(n_97),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_835),
.B(n_31),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_851),
.B(n_36),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_890),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_811),
.A2(n_85),
.B(n_92),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_795),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_853),
.A2(n_956),
.B1(n_927),
.B2(n_945),
.C(n_884),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_822),
.A2(n_48),
.B(n_90),
.C(n_94),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_886),
.A2(n_888),
.B1(n_837),
.B2(n_804),
.Y(n_1064)
);

CKINVDCx8_ASAP7_75t_R g1065 ( 
.A(n_846),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_836),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_L g1067 ( 
.A1(n_878),
.A2(n_917),
.B(n_807),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_934),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_891),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_851),
.B(n_859),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_785),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_900),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_881),
.A2(n_778),
.B(n_903),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_905),
.A2(n_884),
.B1(n_882),
.B2(n_885),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_889),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_812),
.B(n_861),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_891),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_944),
.B(n_941),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_848),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_957),
.A2(n_922),
.B(n_813),
.Y(n_1080)
);

AO21x1_ASAP7_75t_L g1081 ( 
.A1(n_809),
.A2(n_831),
.B(n_932),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_857),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_911),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_895),
.A2(n_824),
.B(n_808),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_812),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_802),
.A2(n_877),
.B(n_825),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_960),
.B(n_838),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_806),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_859),
.B(n_935),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_828),
.A2(n_935),
.B1(n_818),
.B2(n_926),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_931),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_839),
.B(n_929),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_860),
.B(n_952),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_926),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_948),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_941),
.B(n_924),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_812),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_812),
.A2(n_861),
.B1(n_789),
.B2(n_958),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_950),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_867),
.B(n_872),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_879),
.A2(n_896),
.B(n_946),
.C(n_949),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_833),
.B(n_861),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_940),
.Y(n_1103)
);

INVx8_ASAP7_75t_L g1104 ( 
.A(n_861),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_793),
.A2(n_801),
.B(n_809),
.C(n_831),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_854),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_930),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1062),
.A2(n_887),
.B(n_852),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_976),
.B(n_854),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_979),
.A2(n_817),
.B(n_815),
.C(n_955),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1064),
.A2(n_823),
.B(n_868),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1092),
.A2(n_958),
.B1(n_928),
.B2(n_893),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_968),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1077),
.B(n_842),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_968),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_973),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_975),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1064),
.A2(n_794),
.B(n_863),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1054),
.B(n_850),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1015),
.A2(n_823),
.B(n_868),
.C(n_866),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1080),
.A2(n_954),
.B(n_910),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1084),
.A2(n_909),
.B(n_908),
.Y(n_1122)
);

AO21x1_ASAP7_75t_L g1123 ( 
.A1(n_1020),
.A2(n_866),
.B(n_858),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_990),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_1020),
.A2(n_858),
.B(n_930),
.Y(n_1125)
);

AO32x2_ASAP7_75t_L g1126 ( 
.A1(n_1074),
.A2(n_928),
.A3(n_912),
.B1(n_873),
.B2(n_942),
.Y(n_1126)
);

AOI31xp67_ASAP7_75t_L g1127 ( 
.A1(n_1106),
.A2(n_923),
.A3(n_856),
.B(n_869),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_L g1128 ( 
.A(n_1087),
.B(n_938),
.C(n_936),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1105),
.A2(n_959),
.B(n_915),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_974),
.A2(n_855),
.B(n_916),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_962),
.A2(n_951),
.B(n_953),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_970),
.A2(n_972),
.B(n_982),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_984),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1086),
.A2(n_1014),
.B(n_983),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_964),
.A2(n_1101),
.B(n_1007),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1081),
.A2(n_966),
.B(n_1107),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_971),
.A2(n_1100),
.B1(n_1030),
.B2(n_1049),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_978),
.A2(n_1032),
.B1(n_1044),
.B2(n_1057),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1067),
.A2(n_1011),
.B(n_1009),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1074),
.A2(n_1078),
.B1(n_1050),
.B2(n_993),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1065),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1021),
.B(n_967),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1088),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1094),
.B(n_1008),
.Y(n_1144)
);

O2A1O1Ixp5_ASAP7_75t_L g1145 ( 
.A1(n_1050),
.A2(n_1047),
.B(n_1073),
.C(n_1098),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1007),
.A2(n_966),
.B(n_1023),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_999),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1066),
.B(n_1079),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_980),
.A2(n_969),
.B(n_981),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_969),
.A2(n_985),
.B(n_963),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1032),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1052),
.A2(n_1059),
.B1(n_992),
.B2(n_1061),
.C(n_1039),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_968),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_965),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1090),
.A2(n_1026),
.A3(n_1025),
.B(n_1098),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1005),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_997),
.A2(n_1001),
.B(n_1063),
.C(n_1082),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_989),
.B(n_1037),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_961),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1016),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1053),
.A2(n_1010),
.B1(n_1069),
.B2(n_1090),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1018),
.A2(n_1093),
.B(n_1096),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1024),
.A2(n_1041),
.B(n_1006),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_986),
.A2(n_1060),
.B(n_1058),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1027),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_992),
.A2(n_1002),
.B1(n_1019),
.B2(n_1013),
.C(n_1040),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1095),
.A2(n_1096),
.B1(n_1012),
.B2(n_977),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1012),
.B(n_1104),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1093),
.A2(n_1089),
.B(n_1070),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1004),
.B(n_1085),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1029),
.A2(n_1042),
.B(n_1017),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1089),
.A2(n_1103),
.B(n_1042),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1004),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1029),
.A2(n_987),
.B(n_988),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1035),
.Y(n_1175)
);

OAI22x1_ASAP7_75t_L g1176 ( 
.A1(n_1038),
.A2(n_1043),
.B1(n_1046),
.B2(n_1102),
.Y(n_1176)
);

BUFx4f_ASAP7_75t_SL g1177 ( 
.A(n_1000),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1099),
.B(n_1091),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1056),
.A2(n_1104),
.B(n_1033),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1036),
.A2(n_977),
.B(n_1031),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1048),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1104),
.A2(n_1028),
.B(n_994),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_987),
.A2(n_995),
.B(n_1034),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1072),
.Y(n_1184)
);

AO32x2_ASAP7_75t_L g1185 ( 
.A1(n_996),
.A2(n_977),
.A3(n_1019),
.B1(n_1045),
.B2(n_1055),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1028),
.A2(n_1031),
.B(n_1083),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1028),
.A2(n_1034),
.B(n_1022),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1022),
.A2(n_1097),
.B(n_1071),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1051),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1051),
.A2(n_1097),
.B(n_1071),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1075),
.Y(n_1191)
);

NAND3x1_ASAP7_75t_L g1192 ( 
.A(n_991),
.B(n_998),
.C(n_1068),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_1003),
.A2(n_996),
.B(n_1076),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_996),
.A2(n_1051),
.B(n_1071),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1004),
.B(n_1085),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1085),
.B(n_1097),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_991),
.A2(n_865),
.B(n_608),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1064),
.A2(n_725),
.B(n_773),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_SL g1199 ( 
.A1(n_962),
.A2(n_773),
.B(n_788),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_967),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_979),
.A2(n_608),
.B1(n_865),
.B2(n_774),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_976),
.B(n_774),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_973),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_967),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1015),
.A2(n_865),
.B(n_608),
.C(n_871),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1064),
.A2(n_865),
.B(n_608),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_976),
.B(n_774),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_979),
.A2(n_608),
.B1(n_865),
.B2(n_774),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1015),
.A2(n_865),
.B(n_608),
.C(n_871),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1084),
.A2(n_865),
.B(n_773),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1069),
.B(n_905),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_976),
.B(n_774),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_973),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_979),
.A2(n_608),
.B1(n_865),
.B2(n_774),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1065),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_968),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1065),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_968),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1064),
.A2(n_725),
.B(n_773),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_SL g1223 ( 
.A(n_1065),
.B(n_686),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_973),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1092),
.A2(n_608),
.B1(n_865),
.B2(n_883),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1084),
.A2(n_865),
.B(n_773),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1084),
.A2(n_865),
.B(n_773),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1064),
.A2(n_725),
.B(n_773),
.Y(n_1230)
);

OAI21xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1100),
.A2(n_865),
.B(n_608),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_967),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_967),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_976),
.B(n_865),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1064),
.A2(n_725),
.B(n_773),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_990),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_967),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1100),
.A2(n_608),
.B1(n_865),
.B2(n_871),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_976),
.B(n_665),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_979),
.A2(n_608),
.B1(n_865),
.B2(n_774),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_1104),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1084),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_973),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1081),
.A2(n_1106),
.A3(n_1020),
.B(n_1064),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1015),
.A2(n_608),
.B(n_865),
.C(n_883),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_976),
.B(n_665),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1243),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1116),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1133),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1240),
.A2(n_1225),
.B1(n_1217),
.B2(n_1201),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_1220),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1224),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1141),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1117),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1197),
.A2(n_1231),
.B1(n_1210),
.B2(n_1242),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1207),
.A2(n_1211),
.B1(n_1167),
.B2(n_1137),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1147),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1201),
.A2(n_1217),
.B1(n_1242),
.B2(n_1210),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1108),
.A2(n_1236),
.B1(n_1241),
.B2(n_1248),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1156),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1204),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1206),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1247),
.A2(n_1209),
.B1(n_1203),
.B2(n_1215),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1203),
.A2(n_1215),
.B1(n_1209),
.B2(n_1208),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1234),
.Y(n_1267)
);

BUFx4f_ASAP7_75t_L g1268 ( 
.A(n_1221),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1197),
.A2(n_1208),
.B1(n_1168),
.B2(n_1132),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1216),
.Y(n_1270)
);

BUFx8_ASAP7_75t_L g1271 ( 
.A(n_1235),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1166),
.A2(n_1150),
.B1(n_1132),
.B2(n_1140),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1239),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1243),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1218),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1154),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1144),
.B(n_1114),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1245),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1243),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1166),
.A2(n_1150),
.B1(n_1138),
.B2(n_1161),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1148),
.A2(n_1176),
.B1(n_1109),
.B2(n_1135),
.Y(n_1282)
);

BUFx8_ASAP7_75t_L g1283 ( 
.A(n_1159),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1151),
.B(n_1200),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1243),
.B(n_1223),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1124),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1160),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1168),
.A2(n_1112),
.B1(n_1109),
.B2(n_1165),
.Y(n_1288)
);

OAI21xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1119),
.A2(n_1178),
.B(n_1175),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1238),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1221),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1195),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1178),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1136),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1135),
.A2(n_1180),
.B1(n_1125),
.B2(n_1123),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1143),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1162),
.B1(n_1184),
.B2(n_1128),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1196),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1162),
.A2(n_1136),
.B1(n_1193),
.B2(n_1146),
.Y(n_1299)
);

NAND2x1p5_ASAP7_75t_L g1300 ( 
.A(n_1183),
.B(n_1213),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1221),
.Y(n_1301)
);

CKINVDCx6p67_ASAP7_75t_R g1302 ( 
.A(n_1181),
.Y(n_1302)
);

CKINVDCx11_ASAP7_75t_R g1303 ( 
.A(n_1177),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1157),
.A2(n_1158),
.B1(n_1142),
.B2(n_1213),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1182),
.A2(n_1186),
.B1(n_1119),
.B2(n_1169),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1193),
.A2(n_1146),
.B1(n_1164),
.B2(n_1172),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1191),
.A2(n_1152),
.B1(n_1164),
.B2(n_1192),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1198),
.A2(n_1222),
.B1(n_1230),
.B2(n_1237),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1196),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1170),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1212),
.A2(n_1226),
.B1(n_1227),
.B2(n_1131),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1191),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1189),
.Y(n_1313)
);

NAND2x1p5_ASAP7_75t_L g1314 ( 
.A(n_1113),
.B(n_1173),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1179),
.A2(n_1120),
.B1(n_1212),
.B2(n_1226),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1227),
.A2(n_1131),
.B1(n_1152),
.B2(n_1111),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1190),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1170),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1199),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1113),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1115),
.Y(n_1321)
);

CKINVDCx14_ASAP7_75t_R g1322 ( 
.A(n_1115),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1153),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1111),
.A2(n_1129),
.B1(n_1118),
.B2(n_1122),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_1173),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1187),
.A2(n_1219),
.B1(n_1188),
.B2(n_1129),
.Y(n_1326)
);

BUFx8_ASAP7_75t_L g1327 ( 
.A(n_1126),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1219),
.A2(n_1122),
.B1(n_1163),
.B2(n_1130),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1126),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1163),
.A2(n_1194),
.B1(n_1171),
.B2(n_1130),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1194),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1145),
.A2(n_1246),
.B1(n_1126),
.B2(n_1155),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1246),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1246),
.A2(n_1155),
.B1(n_1110),
.B2(n_1185),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1127),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1174),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1139),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_1134),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1202),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1205),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1214),
.B(n_1229),
.Y(n_1341)
);

INVx4_ASAP7_75t_SL g1342 ( 
.A(n_1185),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1185),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1121),
.A2(n_1228),
.B1(n_1232),
.B2(n_1233),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1244),
.A2(n_1240),
.B1(n_608),
.B2(n_1225),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1197),
.A2(n_608),
.B1(n_865),
.B2(n_871),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1225),
.B(n_608),
.Y(n_1347)
);

CKINVDCx16_ASAP7_75t_R g1348 ( 
.A(n_1124),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1240),
.A2(n_865),
.B1(n_608),
.B2(n_1225),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1220),
.Y(n_1350)
);

BUFx4f_ASAP7_75t_SL g1351 ( 
.A(n_1191),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1116),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1240),
.A2(n_865),
.B1(n_608),
.B2(n_1225),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1220),
.Y(n_1354)
);

OAI21xp33_ASAP7_75t_L g1355 ( 
.A1(n_1240),
.A2(n_608),
.B(n_865),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1220),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1220),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1206),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1225),
.A2(n_608),
.B1(n_865),
.B2(n_1201),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1240),
.A2(n_865),
.B1(n_608),
.B2(n_1225),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1197),
.A2(n_608),
.B1(n_865),
.B2(n_871),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1243),
.B(n_785),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1197),
.A2(n_608),
.B1(n_865),
.B2(n_871),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1220),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1225),
.B(n_608),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1243),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1116),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1240),
.A2(n_608),
.B1(n_1225),
.B2(n_865),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1240),
.A2(n_865),
.B1(n_608),
.B2(n_1225),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1220),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1243),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1116),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1294),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1294),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1333),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1309),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1328),
.A2(n_1344),
.B(n_1341),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1342),
.B(n_1260),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1337),
.Y(n_1379)
);

BUFx4f_ASAP7_75t_SL g1380 ( 
.A(n_1370),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1344),
.A2(n_1315),
.B(n_1308),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1368),
.A2(n_1347),
.B1(n_1365),
.B2(n_1258),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1262),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1335),
.A2(n_1288),
.B(n_1305),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1345),
.A2(n_1340),
.B(n_1339),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1288),
.A2(n_1332),
.B(n_1359),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1338),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1283),
.Y(n_1388)
);

BUFx2_ASAP7_75t_SL g1389 ( 
.A(n_1310),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1330),
.A2(n_1311),
.B(n_1340),
.Y(n_1390)
);

NOR2x1_ASAP7_75t_L g1391 ( 
.A(n_1281),
.B(n_1265),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1253),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1338),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1262),
.B(n_1278),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1260),
.B(n_1295),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1327),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1329),
.B(n_1326),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1331),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1330),
.A2(n_1311),
.B(n_1324),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1342),
.B(n_1257),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1334),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1300),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1346),
.A2(n_1363),
.B(n_1361),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1342),
.B(n_1295),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1300),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1327),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1252),
.B(n_1272),
.Y(n_1407)
);

AND2x6_ASAP7_75t_L g1408 ( 
.A(n_1274),
.B(n_1371),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1256),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1289),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1336),
.B(n_1297),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1355),
.B(n_1349),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1259),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1292),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1263),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1270),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1313),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1284),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1343),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1324),
.A2(n_1297),
.B(n_1306),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1304),
.A2(n_1317),
.B1(n_1360),
.B2(n_1353),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1317),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1282),
.B(n_1299),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1317),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1310),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1252),
.B(n_1272),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_SL g1427 ( 
.A1(n_1280),
.A2(n_1282),
.B(n_1352),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1349),
.B(n_1353),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1250),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1251),
.A2(n_1372),
.B(n_1254),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1298),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1293),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1367),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1318),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1360),
.A2(n_1369),
.B1(n_1359),
.B2(n_1269),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1369),
.B(n_1261),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1299),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1306),
.A2(n_1316),
.B(n_1280),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1266),
.A2(n_1321),
.B(n_1320),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1266),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1316),
.B(n_1307),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1319),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1318),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1264),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1314),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1362),
.A2(n_1285),
.B(n_1291),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1362),
.A2(n_1285),
.B(n_1291),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1277),
.A2(n_1249),
.B(n_1366),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1325),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_L g1451 ( 
.A(n_1296),
.B(n_1312),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1279),
.A2(n_1366),
.B(n_1371),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1323),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1267),
.A2(n_1358),
.B1(n_1273),
.B2(n_1271),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1382),
.B(n_1287),
.Y(n_1455)
);

AOI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1403),
.A2(n_1436),
.B(n_1412),
.C(n_1441),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1418),
.B(n_1348),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1434),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1396),
.B(n_1400),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1435),
.A2(n_1322),
.B1(n_1286),
.B2(n_1351),
.Y(n_1460)
);

OAI211xp5_ASAP7_75t_L g1461 ( 
.A1(n_1421),
.A2(n_1354),
.B(n_1356),
.C(n_1303),
.Y(n_1461)
);

NAND4xp25_ASAP7_75t_SL g1462 ( 
.A(n_1441),
.B(n_1357),
.C(n_1350),
.D(n_1351),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1404),
.B(n_1325),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_SL g1464 ( 
.A1(n_1442),
.A2(n_1428),
.B(n_1395),
.C(n_1406),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1442),
.A2(n_1276),
.B1(n_1290),
.B2(n_1302),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1444),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1407),
.A2(n_1426),
.B(n_1395),
.C(n_1427),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1417),
.B(n_1413),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1381),
.A2(n_1301),
.B(n_1268),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1378),
.B(n_1276),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1391),
.A2(n_1268),
.B(n_1290),
.Y(n_1471)
);

OAI211xp5_ASAP7_75t_L g1472 ( 
.A1(n_1391),
.A2(n_1283),
.B(n_1271),
.C(n_1364),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1410),
.A2(n_1255),
.B(n_1275),
.C(n_1407),
.Y(n_1473)
);

NOR2x1_ASAP7_75t_SL g1474 ( 
.A(n_1397),
.B(n_1389),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1410),
.B(n_1426),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1378),
.B(n_1400),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1409),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1437),
.B(n_1415),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1376),
.B(n_1431),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1454),
.A2(n_1397),
.B1(n_1422),
.B2(n_1424),
.C(n_1440),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1437),
.B(n_1415),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1438),
.A2(n_1420),
.B(n_1399),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1405),
.B(n_1402),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1394),
.B(n_1414),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1396),
.B(n_1414),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1397),
.A2(n_1422),
.B1(n_1424),
.B2(n_1406),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1377),
.A2(n_1390),
.B(n_1385),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1397),
.A2(n_1420),
.B(n_1399),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1419),
.B(n_1386),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1438),
.A2(n_1423),
.B(n_1411),
.C(n_1440),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1416),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1386),
.B(n_1394),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1385),
.A2(n_1390),
.B(n_1377),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1394),
.B(n_1432),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1397),
.B(n_1402),
.Y(n_1495)
);

OAI21xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1447),
.A2(n_1448),
.B(n_1446),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1386),
.B(n_1416),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1392),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1383),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1430),
.A2(n_1387),
.B(n_1393),
.Y(n_1500)
);

AOI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1427),
.A2(n_1401),
.B1(n_1423),
.B2(n_1411),
.C(n_1433),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1383),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1398),
.B(n_1429),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1380),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1405),
.B(n_1402),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1453),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1422),
.A2(n_1424),
.B(n_1450),
.C(n_1443),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_L g1509 ( 
.A(n_1445),
.B(n_1389),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1492),
.B(n_1384),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1492),
.B(n_1384),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1497),
.B(n_1398),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1483),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1499),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1458),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1507),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1455),
.A2(n_1411),
.B1(n_1388),
.B2(n_1402),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1482),
.B(n_1384),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1483),
.B(n_1379),
.Y(n_1520)
);

INVxp67_ASAP7_75t_SL g1521 ( 
.A(n_1500),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1478),
.B(n_1439),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1477),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1475),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1458),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1468),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1495),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1481),
.B(n_1439),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1489),
.B(n_1373),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1491),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1489),
.B(n_1374),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1502),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1488),
.B(n_1375),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1500),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1534),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1515),
.A2(n_1475),
.B(n_1464),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1534),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1534),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1522),
.B(n_1494),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1523),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1510),
.B(n_1476),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1521),
.A2(n_1487),
.B(n_1493),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1527),
.B(n_1506),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1513),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1476),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1527),
.B(n_1469),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1511),
.B(n_1493),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

INVx5_ASAP7_75t_L g1552 ( 
.A(n_1527),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1511),
.B(n_1490),
.Y(n_1553)
);

AOI31xp33_ASAP7_75t_L g1554 ( 
.A1(n_1518),
.A2(n_1456),
.A3(n_1473),
.B(n_1472),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1532),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1514),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1532),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1522),
.B(n_1484),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1514),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1513),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1514),
.Y(n_1561)
);

BUFx2_ASAP7_75t_SL g1562 ( 
.A(n_1516),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1479),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1529),
.B(n_1501),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1512),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1531),
.B(n_1504),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1563),
.B(n_1524),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1541),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1537),
.B(n_1515),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1555),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1563),
.B(n_1524),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1563),
.B(n_1531),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1555),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1557),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1557),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1565),
.A2(n_1455),
.B1(n_1527),
.B2(n_1480),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1535),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1566),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1566),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1513),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1513),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1498),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1545),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1513),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1543),
.B(n_1520),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1559),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1559),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1565),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1535),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1553),
.B(n_1545),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1537),
.B(n_1512),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1540),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1545),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1561),
.Y(n_1600)
);

OAI33xp33_ASAP7_75t_L g1601 ( 
.A1(n_1540),
.A2(n_1466),
.A3(n_1558),
.B1(n_1528),
.B2(n_1465),
.B3(n_1530),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1561),
.Y(n_1602)
);

NAND4xp25_ASAP7_75t_L g1603 ( 
.A(n_1536),
.B(n_1461),
.C(n_1467),
.D(n_1473),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1540),
.B(n_1526),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1558),
.B(n_1526),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1579),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1579),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1553),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_SL g1609 ( 
.A(n_1596),
.B(n_1562),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1596),
.B(n_1564),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1572),
.Y(n_1612)
);

NAND2x2_ASAP7_75t_L g1613 ( 
.A(n_1603),
.B(n_1388),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1580),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1599),
.B(n_1564),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1599),
.B(n_1564),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1552),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1550),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1585),
.B(n_1536),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_1593),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1601),
.A2(n_1554),
.B1(n_1550),
.B2(n_1519),
.C(n_1464),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1575),
.Y(n_1624)
);

NOR2x1_ASAP7_75t_R g1625 ( 
.A(n_1603),
.B(n_1505),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1576),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1568),
.B(n_1517),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1576),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1577),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1577),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1569),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1568),
.B(n_1517),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1550),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1580),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1580),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1569),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1581),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1590),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1601),
.B(n_1498),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1590),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1597),
.B(n_1558),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1592),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1588),
.B(n_1552),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1581),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1592),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1588),
.B(n_1545),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1573),
.B(n_1549),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1609),
.B(n_1589),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1611),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1618),
.B(n_1552),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1573),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1647),
.B(n_1571),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1627),
.B(n_1571),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1646),
.B(n_1589),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1612),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1612),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1591),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1606),
.B(n_1607),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1591),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1611),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1641),
.B(n_1605),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1631),
.B(n_1598),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1641),
.B(n_1636),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1643),
.B(n_1595),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1637),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1625),
.B(n_1505),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1639),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1620),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1615),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1644),
.B(n_1582),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1618),
.B(n_1643),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1643),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1644),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1622),
.B(n_1582),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1623),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1656),
.Y(n_1683)
);

O2A1O1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1670),
.A2(n_1611),
.B(n_1613),
.C(n_1578),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1670),
.A2(n_1679),
.B1(n_1671),
.B2(n_1613),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1671),
.B(n_1623),
.C(n_1626),
.Y(n_1686)
);

OAI321xp33_ASAP7_75t_L g1687 ( 
.A1(n_1679),
.A2(n_1460),
.A3(n_1471),
.B1(n_1633),
.B2(n_1519),
.C(n_1616),
.Y(n_1687)
);

XNOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1651),
.B(n_1457),
.Y(n_1688)
);

AOI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1660),
.A2(n_1629),
.B(n_1628),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1610),
.Y(n_1690)
);

OAI211xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1677),
.A2(n_1630),
.B(n_1642),
.C(n_1640),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1669),
.A2(n_1633),
.B(n_1548),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1678),
.A2(n_1673),
.B1(n_1668),
.B2(n_1653),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1657),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1658),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1665),
.A2(n_1551),
.B1(n_1645),
.B2(n_1640),
.C(n_1638),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1665),
.B(n_1642),
.C(n_1638),
.Y(n_1697)
);

OAI22xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1650),
.A2(n_1645),
.B1(n_1604),
.B2(n_1552),
.Y(n_1698)
);

AOI322xp5_ASAP7_75t_L g1699 ( 
.A1(n_1678),
.A2(n_1619),
.A3(n_1616),
.B1(n_1617),
.B2(n_1574),
.C1(n_1604),
.C2(n_1584),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1672),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_SL g1702 ( 
.A1(n_1649),
.A2(n_1560),
.B(n_1546),
.C(n_1574),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1661),
.Y(n_1703)
);

OAI33xp33_ASAP7_75t_L g1704 ( 
.A1(n_1661),
.A2(n_1635),
.A3(n_1634),
.B1(n_1614),
.B2(n_1602),
.B3(n_1600),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1619),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1663),
.A2(n_1634),
.B(n_1614),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1617),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1683),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1685),
.A2(n_1676),
.B1(n_1659),
.B2(n_1648),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1707),
.B(n_1676),
.Y(n_1710)
);

AOI21xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1684),
.A2(n_1650),
.B(n_1648),
.Y(n_1711)
);

AOI32xp33_ASAP7_75t_L g1712 ( 
.A1(n_1687),
.A2(n_1691),
.A3(n_1693),
.B1(n_1690),
.B2(n_1696),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1693),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1694),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1695),
.Y(n_1715)
);

OAI21xp33_ASAP7_75t_L g1716 ( 
.A1(n_1699),
.A2(n_1664),
.B(n_1652),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1687),
.A2(n_1675),
.B1(n_1659),
.B2(n_1681),
.C(n_1674),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1686),
.A2(n_1675),
.B(n_1655),
.C(n_1551),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1700),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1701),
.Y(n_1720)
);

OAI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1688),
.A2(n_1674),
.B(n_1682),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1703),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1697),
.A2(n_1551),
.B1(n_1552),
.B2(n_1462),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1689),
.A2(n_1635),
.B1(n_1662),
.B2(n_1654),
.C(n_1533),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1705),
.B(n_1587),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1698),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1692),
.A2(n_1548),
.B(n_1486),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1713),
.B(n_1712),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1710),
.B(n_1709),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1723),
.A2(n_1552),
.B1(n_1706),
.B2(n_1551),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1711),
.A2(n_1717),
.B1(n_1716),
.B2(n_1721),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1726),
.Y(n_1732)
);

NAND2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1708),
.B(n_1388),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1714),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1725),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1715),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1722),
.B(n_1702),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1731),
.A2(n_1718),
.B1(n_1727),
.B2(n_1724),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1728),
.B(n_1720),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1732),
.A2(n_1727),
.B(n_1551),
.C(n_1704),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1737),
.B(n_1552),
.Y(n_1742)
);

NOR2xp67_ASAP7_75t_L g1743 ( 
.A(n_1729),
.B(n_1600),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1733),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1733),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_L g1746 ( 
.A(n_1735),
.B(n_1738),
.C(n_1734),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_SL g1747 ( 
.A1(n_1730),
.A2(n_1450),
.B(n_1474),
.Y(n_1747)
);

NAND4xp25_ASAP7_75t_L g1748 ( 
.A(n_1740),
.B(n_1736),
.C(n_1485),
.D(n_1470),
.Y(n_1748)
);

AND4x1_ASAP7_75t_L g1749 ( 
.A(n_1746),
.B(n_1736),
.C(n_1509),
.D(n_1451),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1739),
.A2(n_1741),
.B1(n_1745),
.B2(n_1744),
.C(n_1747),
.Y(n_1750)
);

XOR2xp5_ASAP7_75t_L g1751 ( 
.A(n_1742),
.B(n_1545),
.Y(n_1751)
);

AOI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1743),
.A2(n_1508),
.B(n_1459),
.C(n_1496),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1750),
.A2(n_1602),
.B1(n_1521),
.B2(n_1594),
.C(n_1562),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1748),
.A2(n_1594),
.B1(n_1533),
.B2(n_1583),
.C(n_1584),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1752),
.A2(n_1470),
.B(n_1583),
.C(n_1533),
.Y(n_1755)
);

OAI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1751),
.A2(n_1560),
.B(n_1546),
.C(n_1594),
.Y(n_1756)
);

AOI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1749),
.A2(n_1546),
.B1(n_1560),
.B2(n_1544),
.C(n_1538),
.Y(n_1757)
);

OAI221xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1750),
.A2(n_1495),
.B1(n_1516),
.B2(n_1525),
.C(n_1463),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1758),
.B(n_1567),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1753),
.B(n_1549),
.Y(n_1760)
);

NAND4xp75_ASAP7_75t_L g1761 ( 
.A(n_1757),
.B(n_1516),
.C(n_1463),
.D(n_1469),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1756),
.B(n_1449),
.C(n_1503),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1755),
.Y(n_1763)
);

XNOR2xp5_ASAP7_75t_L g1764 ( 
.A(n_1763),
.B(n_1754),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1759),
.A2(n_1548),
.B1(n_1495),
.B2(n_1525),
.C(n_1535),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1760),
.A2(n_1544),
.B(n_1539),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1764),
.B(n_1762),
.Y(n_1767)
);

AO22x2_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1766),
.B1(n_1761),
.B2(n_1765),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1768),
.B(n_1544),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1770),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1769),
.Y(n_1772)
);

AOI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1535),
.B1(n_1539),
.B2(n_1538),
.C(n_1556),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1772),
.A2(n_1548),
.B1(n_1539),
.B2(n_1538),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1774),
.B(n_1544),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1773),
.B(n_1452),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1776),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_R g1778 ( 
.A1(n_1777),
.A2(n_1544),
.B1(n_1525),
.B2(n_1538),
.C(n_1539),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1408),
.B1(n_1425),
.B2(n_1556),
.Y(n_1779)
);


endmodule