module fake_jpeg_5815_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_19),
.B(n_9),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_35),
.B1(n_25),
.B2(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_30),
.C(n_33),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_59),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_22),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_26),
.B1(n_35),
.B2(n_34),
.Y(n_86)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_60),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_34),
.B1(n_22),
.B2(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_73),
.Y(n_100)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_80),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_30),
.Y(n_84)
);

NOR2x1_ASAP7_75t_R g107 ( 
.A(n_84),
.B(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_87),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_93),
.B1(n_19),
.B2(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_46),
.B1(n_41),
.B2(n_45),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_90),
.B1(n_67),
.B2(n_46),
.Y(n_108)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_91),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_46),
.B1(n_40),
.B2(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_44),
.B1(n_19),
.B2(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_119),
.B1(n_123),
.B2(n_36),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_50),
.C(n_60),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_88),
.C(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_111),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_68),
.B(n_37),
.C(n_40),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_59),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_118),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_46),
.B1(n_44),
.B2(n_67),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_122),
.B1(n_73),
.B2(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_45),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_20),
.B1(n_24),
.B2(n_45),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_44),
.B1(n_47),
.B2(n_37),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_47),
.B1(n_40),
.B2(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_47),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_130),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_116),
.B1(n_112),
.B2(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_42),
.C(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_139),
.Y(n_183)
);

XOR2x2_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_39),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_147),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_44),
.B1(n_65),
.B2(n_70),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_48),
.B(n_28),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_153),
.B1(n_114),
.B2(n_113),
.Y(n_174)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_68),
.B(n_37),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_75),
.B1(n_81),
.B2(n_85),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_80),
.B1(n_98),
.B2(n_96),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_150),
.B1(n_157),
.B2(n_105),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_39),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_91),
.B1(n_40),
.B2(n_36),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_158),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_103),
.B(n_48),
.CI(n_42),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_61),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_116),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_40),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_42),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_163),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_154),
.B(n_48),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_185),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_117),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_167),
.C(n_173),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_128),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_175),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_65),
.B1(n_127),
.B2(n_124),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_65),
.B1(n_124),
.B2(n_83),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_140),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_20),
.B1(n_32),
.B2(n_113),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_31),
.B1(n_114),
.B2(n_28),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_136),
.B1(n_149),
.B2(n_131),
.Y(n_199)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_42),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_182),
.B(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_61),
.C(n_42),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_181),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_31),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_48),
.C(n_78),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_17),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_21),
.B(n_28),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_135),
.B1(n_142),
.B2(n_156),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_189),
.B1(n_147),
.B2(n_129),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_17),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_154),
.A3(n_141),
.B1(n_133),
.B2(n_132),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_197),
.B(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_211),
.B1(n_171),
.B2(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_160),
.B(n_132),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_178),
.CI(n_186),
.CON(n_226),
.SN(n_226)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_204),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_21),
.B(n_17),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_161),
.A2(n_28),
.B1(n_120),
.B2(n_17),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_212),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_21),
.B(n_1),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_169),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_0),
.B(n_1),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_11),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_163),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_241),
.CI(n_197),
.CON(n_250),
.SN(n_250)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_167),
.C(n_166),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_240),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_173),
.C(n_184),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_246),
.B1(n_247),
.B2(n_199),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_190),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_174),
.B1(n_159),
.B2(n_190),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_242),
.B1(n_211),
.B2(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_182),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_172),
.B1(n_175),
.B2(n_120),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_78),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_102),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_226),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_256),
.B1(n_264),
.B2(n_242),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_198),
.B(n_194),
.C(n_201),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_255),
.A2(n_260),
.B1(n_265),
.B2(n_245),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_195),
.B1(n_201),
.B2(n_219),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_248),
.B(n_236),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_220),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_259),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_203),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_193),
.B1(n_217),
.B2(n_210),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_261),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_233),
.A2(n_195),
.B1(n_193),
.B2(n_214),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_216),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_268),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_221),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_269),
.C(n_262),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_207),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_207),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_11),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_278),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_241),
.C(n_228),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_279),
.C(n_283),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_239),
.C(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_229),
.C(n_225),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_247),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_267),
.B(n_246),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_251),
.A2(n_257),
.B1(n_249),
.B2(n_270),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_222),
.B1(n_212),
.B2(n_253),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_248),
.B1(n_269),
.B2(n_238),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_289),
.B(n_293),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_250),
.B(n_226),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_279),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_12),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_213),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_300),
.C(n_302),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_276),
.B(n_282),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_276),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_213),
.C(n_2),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_12),
.B1(n_15),
.B2(n_9),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_289),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_271),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_308),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_315),
.B1(n_14),
.B2(n_16),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_6),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_312),
.C(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_12),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_11),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_320),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_319),
.B(n_9),
.C(n_10),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_290),
.CI(n_295),
.CON(n_320),
.SN(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_290),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_323),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_6),
.C(n_7),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_306),
.B1(n_311),
.B2(n_310),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_320),
.B(n_316),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_307),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_330),
.B(n_319),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_327),
.A2(n_329),
.B(n_323),
.Y(n_332)
);

AOI221xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.C(n_16),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_13),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_328),
.C(n_334),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.C(n_331),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_327),
.C(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_10),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_13),
.B(n_7),
.Y(n_340)
);


endmodule