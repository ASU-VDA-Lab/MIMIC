module fake_jpeg_757_n_494 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_7),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_49),
.Y(n_113)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_51),
.B(n_52),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_7),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_53),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_61),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_68),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_72),
.B(n_96),
.Y(n_154)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_87),
.B(n_93),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_14),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_100),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_15),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_20),
.B1(n_15),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_103),
.A2(n_116),
.B1(n_124),
.B2(n_136),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_110),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_41),
.B1(n_46),
.B2(n_15),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_46),
.B1(n_41),
.B2(n_43),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_162),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_47),
.B1(n_48),
.B2(n_45),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_47),
.B1(n_45),
.B2(n_34),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_126),
.A2(n_139),
.B1(n_16),
.B2(n_2),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_32),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_146),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_76),
.A2(n_23),
.B1(n_36),
.B2(n_43),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_54),
.A2(n_43),
.B1(n_32),
.B2(n_23),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_82),
.A2(n_29),
.B1(n_19),
.B2(n_34),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_67),
.B1(n_63),
.B2(n_62),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_31),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_58),
.B(n_31),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_151),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_65),
.B(n_19),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_56),
.A2(n_29),
.B1(n_39),
.B2(n_42),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_79),
.B1(n_75),
.B2(n_71),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_97),
.A2(n_42),
.B1(n_39),
.B2(n_24),
.Y(n_162)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_82),
.B1(n_77),
.B2(n_87),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_24),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_172),
.B(n_178),
.Y(n_257)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_176),
.A2(n_181),
.B1(n_196),
.B2(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_22),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_22),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_188),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_90),
.B1(n_101),
.B2(n_100),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_182),
.A2(n_190),
.B1(n_208),
.B2(n_215),
.Y(n_225)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_1),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_204),
.A3(n_117),
.B1(n_104),
.B2(n_4),
.Y(n_226)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_133),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_115),
.B(n_69),
.C(n_68),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_192),
.C(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_118),
.B(n_61),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_110),
.A2(n_16),
.B(n_9),
.C(n_14),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_193),
.A2(n_217),
.B(n_218),
.Y(n_246)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_198),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_113),
.A2(n_57),
.B1(n_16),
.B2(n_9),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_1),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_126),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_105),
.B1(n_130),
.B2(n_121),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_203),
.A2(n_214),
.B1(n_187),
.B2(n_193),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_1),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_141),
.A2(n_16),
.B(n_10),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_105),
.B(n_108),
.Y(n_239)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_207),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_124),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_103),
.A2(n_116),
.B1(n_136),
.B2(n_114),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_114),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_104),
.B1(n_106),
.B2(n_113),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_133),
.B(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_164),
.B1(n_155),
.B2(n_106),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_219),
.A2(n_221),
.B1(n_230),
.B2(n_242),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_237),
.B1(n_249),
.B2(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_192),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_157),
.B1(n_127),
.B2(n_130),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_144),
.B1(n_149),
.B2(n_166),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_212),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_175),
.A2(n_144),
.B1(n_121),
.B2(n_108),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_149),
.B1(n_165),
.B2(n_129),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_215),
.B1(n_180),
.B2(n_202),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_132),
.B(n_112),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_217),
.B(n_200),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_175),
.A2(n_122),
.B1(n_165),
.B2(n_4),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_255),
.A2(n_186),
.B1(n_216),
.B2(n_172),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_265),
.B1(n_268),
.B2(n_275),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_178),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_229),
.C(n_244),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_186),
.B(n_188),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_261),
.A2(n_281),
.B(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_249),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_263),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_269),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_246),
.B1(n_186),
.B2(n_247),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_176),
.B1(n_199),
.B2(n_183),
.Y(n_266)
);

BUFx4f_ASAP7_75t_SL g301 ( 
.A(n_266),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_225),
.A2(n_192),
.B1(n_204),
.B2(n_169),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_224),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_277),
.C(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_184),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_273),
.B(n_242),
.Y(n_307)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_213),
.B1(n_200),
.B2(n_218),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_224),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_241),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_237),
.B(n_257),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_217),
.B(n_185),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_284),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_241),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_228),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_223),
.Y(n_287)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_303),
.C(n_314),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_236),
.B1(n_226),
.B2(n_250),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_308),
.B1(n_280),
.B2(n_265),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_302),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_258),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_263),
.A2(n_219),
.B1(n_220),
.B2(n_232),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_259),
.A2(n_232),
.B1(n_256),
.B2(n_251),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_279),
.B1(n_274),
.B2(n_262),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_288),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_177),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_280),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_317),
.A2(n_327),
.B1(n_333),
.B2(n_340),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_263),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_328),
.C(n_341),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_306),
.A2(n_263),
.B1(n_281),
.B2(n_259),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_331),
.B1(n_335),
.B2(n_336),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_282),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_324),
.B(n_293),
.Y(n_366)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_300),
.Y(n_326)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_298),
.A2(n_281),
.B1(n_268),
.B2(n_282),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_272),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_332),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_268),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_282),
.B1(n_275),
.B2(n_261),
.Y(n_333)
);

NAND3xp33_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_179),
.C(n_275),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_297),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_306),
.A2(n_261),
.B1(n_284),
.B2(n_279),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_291),
.A2(n_279),
.B1(n_284),
.B2(n_266),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_310),
.A2(n_267),
.B1(n_283),
.B2(n_278),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_337),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_277),
.B(n_271),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_339),
.A2(n_324),
.B(n_323),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_287),
.B1(n_269),
.B2(n_256),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_228),
.C(n_189),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_302),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_351),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_345),
.B(n_362),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_310),
.B1(n_296),
.B2(n_301),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_347),
.A2(n_349),
.B1(n_337),
.B2(n_338),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_320),
.A2(n_310),
.B1(n_296),
.B2(n_301),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_313),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_325),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_355),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_289),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_351),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_339),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_289),
.C(n_290),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_359),
.C(n_363),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_290),
.C(n_304),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_330),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_360),
.A2(n_321),
.B1(n_294),
.B2(n_301),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_326),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_295),
.C(n_309),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_323),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_364),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_365),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_366),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_305),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_329),
.C(n_336),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_373),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_363),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_385),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_343),
.B(n_317),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_382),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_327),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_386),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_316),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_378),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_353),
.A2(n_346),
.B(n_368),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_379),
.A2(n_299),
.B1(n_287),
.B2(n_223),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_350),
.B(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_384),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_342),
.A2(n_367),
.B1(n_361),
.B2(n_356),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_322),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_332),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_390),
.Y(n_413)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_338),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_344),
.B(n_324),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_393),
.Y(n_414)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_394),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_397),
.A2(n_412),
.B1(n_372),
.B2(n_371),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_391),
.A2(n_367),
.B(n_342),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_403),
.A2(n_406),
.B(n_409),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_365),
.C(n_321),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_408),
.C(n_369),
.Y(n_416)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_405),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_301),
.B(n_299),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_392),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_252),
.C(n_235),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_388),
.A2(n_252),
.B(n_235),
.Y(n_409)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_380),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_410),
.Y(n_424)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_411),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_378),
.A2(n_222),
.B1(n_245),
.B2(n_251),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_404),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_415),
.B(n_370),
.Y(n_418)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_425),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_376),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_428),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_403),
.A2(n_397),
.B(n_400),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_427),
.Y(n_443)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_382),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_386),
.C(n_374),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_433),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_393),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_222),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_431),
.A2(n_414),
.B1(n_399),
.B2(n_413),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_406),
.A2(n_372),
.B(n_387),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_432),
.A2(n_412),
.B(n_409),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_381),
.C(n_238),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_446),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_445),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_437),
.A2(n_428),
.B1(n_429),
.B2(n_431),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_425),
.A2(n_419),
.B1(n_432),
.B2(n_421),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_444),
.B1(n_448),
.B2(n_234),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_418),
.A2(n_414),
.B(n_413),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_238),
.B(n_168),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_417),
.A2(n_399),
.B1(n_381),
.B2(n_222),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_423),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_174),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_420),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_420),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_455),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_433),
.C(n_422),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_454),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_449),
.B(n_424),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_210),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_458),
.Y(n_468)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_457),
.A2(n_462),
.B(n_439),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_227),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_211),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_460),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_227),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_191),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_463),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_197),
.Y(n_463)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_450),
.A2(n_441),
.B(n_452),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_467),
.A2(n_470),
.B(n_471),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_439),
.B(n_437),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g471 ( 
.A1(n_453),
.A2(n_446),
.B(n_194),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_234),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_473),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_212),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_466),
.A2(n_173),
.B(n_212),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_476),
.A2(n_465),
.B(n_474),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_167),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_481),
.B(n_474),
.Y(n_484)
);

OAI31xp33_ASAP7_75t_SL g479 ( 
.A1(n_469),
.A2(n_207),
.A3(n_170),
.B(n_209),
.Y(n_479)
);

O2A1O1Ixp33_ASAP7_75t_SL g486 ( 
.A1(n_479),
.A2(n_209),
.B(n_3),
.C(n_5),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_209),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_483),
.Y(n_489)
);

O2A1O1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_484),
.A2(n_486),
.B(n_2),
.C(n_3),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_485),
.A2(n_480),
.B(n_479),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_487),
.A2(n_2),
.B(n_3),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_488),
.B(n_5),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_490),
.B(n_491),
.C(n_489),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_492),
.A2(n_5),
.B(n_6),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_5),
.Y(n_494)
);


endmodule