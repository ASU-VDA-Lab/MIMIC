module fake_jpeg_21096_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_70),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_57),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_64),
.CI(n_46),
.CON(n_98),
.SN(n_98)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_60),
.B1(n_47),
.B2(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_89),
.B1(n_71),
.B2(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_47),
.B1(n_51),
.B2(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_98),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_88),
.B(n_89),
.C(n_83),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_0),
.B(n_1),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_67),
.B1(n_68),
.B2(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_54),
.B1(n_48),
.B2(n_44),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_64),
.B1(n_46),
.B2(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_59),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_66),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_0),
.Y(n_126)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_63),
.B1(n_53),
.B2(n_55),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_8),
.Y(n_131)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_12),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_132),
.B(n_130),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_105),
.C(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_135),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_115),
.B(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_132),
.B(n_134),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_137),
.B(n_139),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_138),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_128),
.B(n_125),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_124),
.B1(n_122),
.B2(n_109),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_107),
.A3(n_118),
.B1(n_113),
.B2(n_16),
.C1(n_17),
.C2(n_22),
.Y(n_147)
);

AOI332xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_118),
.A3(n_14),
.B1(n_15),
.B2(n_23),
.B3(n_24),
.C1(n_25),
.C2(n_26),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_113),
.Y(n_149)
);

AOI321xp33_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_13),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.C(n_39),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_40),
.Y(n_151)
);


endmodule