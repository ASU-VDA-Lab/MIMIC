module fake_jpeg_24432_n_18 (n_3, n_2, n_1, n_0, n_4, n_5, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_18;

wire n_13;
wire n_11;
wire n_14;
wire n_17;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_8),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_12),
.B(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_10),
.B(n_14),
.Y(n_16)
);

AO221x1_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_1),
.C(n_2),
.Y(n_18)
);


endmodule