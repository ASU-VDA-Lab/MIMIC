module fake_netlist_5_2406_n_4251 (n_924, n_1263, n_977, n_611, n_1126, n_1166, n_469, n_82, n_785, n_549, n_532, n_1161, n_1150, n_226, n_667, n_790, n_1055, n_111, n_880, n_544, n_1007, n_155, n_552, n_1292, n_1198, n_1360, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_1323, n_688, n_1353, n_800, n_1347, n_671, n_819, n_1022, n_915, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_292, n_625, n_854, n_674, n_417, n_516, n_933, n_1152, n_497, n_606, n_275, n_26, n_877, n_2, n_755, n_1118, n_6, n_947, n_1285, n_373, n_307, n_1359, n_530, n_87, n_150, n_1107, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_191, n_1104, n_1294, n_659, n_51, n_1257, n_171, n_1182, n_579, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_1314, n_709, n_317, n_1236, n_569, n_227, n_920, n_1289, n_94, n_335, n_370, n_976, n_343, n_308, n_297, n_156, n_1078, n_775, n_219, n_157, n_600, n_1328, n_223, n_264, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_436, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_1267, n_496, n_958, n_1034, n_670, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_395, n_164, n_553, n_901, n_813, n_1284, n_214, n_675, n_888, n_1167, n_637, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_468, n_213, n_129, n_342, n_464, n_363, n_197, n_1069, n_1075, n_1322, n_460, n_889, n_973, n_477, n_571, n_461, n_1211, n_1197, n_907, n_190, n_989, n_1039, n_34, n_228, n_283, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_440, n_793, n_478, n_476, n_534, n_884, n_345, n_944, n_91, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_1319, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_596, n_558, n_702, n_1276, n_822, n_728, n_266, n_1162, n_272, n_1199, n_352, n_53, n_1038, n_520, n_409, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_434, n_868, n_639, n_914, n_411, n_414, n_1293, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_64, n_759, n_28, n_806, n_324, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_706, n_746, n_747, n_52, n_784, n_110, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_776, n_367, n_452, n_525, n_1260, n_649, n_547, n_43, n_1191, n_116, n_284, n_1128, n_139, n_744, n_590, n_629, n_1308, n_254, n_1233, n_23, n_526, n_293, n_372, n_677, n_244, n_47, n_1333, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1008, n_946, n_1001, n_498, n_689, n_738, n_640, n_252, n_624, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1195, n_610, n_936, n_568, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1158, n_563, n_1145, n_878, n_524, n_204, n_394, n_1049, n_1153, n_741, n_1306, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_1362, n_456, n_959, n_535, n_152, n_940, n_9, n_592, n_1169, n_45, n_1017, n_123, n_978, n_1054, n_1269, n_1095, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_484, n_1033, n_442, n_131, n_636, n_660, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_374, n_185, n_396, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_723, n_1065, n_1336, n_473, n_1309, n_1043, n_355, n_486, n_614, n_337, n_88, n_1286, n_1177, n_1355, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_361, n_700, n_1237, n_573, n_69, n_1132, n_388, n_1300, n_1127, n_761, n_1006, n_329, n_274, n_1270, n_582, n_1332, n_73, n_19, n_309, n_30, n_512, n_84, n_130, n_322, n_1249, n_652, n_1111, n_25, n_1349, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_44, n_224, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_1304, n_1324, n_987, n_261, n_174, n_767, n_993, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_83, n_513, n_1094, n_1354, n_560, n_340, n_1351, n_1044, n_1205, n_346, n_1209, n_495, n_602, n_574, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_490, n_1327, n_996, n_921, n_233, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1037, n_1080, n_1274, n_1316, n_426, n_1082, n_589, n_716, n_562, n_62, n_952, n_1229, n_391, n_701, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_162, n_960, n_222, n_1290, n_1123, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1029, n_925, n_1206, n_424, n_1311, n_256, n_950, n_380, n_419, n_1346, n_444, n_1299, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_376, n_967, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_1357, n_483, n_683, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_983, n_38, n_280, n_1305, n_873, n_378, n_1112, n_762, n_1283, n_17, n_690, n_33, n_583, n_302, n_1343, n_1203, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1288, n_212, n_385, n_507, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1301, n_1363, n_1185, n_991, n_828, n_779, n_576, n_1143, n_1329, n_1312, n_804, n_537, n_945, n_492, n_153, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_883, n_470, n_325, n_449, n_132, n_1214, n_1342, n_900, n_856, n_918, n_942, n_189, n_1147, n_13, n_1077, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_831, n_964, n_1350, n_1096, n_234, n_833, n_5, n_225, n_1307, n_988, n_814, n_192, n_1201, n_1114, n_655, n_669, n_472, n_1176, n_387, n_1149, n_398, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_50, n_430, n_510, n_216, n_311, n_830, n_1296, n_801, n_241, n_875, n_357, n_1110, n_445, n_749, n_1134, n_1358, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_734, n_638, n_866, n_107, n_969, n_1019, n_1105, n_249, n_304, n_1338, n_577, n_338, n_149, n_693, n_14, n_836, n_990, n_975, n_1256, n_567, n_778, n_1122, n_151, n_306, n_458, n_770, n_1102, n_711, n_85, n_1187, n_1164, n_489, n_1174, n_617, n_1303, n_876, n_1190, n_118, n_601, n_917, n_966, n_253, n_1116, n_1212, n_172, n_206, n_217, n_726, n_982, n_818, n_861, n_1183, n_899, n_1253, n_210, n_774, n_1335, n_1059, n_1345, n_176, n_1133, n_557, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_393, n_108, n_487, n_665, n_66, n_177, n_421, n_1356, n_910, n_768, n_1302, n_205, n_1136, n_1313, n_754, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_1310, n_202, n_427, n_791, n_732, n_193, n_808, n_797, n_1025, n_500, n_1067, n_148, n_435, n_159, n_766, n_541, n_538, n_1117, n_799, n_687, n_715, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1297, n_1155, n_89, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_1352, n_626, n_1144, n_1137, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_194, n_855, n_1178, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_605, n_1273, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_1318, n_780, n_998, n_467, n_1227, n_840, n_1334, n_501, n_823, n_245, n_725, n_1295, n_672, n_581, n_382, n_554, n_898, n_1013, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_909, n_997, n_932, n_612, n_788, n_1326, n_119, n_1268, n_559, n_825, n_508, n_506, n_1320, n_737, n_986, n_509, n_1317, n_147, n_1281, n_67, n_1192, n_1024, n_1063, n_209, n_733, n_941, n_981, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1108, n_782, n_1100, n_862, n_760, n_381, n_220, n_390, n_1330, n_31, n_481, n_769, n_42, n_1046, n_271, n_934, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_1341, n_570, n_1361, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1225, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_221, n_622, n_1087, n_386, n_994, n_848, n_1223, n_1272, n_104, n_682, n_56, n_141, n_1247, n_922, n_816, n_591, n_145, n_1344, n_313, n_631, n_479, n_1246, n_1339, n_432, n_839, n_1210, n_328, n_140, n_1250, n_369, n_871, n_598, n_685, n_928, n_608, n_78, n_772, n_499, n_517, n_98, n_402, n_413, n_1086, n_796, n_236, n_1012, n_1, n_1348, n_903, n_740, n_203, n_384, n_80, n_35, n_1315, n_277, n_1061, n_92, n_333, n_1298, n_462, n_1193, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_40, n_1028, n_781, n_474, n_542, n_463, n_595, n_502, n_466, n_420, n_1337, n_632, n_699, n_979, n_1245, n_846, n_465, n_76, n_362, n_1321, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1103, n_648, n_312, n_1076, n_1091, n_494, n_641, n_730, n_1325, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1220, n_37, n_229, n_437, n_60, n_403, n_453, n_1130, n_720, n_0, n_863, n_805, n_1275, n_113, n_712, n_246, n_1042, n_269, n_285, n_412, n_657, n_644, n_1160, n_491, n_1258, n_1074, n_251, n_160, n_566, n_565, n_597, n_1181, n_1196, n_651, n_1340, n_334, n_811, n_807, n_835, n_175, n_666, n_262, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1018, n_438, n_713, n_904, n_166, n_1180, n_1271, n_533, n_1251, n_278, n_4251);

input n_924;
input n_1263;
input n_977;
input n_611;
input n_1126;
input n_1166;
input n_469;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1150;
input n_226;
input n_667;
input n_790;
input n_1055;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1292;
input n_1198;
input n_1360;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_1323;
input n_688;
input n_1353;
input n_800;
input n_1347;
input n_671;
input n_819;
input n_1022;
input n_915;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_292;
input n_625;
input n_854;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_755;
input n_1118;
input n_6;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_1314;
input n_709;
input n_317;
input n_1236;
input n_569;
input n_227;
input n_920;
input n_1289;
input n_94;
input n_335;
input n_370;
input n_976;
input n_343;
input n_308;
input n_297;
input n_156;
input n_1078;
input n_775;
input n_219;
input n_157;
input n_600;
input n_1328;
input n_223;
input n_264;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_436;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_496;
input n_958;
input n_1034;
input n_670;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1284;
input n_214;
input n_675;
input n_888;
input n_1167;
input n_637;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_197;
input n_1069;
input n_1075;
input n_1322;
input n_460;
input n_889;
input n_973;
input n_477;
input n_571;
input n_461;
input n_1211;
input n_1197;
input n_907;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_440;
input n_793;
input n_478;
input n_476;
input n_534;
input n_884;
input n_345;
input n_944;
input n_91;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_1319;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_596;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_409;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_434;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_1293;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_64;
input n_759;
input n_28;
input n_806;
input n_324;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_706;
input n_746;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_776;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_649;
input n_547;
input n_43;
input n_1191;
input n_116;
input n_284;
input n_1128;
input n_139;
input n_744;
input n_590;
input n_629;
input n_1308;
input n_254;
input n_1233;
input n_23;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1008;
input n_946;
input n_1001;
input n_498;
input n_689;
input n_738;
input n_640;
input n_252;
input n_624;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1158;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1049;
input n_1153;
input n_741;
input n_1306;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_1362;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_9;
input n_592;
input n_1169;
input n_45;
input n_1017;
input n_123;
input n_978;
input n_1054;
input n_1269;
input n_1095;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_484;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_374;
input n_185;
input n_396;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_723;
input n_1065;
input n_1336;
input n_473;
input n_1309;
input n_1043;
input n_355;
input n_486;
input n_614;
input n_337;
input n_88;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1132;
input n_388;
input n_1300;
input n_1127;
input n_761;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_582;
input n_1332;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_84;
input n_130;
input n_322;
input n_1249;
input n_652;
input n_1111;
input n_25;
input n_1349;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_44;
input n_224;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1304;
input n_1324;
input n_987;
input n_261;
input n_174;
input n_767;
input n_993;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_83;
input n_513;
input n_1094;
input n_1354;
input n_560;
input n_340;
input n_1351;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_495;
input n_602;
input n_574;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_490;
input n_1327;
input n_996;
input n_921;
input n_233;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1037;
input n_1080;
input n_1274;
input n_1316;
input n_426;
input n_1082;
input n_589;
input n_716;
input n_562;
input n_62;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_162;
input n_960;
input n_222;
input n_1290;
input n_1123;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_1311;
input n_256;
input n_950;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_376;
input n_967;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1357;
input n_483;
input n_683;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_983;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1343;
input n_1203;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1301;
input n_1363;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_1329;
input n_1312;
input n_804;
input n_537;
input n_945;
input n_492;
input n_153;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_883;
input n_470;
input n_325;
input n_449;
input n_132;
input n_1214;
input n_1342;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_13;
input n_1077;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_831;
input n_964;
input n_1350;
input n_1096;
input n_234;
input n_833;
input n_5;
input n_225;
input n_1307;
input n_988;
input n_814;
input n_192;
input n_1201;
input n_1114;
input n_655;
input n_669;
input n_472;
input n_1176;
input n_387;
input n_1149;
input n_398;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_1296;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_445;
input n_749;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_1338;
input n_577;
input n_338;
input n_149;
input n_693;
input n_14;
input n_836;
input n_990;
input n_975;
input n_1256;
input n_567;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1102;
input n_711;
input n_85;
input n_1187;
input n_1164;
input n_489;
input n_1174;
input n_617;
input n_1303;
input n_876;
input n_1190;
input n_118;
input n_601;
input n_917;
input n_966;
input n_253;
input n_1116;
input n_1212;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_818;
input n_861;
input n_1183;
input n_899;
input n_1253;
input n_210;
input n_774;
input n_1335;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_557;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_393;
input n_108;
input n_487;
input n_665;
input n_66;
input n_177;
input n_421;
input n_1356;
input n_910;
input n_768;
input n_1302;
input n_205;
input n_1136;
input n_1313;
input n_754;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_1310;
input n_202;
input n_427;
input n_791;
input n_732;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_148;
input n_435;
input n_159;
input n_766;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1155;
input n_89;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1352;
input n_626;
input n_1144;
input n_1137;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_194;
input n_855;
input n_1178;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_605;
input n_1273;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_1318;
input n_780;
input n_998;
input n_467;
input n_1227;
input n_840;
input n_1334;
input n_501;
input n_823;
input n_245;
input n_725;
input n_1295;
input n_672;
input n_581;
input n_382;
input n_554;
input n_898;
input n_1013;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_909;
input n_997;
input n_932;
input n_612;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_1320;
input n_737;
input n_986;
input n_509;
input n_1317;
input n_147;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_733;
input n_941;
input n_981;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1108;
input n_782;
input n_1100;
input n_862;
input n_760;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_31;
input n_481;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_1341;
input n_570;
input n_1361;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1225;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_221;
input n_622;
input n_1087;
input n_386;
input n_994;
input n_848;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_591;
input n_145;
input n_1344;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_432;
input n_839;
input n_1210;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_78;
input n_772;
input n_499;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_236;
input n_1012;
input n_1;
input n_1348;
input n_903;
input n_740;
input n_203;
input n_384;
input n_80;
input n_35;
input n_1315;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_1298;
input n_462;
input n_1193;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_40;
input n_1028;
input n_781;
input n_474;
input n_542;
input n_463;
input n_595;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_632;
input n_699;
input n_979;
input n_1245;
input n_846;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1103;
input n_648;
input n_312;
input n_1076;
input n_1091;
input n_494;
input n_641;
input n_730;
input n_1325;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1220;
input n_37;
input n_229;
input n_437;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_863;
input n_805;
input n_1275;
input n_113;
input n_712;
input n_246;
input n_1042;
input n_269;
input n_285;
input n_412;
input n_657;
input n_644;
input n_1160;
input n_491;
input n_1258;
input n_1074;
input n_251;
input n_160;
input n_566;
input n_565;
input n_597;
input n_1181;
input n_1196;
input n_651;
input n_1340;
input n_334;
input n_811;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1018;
input n_438;
input n_713;
input n_904;
input n_166;
input n_1180;
input n_1271;
input n_533;
input n_1251;
input n_278;

output n_4251;

wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_3912;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_4129;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_2955;
wire n_2899;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_3906;
wire n_4127;
wire n_4138;
wire n_3086;
wire n_3297;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_4217;
wire n_2683;
wire n_1370;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_2388;
wire n_2568;
wire n_3641;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3766;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4238;
wire n_1451;
wire n_4038;
wire n_2302;
wire n_4109;
wire n_2374;
wire n_1545;
wire n_3341;
wire n_1947;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4227;
wire n_4033;
wire n_2538;
wire n_2105;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1686;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_2543;
wire n_1860;
wire n_4155;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_3036;
wire n_2482;
wire n_3891;
wire n_4145;
wire n_2677;
wire n_4144;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_3532;
wire n_2770;
wire n_3987;
wire n_4061;
wire n_4131;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_1705;
wire n_2584;
wire n_2639;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_1698;
wire n_3880;
wire n_2329;
wire n_2963;
wire n_3834;
wire n_3624;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_3283;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_2091;
wire n_2466;
wire n_1517;
wire n_2652;
wire n_2635;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_2149;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_3947;
wire n_3490;
wire n_3656;
wire n_2071;
wire n_1484;
wire n_2643;
wire n_1374;
wire n_2561;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_2384;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_4135;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1547;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_3985;
wire n_1801;
wire n_1391;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_3744;
wire n_2235;
wire n_1862;
wire n_3980;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_2551;
wire n_1796;
wire n_3291;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_1521;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2506;
wire n_2699;
wire n_4064;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_3550;
wire n_1626;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_2118;
wire n_2985;
wire n_2944;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_2358;
wire n_3986;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3837;
wire n_1971;
wire n_1599;
wire n_3936;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_3096;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_2544;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_4069;
wire n_1667;
wire n_3359;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_3470;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_4195;
wire n_4218;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_3781;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_3328;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_3433;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_2305;
wire n_3392;
wire n_3430;
wire n_3975;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_3992;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_4148;
wire n_4151;
wire n_1883;
wire n_1906;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_4160;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_3989;
wire n_2837;
wire n_3804;
wire n_4051;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_3655;
wire n_2808;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_1538;
wire n_2930;
wire n_4206;
wire n_1838;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_2434;
wire n_1884;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_2967;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_3923;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_2454;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_2801;
wire n_3120;
wire n_1876;
wire n_4007;
wire n_1743;
wire n_3790;
wire n_4011;
wire n_3491;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_1888;
wire n_2009;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_2690;
wire n_4082;
wire n_4028;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_1690;
wire n_3819;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_2064;
wire n_3978;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_3500;
wire n_2413;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_1759;
wire n_2491;
wire n_2177;
wire n_1788;
wire n_3747;
wire n_1537;
wire n_3833;
wire n_3775;
wire n_2227;
wire n_4133;
wire n_2671;
wire n_4184;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_2022;
wire n_1798;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_3484;
wire n_3620;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_2469;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_3855;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1994;
wire n_3113;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_2960;
wire n_1500;
wire n_2796;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_3205;
wire n_4156;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_3856;
wire n_2145;
wire n_1639;
wire n_3703;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_3271;
wire n_2039;
wire n_4086;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_3753;
wire n_2084;
wire n_1781;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_3396;
wire n_3701;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_2320;
wire n_2339;
wire n_2473;
wire n_2038;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_3767;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_2847;
wire n_2051;
wire n_2029;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_4232;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_2457;
wire n_2346;
wire n_2312;
wire n_3990;
wire n_3475;
wire n_3015;
wire n_4170;
wire n_1578;
wire n_1920;
wire n_2536;
wire n_1592;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_2338;
wire n_1758;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_3730;
wire n_3883;
wire n_3276;
wire n_2565;
wire n_4152;
wire n_3897;
wire n_3845;
wire n_3787;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_3149;
wire n_2156;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_2418;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_2111;
wire n_2521;
wire n_1724;
wire n_3301;
wire n_3466;
wire n_3458;
wire n_1420;
wire n_3185;
wire n_3330;
wire n_1366;
wire n_3960;
wire n_2595;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_3586;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_2033;
wire n_1591;
wire n_4071;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_3399;
wire n_2896;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_2400;
wire n_3645;
wire n_3838;
wire n_3223;
wire n_1909;
wire n_3929;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_3474;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_3984;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_3679;
wire n_3779;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_2831;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_4110;
wire n_2803;
wire n_2851;
wire n_3707;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_1961;
wire n_4037;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_2436;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_4015;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_2301;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_3961;
wire n_2122;
wire n_1630;
wire n_2512;
wire n_3589;
wire n_4102;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1437;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_1424;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_3886;
wire n_1467;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_3860;
wire n_1382;
wire n_3546;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_2191;
wire n_2969;
wire n_2864;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_3053;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3548;
wire n_2440;
wire n_1699;
wire n_1386;
wire n_3334;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_3953;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_4003;
wire n_3800;
wire n_2402;
wire n_3073;
wire n_2403;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_3749;
wire n_3178;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1644;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_2475;
wire n_2733;
wire n_1719;
wire n_2993;
wire n_3864;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_3417;
wire n_3482;
wire n_2903;
wire n_3866;
wire n_3921;
wire n_1967;
wire n_2233;
wire n_1579;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1439;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_3734;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_1400;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_3529;
wire n_3854;
wire n_2169;
wire n_1804;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_4201;
wire n_1610;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_1636;
wire n_3253;
wire n_2056;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1865;
wire n_1511;
wire n_2973;
wire n_1470;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_2318;
wire n_2393;
wire n_1697;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_3372;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_2707;
wire n_2751;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_3950;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_2285;
wire n_1446;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_3869;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_2795;
wire n_4091;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_2098;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_3697;
wire n_2361;
wire n_3393;
wire n_1603;
wire n_4247;
wire n_2638;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1998;
wire n_3759;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_2034;
wire n_1637;
wire n_1419;
wire n_2711;
wire n_3933;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_2259;
wire n_1702;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_4068;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_2097;
wire n_1834;
wire n_1659;
wire n_2313;
wire n_2542;
wire n_3324;
wire n_2431;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_3736;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_3450;
wire n_1714;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_3174;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_2217;
wire n_3746;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_2745;
wire n_2201;
wire n_1737;
wire n_2722;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_3090;
wire n_2067;
wire n_2437;
wire n_2219;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1774;
wire n_1725;
wire n_3972;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_2532;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1991;
wire n_2224;
wire n_1399;
wire n_1979;
wire n_1543;
wire n_3368;
wire n_1533;
wire n_2924;
wire n_3467;
wire n_2484;
wire n_4111;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_3928;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_2264;
wire n_2754;
wire n_3534;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_2489;
wire n_3970;
wire n_3757;
wire n_3438;
wire n_4098;
wire n_2012;
wire n_3792;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_2245;
wire n_1782;
wire n_3561;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_2184;
wire n_2917;
wire n_1855;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_2965;
wire n_3635;
wire n_4150;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_3973;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_3934;
wire n_2213;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_3968;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1461;
wire n_2697;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1783;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1531;
wire n_1907;
wire n_3600;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_3239;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_4220;
wire n_1683;
wire n_1817;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_3431;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_2996;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1663;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_2315;
wire n_3228;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_2221;
wire n_3576;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_2326;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_2448;
wire n_3140;
wire n_3852;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_2898;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_3584;
wire n_1425;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_2447;
wire n_1813;
wire n_3761;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_2345;
wire n_2986;
wire n_2535;
wire n_4205;
wire n_2774;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_2376;
wire n_2488;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_3904;
wire n_2778;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_2691;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_1567;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_1648;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_2041;
wire n_3627;
wire n_3840;
wire n_1478;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_3903;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_2173;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_3464;
wire n_2018;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_3428;
wire n_2961;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1396;
wire n_2744;
wire n_2030;
wire n_2453;
wire n_2883;
wire n_1752;
wire n_1525;
wire n_2397;
wire n_3115;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_2234;
wire n_3251;
wire n_1910;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2050;
wire n_2809;
wire n_2797;
wire n_1676;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_3384;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1495;
wire n_4231;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_3250;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_3114;
wire n_2594;
wire n_3125;
wire n_3234;
wire n_2394;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_2823;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_3930;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_4212;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1397;
wire n_4057;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4245;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_1879;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1505;
wire n_4222;
wire n_4216;
wire n_1634;
wire n_3939;
wire n_4012;
wire n_2019;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_1558;
wire n_4241;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_3594;
wire n_1433;
wire n_2256;
wire n_1704;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_3799;
wire n_4119;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_2109;
wire n_2044;
wire n_2013;
wire n_2689;
wire n_1990;
wire n_2920;
wire n_3259;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_3693;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_569),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_740),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_638),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_114),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_872),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_341),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_745),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_304),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_492),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_889),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1006),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_892),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_590),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1275),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_440),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_703),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_90),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1213),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1229),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_165),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1303),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1242),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_58),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1221),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_383),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1280),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_385),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_934),
.Y(n_1391)
);

BUFx5_ASAP7_75t_L g1392 ( 
.A(n_850),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_469),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_399),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_818),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_516),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_290),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1336),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1048),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_221),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_278),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1186),
.Y(n_1402)
);

BUFx10_ASAP7_75t_L g1403 ( 
.A(n_1225),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_125),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_675),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1222),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1128),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1308),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_84),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_597),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_995),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_164),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_807),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_531),
.Y(n_1414)
);

BUFx10_ASAP7_75t_L g1415 ( 
.A(n_537),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1253),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1145),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_937),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1276),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1015),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_529),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_415),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1011),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_937),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1282),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1236),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_230),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1027),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1043),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1275),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1307),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_916),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1053),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1076),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_593),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_496),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_367),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1230),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1322),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1221),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_947),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_351),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_315),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_240),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_886),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_621),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_960),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_958),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1168),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_25),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1315),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_640),
.Y(n_1452)
);

BUFx10_ASAP7_75t_L g1453 ( 
.A(n_1255),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1239),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1087),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1044),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_270),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_500),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_391),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1108),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1310),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1156),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_583),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1258),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_960),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1088),
.Y(n_1466)
);

BUFx10_ASAP7_75t_L g1467 ( 
.A(n_1113),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_478),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_823),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_852),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1312),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_796),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_301),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1360),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_890),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_48),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_94),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_414),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_37),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1316),
.Y(n_1480)
);

BUFx2_ASAP7_75t_SL g1481 ( 
.A(n_1268),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1313),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_795),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_327),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1306),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_465),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_827),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1362),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_184),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1213),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_249),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_116),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1270),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1132),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1045),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1227),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_307),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1123),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_712),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1342),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1226),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1217),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_250),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_424),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_253),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_387),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_608),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_210),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_334),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_550),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_787),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_412),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_887),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1254),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_242),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_329),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_920),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1271),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1265),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_897),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_532),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_90),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1283),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_96),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_750),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_946),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_303),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_829),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1257),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1234),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_435),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1244),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_253),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1107),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_919),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1273),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1291),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_880),
.Y(n_1538)
);

BUFx10_ASAP7_75t_L g1539 ( 
.A(n_801),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_698),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1143),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_627),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1257),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_643),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_290),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_656),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_853),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1111),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_775),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1317),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_580),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1248),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_771),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_983),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1262),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1318),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_63),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1272),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1297),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1126),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_371),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1262),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_243),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_862),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1332),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_992),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_596),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1202),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1311),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1039),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_12),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_631),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1237),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1260),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1264),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1277),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1000),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_462),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_394),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_362),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1286),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_392),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_108),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1320),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1062),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1301),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_198),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1321),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1333),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_796),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1222),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1256),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_654),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_323),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_982),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1214),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_912),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_934),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1241),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1144),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_70),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_163),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_563),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_472),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_561),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_111),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1355),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_949),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1243),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_590),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1073),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1292),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_979),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_158),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_274),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_93),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1063),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1216),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_945),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_173),
.Y(n_1620)
);

BUFx5_ASAP7_75t_L g1621 ( 
.A(n_566),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_388),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1155),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1309),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1259),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_378),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1362),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_619),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_542),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1240),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1235),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_220),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_847),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_96),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_858),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1020),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_740),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_542),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1047),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1241),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_522),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_483),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1252),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1146),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1048),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1359),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1212),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_778),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_871),
.Y(n_1649)
);

BUFx10_ASAP7_75t_L g1650 ( 
.A(n_1070),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_517),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1266),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_201),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_626),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_1201),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_403),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_232),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1187),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1194),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1285),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_923),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_317),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1105),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_343),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1174),
.Y(n_1665)
);

CKINVDCx14_ASAP7_75t_R g1666 ( 
.A(n_541),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1121),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_224),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1298),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1251),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_479),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_499),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1334),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_268),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1289),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_553),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1290),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1261),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1326),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_431),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1326),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_662),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_137),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_429),
.Y(n_1684)
);

INVx4_ASAP7_75t_R g1685 ( 
.A(n_1253),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_731),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1219),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1054),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_276),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_319),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1295),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1140),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_870),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_846),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1279),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_814),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1072),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_222),
.Y(n_1698)
);

CKINVDCx16_ASAP7_75t_R g1699 ( 
.A(n_581),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1089),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_83),
.Y(n_1701)
);

BUFx10_ASAP7_75t_L g1702 ( 
.A(n_431),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_632),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1071),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1129),
.Y(n_1705)
);

BUFx2_ASAP7_75t_SL g1706 ( 
.A(n_1288),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_518),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_624),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1018),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_236),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1232),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1101),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_972),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_918),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_468),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_611),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_37),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_409),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1042),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1061),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_69),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1314),
.Y(n_1722)
);

CKINVDCx14_ASAP7_75t_R g1723 ( 
.A(n_973),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_551),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_95),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_383),
.Y(n_1726)
);

INVx4_ASAP7_75t_R g1727 ( 
.A(n_113),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1163),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_398),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_766),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_879),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_160),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_244),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_309),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_723),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_601),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_633),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_159),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_697),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1038),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1082),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_286),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_59),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_190),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_845),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_957),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1300),
.Y(n_1747)
);

BUFx2_ASAP7_75t_SL g1748 ( 
.A(n_92),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1130),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1296),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1224),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1331),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_645),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_137),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_672),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_514),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1238),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_547),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_207),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_58),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_875),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_225),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1263),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1305),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1285),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_603),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_157),
.Y(n_1767)
);

BUFx8_ASAP7_75t_SL g1768 ( 
.A(n_1155),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_591),
.Y(n_1769)
);

BUFx10_ASAP7_75t_L g1770 ( 
.A(n_638),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1056),
.Y(n_1771)
);

CKINVDCx14_ASAP7_75t_R g1772 ( 
.A(n_574),
.Y(n_1772)
);

CKINVDCx16_ASAP7_75t_R g1773 ( 
.A(n_100),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_389),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_192),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_134),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1147),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_219),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_238),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_830),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1250),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1218),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_97),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_151),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_117),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_122),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_527),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1284),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_880),
.Y(n_1789)
);

BUFx5_ASAP7_75t_L g1790 ( 
.A(n_1304),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_240),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_813),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1287),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_95),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_741),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_277),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_255),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_28),
.Y(n_1798)
);

BUFx10_ASAP7_75t_L g1799 ( 
.A(n_1302),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_193),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1271),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1269),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1215),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_915),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_449),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_285),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_551),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1013),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1313),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_441),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_318),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1274),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1036),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_SL g1814 ( 
.A(n_657),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_404),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_614),
.Y(n_1816)
);

CKINVDCx20_ASAP7_75t_R g1817 ( 
.A(n_19),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_301),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_983),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_363),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1220),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1171),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_538),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1074),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1150),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_221),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_476),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1160),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_43),
.Y(n_1829)
);

BUFx5_ASAP7_75t_L g1830 ( 
.A(n_958),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_799),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_951),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_677),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1278),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1299),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_103),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1017),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_497),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1290),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_24),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1025),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1245),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_968),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1117),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_189),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_634),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_275),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1267),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_974),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_895),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_525),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_800),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_596),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_493),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1249),
.Y(n_1855)
);

BUFx10_ASAP7_75t_L g1856 ( 
.A(n_1004),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_15),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_166),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_803),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_336),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_211),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_223),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1009),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1223),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_192),
.Y(n_1865)
);

BUFx8_ASAP7_75t_SL g1866 ( 
.A(n_445),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_43),
.Y(n_1867)
);

CKINVDCx20_ASAP7_75t_R g1868 ( 
.A(n_35),
.Y(n_1868)
);

BUFx2_ASAP7_75t_SL g1869 ( 
.A(n_1293),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_993),
.Y(n_1870)
);

BUFx10_ASAP7_75t_L g1871 ( 
.A(n_1095),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_764),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1344),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_458),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_462),
.Y(n_1875)
);

CKINVDCx16_ASAP7_75t_R g1876 ( 
.A(n_867),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_128),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_689),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1348),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_37),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_99),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1207),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_675),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_765),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1016),
.Y(n_1885)
);

BUFx10_ASAP7_75t_L g1886 ( 
.A(n_520),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_829),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_166),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1294),
.Y(n_1889)
);

BUFx10_ASAP7_75t_L g1890 ( 
.A(n_481),
.Y(n_1890)
);

INVxp33_ASAP7_75t_R g1891 ( 
.A(n_1341),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_486),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1055),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_6),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_721),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1000),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_718),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1012),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_669),
.Y(n_1899)
);

BUFx10_ASAP7_75t_L g1900 ( 
.A(n_773),
.Y(n_1900)
);

CKINVDCx20_ASAP7_75t_R g1901 ( 
.A(n_206),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1281),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_227),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1242),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1119),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1233),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_581),
.Y(n_1907)
);

CKINVDCx16_ASAP7_75t_R g1908 ( 
.A(n_575),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_11),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_180),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_93),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1228),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1170),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1231),
.Y(n_1914)
);

BUFx10_ASAP7_75t_L g1915 ( 
.A(n_338),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_174),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_1008),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_640),
.Y(n_1918)
);

BUFx5_ASAP7_75t_L g1919 ( 
.A(n_266),
.Y(n_1919)
);

BUFx2_ASAP7_75t_SL g1920 ( 
.A(n_418),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_255),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_387),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_281),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_896),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_886),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1049),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_788),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_1080),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_362),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_168),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1263),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_16),
.Y(n_1932)
);

CKINVDCx14_ASAP7_75t_R g1933 ( 
.A(n_1246),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1247),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_864),
.Y(n_1935)
);

CKINVDCx20_ASAP7_75t_R g1936 ( 
.A(n_1933),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1524),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1392),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1392),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1392),
.Y(n_1940)
);

INVxp33_ASAP7_75t_L g1941 ( 
.A(n_1653),
.Y(n_1941)
);

BUFx10_ASAP7_75t_L g1942 ( 
.A(n_1367),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1621),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1621),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1621),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1790),
.Y(n_1946)
);

INVxp67_ASAP7_75t_SL g1947 ( 
.A(n_1722),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1666),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1790),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1394),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1790),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1830),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1830),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1459),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1830),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1768),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1866),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1773),
.Y(n_1958)
);

CKINVDCx20_ASAP7_75t_R g1959 ( 
.A(n_1723),
.Y(n_1959)
);

CKINVDCx14_ASAP7_75t_R g1960 ( 
.A(n_1772),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1919),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1919),
.Y(n_1962)
);

CKINVDCx20_ASAP7_75t_R g1963 ( 
.A(n_1388),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1754),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1383),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1655),
.Y(n_1966)
);

INVxp33_ASAP7_75t_SL g1967 ( 
.A(n_1374),
.Y(n_1967)
);

CKINVDCx16_ASAP7_75t_R g1968 ( 
.A(n_1699),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1444),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1412),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1476),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1903),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1587),
.Y(n_1973)
);

INVxp33_ASAP7_75t_L g1974 ( 
.A(n_1391),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1601),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1876),
.Y(n_1976)
);

CKINVDCx20_ASAP7_75t_R g1977 ( 
.A(n_1908),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1698),
.Y(n_1978)
);

INVxp33_ASAP7_75t_L g1979 ( 
.A(n_1429),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1701),
.Y(n_1980)
);

NOR2xp67_ASAP7_75t_L g1981 ( 
.A(n_1844),
.B(n_0),
.Y(n_1981)
);

INVxp33_ASAP7_75t_SL g1982 ( 
.A(n_1780),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1738),
.Y(n_1983)
);

CKINVDCx20_ASAP7_75t_R g1984 ( 
.A(n_1382),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1760),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1779),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1783),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1786),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1380),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1791),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1836),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1840),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1857),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1867),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1877),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1888),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1387),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1386),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1393),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1894),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1412),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1498),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1657),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1657),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1794),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1794),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1634),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1394),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1394),
.Y(n_2009)
);

BUFx3_ASAP7_75t_L g2010 ( 
.A(n_1402),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1430),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1430),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1400),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1472),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1404),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1472),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1528),
.Y(n_2017)
);

CKINVDCx16_ASAP7_75t_R g2018 ( 
.A(n_1814),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1682),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1409),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1682),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_1682),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1421),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1709),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1709),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1709),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_1740),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_1673),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1427),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1440),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1747),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1747),
.Y(n_2032)
);

INVxp33_ASAP7_75t_L g2033 ( 
.A(n_1690),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1769),
.Y(n_2034)
);

INVxp67_ASAP7_75t_SL g2035 ( 
.A(n_1807),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1812),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1456),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_1917),
.Y(n_2038)
);

INVxp33_ASAP7_75t_SL g2039 ( 
.A(n_1450),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1477),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1833),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1479),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1853),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1405),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_1930),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1492),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1417),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_1426),
.Y(n_2048)
);

NOR2xp67_ASAP7_75t_L g2049 ( 
.A(n_1436),
.B(n_0),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1503),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1508),
.Y(n_2051)
);

INVx1_ASAP7_75t_SL g2052 ( 
.A(n_1935),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1569),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1675),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1678),
.Y(n_2055)
);

INVxp67_ASAP7_75t_SL g2056 ( 
.A(n_1687),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1695),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1703),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1708),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1728),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1731),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1749),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1804),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1815),
.Y(n_2064)
);

INVxp67_ASAP7_75t_SL g2065 ( 
.A(n_1863),
.Y(n_2065)
);

INVxp67_ASAP7_75t_SL g2066 ( 
.A(n_1899),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1557),
.Y(n_2067)
);

INVxp33_ASAP7_75t_SL g2068 ( 
.A(n_1571),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_1379),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1931),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1934),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1583),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1366),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1925),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1926),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1602),
.Y(n_2076)
);

BUFx2_ASAP7_75t_L g2077 ( 
.A(n_1606),
.Y(n_2077)
);

INVxp67_ASAP7_75t_SL g2078 ( 
.A(n_1437),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1403),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1368),
.Y(n_2080)
);

OA21x2_ASAP7_75t_L g2081 ( 
.A1(n_1938),
.A2(n_1469),
.B(n_1435),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1970),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2017),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1960),
.B(n_1460),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2022),
.Y(n_2085)
);

OA21x2_ASAP7_75t_L g2086 ( 
.A1(n_1939),
.A2(n_1478),
.B(n_1471),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_2018),
.Y(n_2087)
);

BUFx2_ASAP7_75t_L g2088 ( 
.A(n_1963),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1970),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1967),
.A2(n_1614),
.B1(n_1620),
.B2(n_1616),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2027),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1947),
.B(n_1705),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1937),
.B(n_1725),
.Y(n_2093)
);

CKINVDCx8_ASAP7_75t_R g2094 ( 
.A(n_1968),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2035),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_2079),
.B(n_1411),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_2069),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2001),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2003),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_2069),
.Y(n_2100)
);

OAI21x1_ASAP7_75t_L g2101 ( 
.A1(n_1940),
.A2(n_1514),
.B(n_1491),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2004),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2005),
.Y(n_2103)
);

BUFx12f_ASAP7_75t_L g2104 ( 
.A(n_1956),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2006),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1954),
.B(n_2002),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1982),
.A2(n_1683),
.B1(n_1710),
.B2(n_1668),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2008),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_2039),
.B(n_1717),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2048),
.B(n_1721),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2009),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2056),
.B(n_1527),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1950),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2065),
.B(n_1406),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2011),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1957),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2012),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2014),
.Y(n_2118)
);

BUFx3_ASAP7_75t_L g2119 ( 
.A(n_1964),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2016),
.Y(n_2120)
);

CKINVDCx16_ASAP7_75t_R g2121 ( 
.A(n_1936),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_1942),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1972),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2066),
.B(n_1743),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2077),
.B(n_1406),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_2068),
.B(n_1744),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_1942),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_SL g2128 ( 
.A1(n_1977),
.A2(n_1732),
.B1(n_1817),
.B2(n_1522),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2078),
.B(n_1759),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_1986),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1992),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1999),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_2010),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_2045),
.B(n_2028),
.Y(n_2134)
);

BUFx2_ASAP7_75t_L g2135 ( 
.A(n_1948),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2019),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1966),
.A2(n_1767),
.B1(n_1775),
.B2(n_1762),
.Y(n_2137)
);

BUFx3_ASAP7_75t_L g2138 ( 
.A(n_2047),
.Y(n_2138)
);

BUFx12f_ASAP7_75t_L g2139 ( 
.A(n_1958),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2021),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2024),
.Y(n_2141)
);

OAI22x1_ASAP7_75t_SL g2142 ( 
.A1(n_1984),
.A2(n_1868),
.B1(n_1901),
.B2(n_1865),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_2025),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2026),
.Y(n_2144)
);

XOR2xp5_ASAP7_75t_L g2145 ( 
.A(n_1997),
.B(n_1488),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2031),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1989),
.B(n_1776),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_2032),
.Y(n_2148)
);

CKINVDCx6p67_ASAP7_75t_R g2149 ( 
.A(n_1959),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_1998),
.Y(n_2150)
);

BUFx6f_ASAP7_75t_L g2151 ( 
.A(n_2034),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_2036),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2041),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_2013),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_2044),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_2050),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_2043),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1965),
.Y(n_2158)
);

AND2x6_ASAP7_75t_L g2159 ( 
.A(n_2053),
.B(n_1489),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2015),
.B(n_1415),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2020),
.B(n_2029),
.Y(n_2161)
);

OAI21x1_ASAP7_75t_L g2162 ( 
.A1(n_1943),
.A2(n_1777),
.B(n_1752),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1945),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1944),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1946),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1949),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2038),
.A2(n_1778),
.B1(n_1785),
.B2(n_1784),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2052),
.A2(n_1800),
.B1(n_1826),
.B2(n_1798),
.Y(n_2168)
);

BUFx3_ASAP7_75t_L g2169 ( 
.A(n_2054),
.Y(n_2169)
);

OA21x2_ASAP7_75t_L g2170 ( 
.A1(n_1951),
.A2(n_1847),
.B(n_1841),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1952),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1969),
.Y(n_2172)
);

AND2x4_ASAP7_75t_SL g2173 ( 
.A(n_1976),
.B(n_1453),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1953),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1955),
.Y(n_2175)
);

AND2x6_ASAP7_75t_L g2176 ( 
.A(n_2055),
.B(n_2057),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_2040),
.A2(n_2046),
.B1(n_2051),
.B2(n_2042),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1961),
.Y(n_2178)
);

OA21x2_ASAP7_75t_L g2179 ( 
.A1(n_1962),
.A2(n_1921),
.B(n_1902),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2067),
.B(n_1829),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1971),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2070),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2072),
.B(n_1845),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2076),
.B(n_1858),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2071),
.Y(n_2185)
);

BUFx2_ASAP7_75t_L g2186 ( 
.A(n_2023),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_2058),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2073),
.Y(n_2188)
);

BUFx8_ASAP7_75t_SL g2189 ( 
.A(n_2030),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_2059),
.B(n_1369),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2060),
.B(n_1861),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_2061),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_2189),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2138),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_2154),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_2177),
.B(n_2109),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2092),
.B(n_1981),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2182),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2185),
.Y(n_2199)
);

CKINVDCx16_ASAP7_75t_R g2200 ( 
.A(n_2121),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_SL g2201 ( 
.A(n_2122),
.Y(n_2201)
);

CKINVDCx20_ASAP7_75t_R g2202 ( 
.A(n_2087),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_2097),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2188),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_2116),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2100),
.Y(n_2206)
);

CKINVDCx20_ASAP7_75t_R g2207 ( 
.A(n_2149),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2158),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2089),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_2132),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_2104),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_2139),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_2150),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_2186),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_2094),
.Y(n_2215)
);

CKINVDCx16_ASAP7_75t_R g2216 ( 
.A(n_2145),
.Y(n_2216)
);

NAND2xp33_ASAP7_75t_R g2217 ( 
.A(n_2088),
.B(n_1862),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_R g2218 ( 
.A(n_2127),
.B(n_2037),
.Y(n_2218)
);

AO22x2_ASAP7_75t_L g2219 ( 
.A1(n_2090),
.A2(n_1748),
.B1(n_1706),
.B2(n_1481),
.Y(n_2219)
);

CKINVDCx20_ASAP7_75t_R g2220 ( 
.A(n_2135),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_2161),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2125),
.B(n_2033),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_SL g2223 ( 
.A1(n_2128),
.A2(n_1495),
.B1(n_1534),
.B2(n_1493),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_2082),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2123),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2083),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_R g2227 ( 
.A(n_2085),
.B(n_2091),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_2133),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_2126),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2172),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_2147),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2180),
.Y(n_2232)
);

BUFx3_ASAP7_75t_L g2233 ( 
.A(n_2155),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_R g2234 ( 
.A(n_2095),
.B(n_2062),
.Y(n_2234)
);

AOI21x1_ASAP7_75t_L g2235 ( 
.A1(n_2165),
.A2(n_2075),
.B(n_2074),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_R g2236 ( 
.A(n_2183),
.B(n_2063),
.Y(n_2236)
);

BUFx3_ASAP7_75t_L g2237 ( 
.A(n_2156),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_2160),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2181),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_2113),
.Y(n_2240)
);

INVxp33_ASAP7_75t_SL g2241 ( 
.A(n_2168),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2114),
.B(n_1941),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_2142),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_2137),
.Y(n_2244)
);

BUFx10_ASAP7_75t_L g2245 ( 
.A(n_2106),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2110),
.B(n_1974),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_2124),
.Y(n_2247)
);

BUFx3_ASAP7_75t_L g2248 ( 
.A(n_2169),
.Y(n_2248)
);

CKINVDCx20_ASAP7_75t_R g2249 ( 
.A(n_2173),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_2084),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_2129),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_2107),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_2192),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2174),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2134),
.B(n_1979),
.Y(n_2255)
);

INVx1_ASAP7_75t_SL g2256 ( 
.A(n_2096),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2178),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_2167),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_R g2259 ( 
.A(n_2191),
.B(n_2064),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_2159),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2164),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2166),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2159),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_2112),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2163),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2171),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2093),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_2176),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_2130),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_2131),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_2081),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2143),
.Y(n_2272)
);

INVxp67_ASAP7_75t_L g2273 ( 
.A(n_2151),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2175),
.Y(n_2274)
);

BUFx2_ASAP7_75t_L g2275 ( 
.A(n_2190),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_2152),
.Y(n_2276)
);

CKINVDCx5p33_ASAP7_75t_R g2277 ( 
.A(n_2157),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2103),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2105),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2187),
.B(n_1973),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2086),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2140),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2148),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_2153),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_2101),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_R g2286 ( 
.A(n_2098),
.B(n_1538),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2108),
.B(n_2111),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2099),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_R g2289 ( 
.A(n_2102),
.B(n_1552),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_2115),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2170),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_2117),
.Y(n_2292)
);

BUFx2_ASAP7_75t_L g2293 ( 
.A(n_2179),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2118),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_2120),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_2136),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2141),
.B(n_2049),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2144),
.B(n_1975),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2146),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2162),
.B(n_1978),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_R g2301 ( 
.A(n_2087),
.B(n_1560),
.Y(n_2301)
);

BUFx6f_ASAP7_75t_SL g2302 ( 
.A(n_2122),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_2189),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_2097),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2147),
.B(n_1880),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_2132),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_2119),
.B(n_1980),
.Y(n_2307)
);

CKINVDCx20_ASAP7_75t_R g2308 ( 
.A(n_2189),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2138),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2110),
.B(n_1983),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2189),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_2184),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2251),
.B(n_1364),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2312),
.B(n_1891),
.Y(n_2314)
);

NOR2x1p5_ASAP7_75t_L g2315 ( 
.A(n_2263),
.B(n_1881),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2300),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2287),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2198),
.Y(n_2318)
);

INVx4_ASAP7_75t_L g2319 ( 
.A(n_2272),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2222),
.B(n_1985),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2210),
.B(n_1987),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2199),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_2240),
.Y(n_2323)
);

OR2x6_ASAP7_75t_L g2324 ( 
.A(n_2306),
.B(n_1869),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2231),
.B(n_2080),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_2225),
.B(n_1988),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2204),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2232),
.B(n_1990),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2247),
.B(n_1407),
.Y(n_2329)
);

BUFx3_ASAP7_75t_L g2330 ( 
.A(n_2269),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2298),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2240),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2305),
.B(n_2197),
.Y(n_2333)
);

AND2x2_ASAP7_75t_SL g2334 ( 
.A(n_2260),
.B(n_1370),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2221),
.B(n_1420),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_2240),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2246),
.B(n_2250),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_L g2338 ( 
.A1(n_2293),
.A2(n_1920),
.B1(n_1375),
.B2(n_1377),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2254),
.B(n_1991),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2294),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_2264),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2257),
.B(n_1993),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2299),
.Y(n_2343)
);

INVx4_ASAP7_75t_L g2344 ( 
.A(n_2276),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2226),
.Y(n_2345)
);

AND2x6_ASAP7_75t_L g2346 ( 
.A(n_2307),
.B(n_1632),
.Y(n_2346)
);

AO22x2_ASAP7_75t_L g2347 ( 
.A1(n_2223),
.A2(n_1484),
.B1(n_1531),
.B2(n_1462),
.Y(n_2347)
);

AND2x2_ASAP7_75t_SL g2348 ( 
.A(n_2200),
.B(n_1372),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2265),
.Y(n_2349)
);

AND2x6_ASAP7_75t_L g2350 ( 
.A(n_2233),
.B(n_1378),
.Y(n_2350)
);

INVx1_ASAP7_75t_SL g2351 ( 
.A(n_2286),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_2224),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2228),
.B(n_1994),
.Y(n_2353)
);

CKINVDCx20_ASAP7_75t_R g2354 ( 
.A(n_2202),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2237),
.B(n_1995),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2229),
.B(n_1533),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2224),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_2248),
.B(n_1996),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_2289),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2280),
.Y(n_2360)
);

INVx2_ASAP7_75t_SL g2361 ( 
.A(n_2245),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2241),
.B(n_1605),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_2203),
.Y(n_2363)
);

INVx4_ASAP7_75t_L g2364 ( 
.A(n_2277),
.Y(n_2364)
);

AND2x6_ASAP7_75t_L g2365 ( 
.A(n_2194),
.B(n_1384),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2203),
.Y(n_2366)
);

INVxp67_ASAP7_75t_L g2367 ( 
.A(n_2255),
.Y(n_2367)
);

OAI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2310),
.A2(n_1619),
.B1(n_1652),
.B2(n_1630),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2278),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2279),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2282),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2281),
.B(n_2000),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2288),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2261),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2236),
.B(n_1365),
.Y(n_2375)
);

NAND2xp33_ASAP7_75t_R g2376 ( 
.A(n_2301),
.B(n_1909),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_R g2377 ( 
.A(n_2193),
.B(n_1910),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2262),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_2206),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_2195),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_2206),
.Y(n_2381)
);

INVx5_ASAP7_75t_L g2382 ( 
.A(n_2206),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2266),
.Y(n_2383)
);

AND2x6_ASAP7_75t_L g2384 ( 
.A(n_2309),
.B(n_1385),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2209),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_2304),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2258),
.B(n_1684),
.Y(n_2387)
);

BUFx3_ASAP7_75t_L g2388 ( 
.A(n_2270),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_2273),
.B(n_2007),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2274),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2291),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2235),
.Y(n_2392)
);

INVx6_ASAP7_75t_L g2393 ( 
.A(n_2304),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2238),
.B(n_1467),
.Y(n_2394)
);

BUFx10_ASAP7_75t_L g2395 ( 
.A(n_2303),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2267),
.Y(n_2396)
);

INVx1_ASAP7_75t_SL g2397 ( 
.A(n_2220),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2285),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2290),
.B(n_1735),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2292),
.B(n_1808),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2285),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2227),
.B(n_1371),
.Y(n_2402)
);

INVx2_ASAP7_75t_SL g2403 ( 
.A(n_2234),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2295),
.B(n_1818),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2213),
.B(n_1467),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2275),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2208),
.B(n_1395),
.Y(n_2407)
);

INVx4_ASAP7_75t_L g2408 ( 
.A(n_2215),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2284),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2259),
.B(n_1373),
.Y(n_2410)
);

AOI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2219),
.A2(n_1398),
.B1(n_1399),
.B2(n_1397),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2283),
.B(n_1376),
.Y(n_2412)
);

AND2x6_ASAP7_75t_L g2413 ( 
.A(n_2230),
.B(n_1410),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2239),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2216),
.B(n_1872),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2296),
.B(n_1381),
.Y(n_2416)
);

BUFx6f_ASAP7_75t_L g2417 ( 
.A(n_2214),
.Y(n_2417)
);

INVxp33_ASAP7_75t_L g2418 ( 
.A(n_2218),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2253),
.Y(n_2419)
);

BUFx6f_ASAP7_75t_L g2420 ( 
.A(n_2212),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2297),
.Y(n_2421)
);

AND2x6_ASAP7_75t_L g2422 ( 
.A(n_2268),
.B(n_1414),
.Y(n_2422)
);

INVx4_ASAP7_75t_L g2423 ( 
.A(n_2211),
.Y(n_2423)
);

AND2x6_ASAP7_75t_L g2424 ( 
.A(n_2201),
.B(n_1418),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2244),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_2249),
.B(n_1419),
.Y(n_2426)
);

OR2x2_ASAP7_75t_SL g2427 ( 
.A(n_2252),
.B(n_1422),
.Y(n_2427)
);

AND2x6_ASAP7_75t_L g2428 ( 
.A(n_2302),
.B(n_1425),
.Y(n_2428)
);

INVx6_ASAP7_75t_L g2429 ( 
.A(n_2207),
.Y(n_2429)
);

INVx1_ASAP7_75t_SL g2430 ( 
.A(n_2205),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2243),
.Y(n_2431)
);

AND2x6_ASAP7_75t_L g2432 ( 
.A(n_2217),
.B(n_1428),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_2311),
.Y(n_2433)
);

AND2x6_ASAP7_75t_L g2434 ( 
.A(n_2308),
.B(n_1434),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2265),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2224),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2265),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2242),
.B(n_1539),
.Y(n_2438)
);

BUFx3_ASAP7_75t_L g2439 ( 
.A(n_2210),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2300),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2300),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2231),
.B(n_1389),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2231),
.B(n_1390),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2265),
.Y(n_2444)
);

HB1xp67_ASAP7_75t_L g2445 ( 
.A(n_2256),
.Y(n_2445)
);

INVxp67_ASAP7_75t_SL g2446 ( 
.A(n_2271),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_2210),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2300),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2231),
.B(n_1396),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2251),
.B(n_1401),
.Y(n_2450)
);

INVx4_ASAP7_75t_L g2451 ( 
.A(n_2272),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2210),
.B(n_1445),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2300),
.Y(n_2453)
);

AOI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2251),
.A2(n_1562),
.B1(n_1564),
.B2(n_1561),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2222),
.Y(n_2455)
);

INVx4_ASAP7_75t_L g2456 ( 
.A(n_2272),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2300),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_2272),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2242),
.B(n_1922),
.Y(n_2459)
);

NOR2x1p5_ASAP7_75t_L g2460 ( 
.A(n_2263),
.B(n_1911),
.Y(n_2460)
);

NAND2x1p5_ASAP7_75t_L g2461 ( 
.A(n_2233),
.B(n_1447),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2231),
.B(n_1408),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2312),
.B(n_1916),
.Y(n_2463)
);

AO22x2_ASAP7_75t_L g2464 ( 
.A1(n_2196),
.A2(n_1452),
.B1(n_1455),
.B2(n_1448),
.Y(n_2464)
);

CKINVDCx16_ASAP7_75t_R g2465 ( 
.A(n_2218),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2242),
.B(n_1650),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2265),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2333),
.B(n_1577),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2318),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2445),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2337),
.B(n_1603),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2446),
.B(n_1413),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2329),
.B(n_1416),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2335),
.B(n_1612),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2349),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2440),
.B(n_1423),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2441),
.B(n_1424),
.Y(n_2477)
);

OR2x2_ASAP7_75t_L g2478 ( 
.A(n_2459),
.B(n_1932),
.Y(n_2478)
);

INVx5_ASAP7_75t_L g2479 ( 
.A(n_2417),
.Y(n_2479)
);

HB1xp67_ASAP7_75t_L g2480 ( 
.A(n_2455),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2448),
.B(n_1431),
.Y(n_2481)
);

NAND3xp33_ASAP7_75t_SL g2482 ( 
.A(n_2454),
.B(n_1704),
.C(n_1693),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2453),
.B(n_1432),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2457),
.B(n_1433),
.Y(n_2484)
);

OR2x6_ASAP7_75t_L g2485 ( 
.A(n_2388),
.B(n_1461),
.Y(n_2485)
);

NOR2xp67_ASAP7_75t_SL g2486 ( 
.A(n_2403),
.B(n_1463),
.Y(n_2486)
);

INVx2_ASAP7_75t_SL g2487 ( 
.A(n_2393),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2322),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2435),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_2352),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2399),
.B(n_1702),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2357),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2437),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2327),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_2387),
.B(n_1789),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2340),
.Y(n_2496)
);

OR2x6_ASAP7_75t_L g2497 ( 
.A(n_2319),
.B(n_1464),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2444),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2360),
.B(n_1438),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_SL g2500 ( 
.A(n_2424),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2328),
.B(n_1439),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2325),
.B(n_1441),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2463),
.B(n_1442),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2343),
.Y(n_2504)
);

INVx8_ASAP7_75t_L g2505 ( 
.A(n_2382),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2391),
.B(n_1443),
.Y(n_2506)
);

INVxp67_ASAP7_75t_L g2507 ( 
.A(n_2400),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2317),
.B(n_2404),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2331),
.B(n_1446),
.Y(n_2509)
);

NAND2x1_ASAP7_75t_L g2510 ( 
.A(n_2398),
.B(n_1727),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_L g2511 ( 
.A1(n_2464),
.A2(n_1928),
.B1(n_1465),
.B2(n_1466),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2320),
.B(n_1702),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2372),
.B(n_1449),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2442),
.B(n_1451),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2443),
.B(n_1454),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2345),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2449),
.B(n_1457),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2467),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_2386),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2415),
.B(n_1458),
.Y(n_2520)
);

A2O1A1Ixp33_ASAP7_75t_L g2521 ( 
.A1(n_2338),
.A2(n_1483),
.B(n_1486),
.C(n_1475),
.Y(n_2521)
);

OAI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2401),
.A2(n_1470),
.B1(n_1473),
.B2(n_1468),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2462),
.B(n_1474),
.Y(n_2523)
);

AOI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2334),
.A2(n_1482),
.B1(n_1485),
.B2(n_1480),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2370),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2369),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2371),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2321),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2351),
.B(n_1490),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2402),
.B(n_2438),
.Y(n_2530)
);

NAND2x1_ASAP7_75t_L g2531 ( 
.A(n_2392),
.B(n_1685),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2390),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2373),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2374),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2378),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2383),
.Y(n_2536)
);

AND2x6_ASAP7_75t_SL g2537 ( 
.A(n_2314),
.B(n_1487),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2409),
.B(n_1494),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2466),
.B(n_1496),
.Y(n_2539)
);

HB1xp67_ASAP7_75t_L g2540 ( 
.A(n_2406),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2355),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2359),
.B(n_1497),
.Y(n_2542)
);

INVx2_ASAP7_75t_SL g2543 ( 
.A(n_2358),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2416),
.B(n_1499),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_L g2545 ( 
.A(n_2418),
.B(n_1501),
.Y(n_2545)
);

OAI221xp5_ASAP7_75t_L g2546 ( 
.A1(n_2411),
.A2(n_1507),
.B1(n_1509),
.B2(n_1502),
.C(n_1500),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2354),
.Y(n_2547)
);

BUFx3_ASAP7_75t_L g2548 ( 
.A(n_2439),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2385),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2421),
.A2(n_1512),
.B(n_1511),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2339),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2367),
.A2(n_1505),
.B1(n_1506),
.B2(n_1504),
.Y(n_2552)
);

INVx2_ASAP7_75t_SL g2553 ( 
.A(n_2326),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2342),
.B(n_1510),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2414),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2412),
.B(n_1513),
.Y(n_2556)
);

O2A1O1Ixp33_ASAP7_75t_L g2557 ( 
.A1(n_2368),
.A2(n_1519),
.B(n_1520),
.C(n_1515),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2394),
.B(n_1770),
.Y(n_2558)
);

AND2x6_ASAP7_75t_SL g2559 ( 
.A(n_2426),
.B(n_1521),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2432),
.B(n_1516),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2313),
.B(n_1517),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2450),
.B(n_1518),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2447),
.Y(n_2563)
);

INVxp67_ASAP7_75t_L g2564 ( 
.A(n_2419),
.Y(n_2564)
);

AO221x1_ASAP7_75t_L g2565 ( 
.A1(n_2347),
.A2(n_1537),
.B1(n_1541),
.B2(n_1536),
.C(n_1535),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2436),
.Y(n_2566)
);

A2O1A1Ixp33_ASAP7_75t_L g2567 ( 
.A1(n_2425),
.A2(n_1548),
.B(n_1550),
.C(n_1544),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2407),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2348),
.B(n_1523),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2375),
.B(n_1525),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2465),
.B(n_1526),
.Y(n_2571)
);

A2O1A1Ixp33_ASAP7_75t_L g2572 ( 
.A1(n_2410),
.A2(n_1574),
.B(n_1579),
.C(n_1568),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2389),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2430),
.B(n_1529),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2341),
.B(n_1530),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_R g2576 ( 
.A(n_2376),
.B(n_1532),
.Y(n_2576)
);

AOI22xp33_ASAP7_75t_L g2577 ( 
.A1(n_2365),
.A2(n_1593),
.B1(n_1594),
.B2(n_1588),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2323),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2405),
.B(n_2365),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2384),
.B(n_1540),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2332),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2397),
.B(n_1542),
.Y(n_2582)
);

INVx8_ASAP7_75t_L g2583 ( 
.A(n_2324),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2408),
.B(n_1543),
.Y(n_2584)
);

AOI22xp33_ASAP7_75t_L g2585 ( 
.A1(n_2384),
.A2(n_1600),
.B1(n_1609),
.B2(n_1599),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2336),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2315),
.A2(n_1546),
.B1(n_1547),
.B2(n_1545),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2363),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2353),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2422),
.B(n_1549),
.Y(n_2590)
);

AOI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2422),
.A2(n_1623),
.B1(n_1625),
.B2(n_1615),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_2344),
.B(n_1551),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2364),
.B(n_1799),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2366),
.B(n_1553),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2379),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2451),
.B(n_1554),
.Y(n_2596)
);

INVxp67_ASAP7_75t_SL g2597 ( 
.A(n_2381),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2350),
.B(n_1555),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2456),
.B(n_1799),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2452),
.Y(n_2600)
);

AOI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2460),
.A2(n_1558),
.B1(n_1559),
.B2(n_1556),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_L g2602 ( 
.A(n_2424),
.B(n_1563),
.Y(n_2602)
);

A2O1A1Ixp33_ASAP7_75t_L g2603 ( 
.A1(n_2361),
.A2(n_1640),
.B(n_1644),
.C(n_1638),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2396),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2350),
.B(n_1565),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2346),
.A2(n_1664),
.B1(n_1665),
.B2(n_1661),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_L g2607 ( 
.A(n_2458),
.B(n_1566),
.Y(n_2607)
);

AOI221xp5_ASAP7_75t_L g2608 ( 
.A1(n_2377),
.A2(n_1670),
.B1(n_1671),
.B2(n_1669),
.C(n_1667),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2346),
.B(n_1567),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2461),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2413),
.B(n_1570),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2428),
.B(n_1572),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2420),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2423),
.B(n_1573),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2429),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2427),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2395),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2431),
.Y(n_2618)
);

INVxp67_ASAP7_75t_L g2619 ( 
.A(n_2434),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2433),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2352),
.Y(n_2621)
);

OAI221xp5_ASAP7_75t_L g2622 ( 
.A1(n_2411),
.A2(n_1688),
.B1(n_1689),
.B2(n_1686),
.C(n_1672),
.Y(n_2622)
);

NOR3xp33_ASAP7_75t_L g2623 ( 
.A(n_2362),
.B(n_1576),
.C(n_1575),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2329),
.B(n_1856),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2318),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2333),
.B(n_1578),
.Y(n_2626)
);

OAI22xp5_ASAP7_75t_SL g2627 ( 
.A1(n_2362),
.A2(n_1581),
.B1(n_1582),
.B2(n_1580),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2333),
.B(n_1584),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2333),
.B(n_1585),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2318),
.Y(n_2630)
);

INVxp67_ASAP7_75t_L g2631 ( 
.A(n_2459),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2318),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2333),
.B(n_1586),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2445),
.Y(n_2634)
);

OR2x6_ASAP7_75t_L g2635 ( 
.A(n_2330),
.B(n_1691),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2333),
.B(n_1589),
.Y(n_2636)
);

INVx5_ASAP7_75t_L g2637 ( 
.A(n_2417),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2333),
.B(n_1590),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2333),
.B(n_1591),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2356),
.B(n_1592),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2333),
.B(n_1595),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2333),
.B(n_1596),
.Y(n_2642)
);

O2A1O1Ixp5_ASAP7_75t_L g2643 ( 
.A1(n_2333),
.A2(n_1694),
.B(n_1707),
.C(n_1692),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2333),
.B(n_1597),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2349),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2333),
.B(n_1598),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2333),
.B(n_1604),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2316),
.A2(n_1714),
.B1(n_1720),
.B2(n_1711),
.Y(n_2648)
);

OR2x6_ASAP7_75t_L g2649 ( 
.A(n_2330),
.B(n_1726),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2356),
.B(n_1607),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2333),
.B(n_1608),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_2380),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2333),
.B(n_1610),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2333),
.A2(n_1613),
.B1(n_1617),
.B2(n_1611),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2333),
.B(n_1618),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2469),
.Y(n_2656)
);

BUFx2_ASAP7_75t_L g2657 ( 
.A(n_2634),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2495),
.B(n_1622),
.Y(n_2658)
);

INVx4_ASAP7_75t_L g2659 ( 
.A(n_2479),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2470),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2551),
.B(n_1624),
.Y(n_2661)
);

AOI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2530),
.A2(n_1746),
.B(n_1745),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2507),
.A2(n_1627),
.B1(n_1628),
.B2(n_1626),
.Y(n_2663)
);

BUFx6f_ASAP7_75t_L g2664 ( 
.A(n_2505),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2508),
.B(n_1629),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2474),
.B(n_1631),
.Y(n_2666)
);

INVxp67_ASAP7_75t_L g2667 ( 
.A(n_2480),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2624),
.B(n_1856),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2505),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2475),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2626),
.B(n_1633),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2488),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2629),
.B(n_1635),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2531),
.A2(n_2556),
.B(n_2472),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2640),
.B(n_1636),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2633),
.B(n_1637),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2494),
.Y(n_2677)
);

AOI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2513),
.A2(n_1811),
.B(n_1803),
.Y(n_2678)
);

AOI21xp33_ASAP7_75t_L g2679 ( 
.A1(n_2650),
.A2(n_1641),
.B(n_1639),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2628),
.A2(n_1823),
.B(n_1821),
.Y(n_2680)
);

AOI21xp5_ASAP7_75t_L g2681 ( 
.A1(n_2636),
.A2(n_1831),
.B(n_1825),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2496),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2638),
.A2(n_1834),
.B(n_1832),
.Y(n_2683)
);

O2A1O1Ixp33_ASAP7_75t_L g2684 ( 
.A1(n_2468),
.A2(n_1839),
.B(n_1842),
.C(n_1838),
.Y(n_2684)
);

BUFx6f_ASAP7_75t_L g2685 ( 
.A(n_2613),
.Y(n_2685)
);

AOI21xp5_ASAP7_75t_L g2686 ( 
.A1(n_2641),
.A2(n_1846),
.B(n_1843),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2473),
.B(n_1642),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2479),
.B(n_1848),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2631),
.B(n_1643),
.Y(n_2689)
);

AO21x1_ASAP7_75t_L g2690 ( 
.A1(n_2503),
.A2(n_1852),
.B(n_1849),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2504),
.Y(n_2691)
);

BUFx2_ASAP7_75t_L g2692 ( 
.A(n_2540),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2639),
.B(n_1645),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2515),
.A2(n_1647),
.B1(n_1648),
.B2(n_1646),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2512),
.B(n_1871),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2489),
.Y(n_2696)
);

INVx3_ASAP7_75t_L g2697 ( 
.A(n_2613),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2493),
.Y(n_2698)
);

OR2x6_ASAP7_75t_L g2699 ( 
.A(n_2583),
.B(n_1864),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2498),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2544),
.B(n_1649),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2642),
.B(n_1651),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2653),
.A2(n_1873),
.B(n_1870),
.Y(n_2703)
);

O2A1O1Ixp5_ASAP7_75t_L g2704 ( 
.A1(n_2643),
.A2(n_1874),
.B(n_1879),
.C(n_1875),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2644),
.B(n_1654),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2625),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2637),
.B(n_1882),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2646),
.B(n_1656),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2630),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2655),
.A2(n_1887),
.B(n_1883),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2647),
.B(n_1658),
.Y(n_2711)
);

OAI21xp33_ASAP7_75t_SL g2712 ( 
.A1(n_2632),
.A2(n_1905),
.B(n_1898),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2490),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2651),
.B(n_1659),
.Y(n_2714)
);

NOR2x2_ASAP7_75t_L g2715 ( 
.A(n_2485),
.B(n_1871),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2490),
.Y(n_2716)
);

BUFx4f_ASAP7_75t_L g2717 ( 
.A(n_2566),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2471),
.B(n_1660),
.Y(n_2718)
);

O2A1O1Ixp33_ASAP7_75t_SL g2719 ( 
.A1(n_2521),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2510),
.A2(n_1663),
.B(n_1662),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2491),
.B(n_1886),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2514),
.A2(n_1676),
.B(n_1674),
.Y(n_2722)
);

AOI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2517),
.A2(n_1679),
.B(n_1677),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2501),
.B(n_1680),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2502),
.B(n_1681),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2523),
.A2(n_1697),
.B(n_1696),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2532),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2555),
.Y(n_2728)
);

OR2x2_ASAP7_75t_L g2729 ( 
.A(n_2478),
.B(n_1700),
.Y(n_2729)
);

AOI21x1_ASAP7_75t_L g2730 ( 
.A1(n_2516),
.A2(n_242),
.B(n_241),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_SL g2731 ( 
.A(n_2652),
.B(n_2547),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2554),
.B(n_1712),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2529),
.B(n_1713),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2549),
.Y(n_2734)
);

OAI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2506),
.A2(n_1716),
.B(n_1715),
.Y(n_2735)
);

AOI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2482),
.A2(n_1719),
.B1(n_1724),
.B2(n_1718),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2597),
.A2(n_1730),
.B(n_1729),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2518),
.A2(n_1734),
.B(n_1733),
.Y(n_2738)
);

OR2x6_ASAP7_75t_L g2739 ( 
.A(n_2583),
.B(n_1886),
.Y(n_2739)
);

A2O1A1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_2623),
.A2(n_1737),
.B(n_1739),
.C(n_1736),
.Y(n_2740)
);

AOI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2525),
.A2(n_1742),
.B(n_1741),
.Y(n_2741)
);

O2A1O1Ixp33_ASAP7_75t_L g2742 ( 
.A1(n_2557),
.A2(n_1900),
.B(n_1915),
.C(n_1890),
.Y(n_2742)
);

OAI321xp33_ASAP7_75t_L g2743 ( 
.A1(n_2627),
.A2(n_1900),
.A3(n_1915),
.B1(n_1890),
.B2(n_1753),
.C(n_1751),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2539),
.B(n_1750),
.Y(n_2744)
);

INVx11_ASAP7_75t_L g2745 ( 
.A(n_2620),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2645),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2564),
.B(n_1755),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2533),
.A2(n_1757),
.B(n_1756),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2604),
.B(n_1758),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2526),
.Y(n_2750)
);

OR2x6_ASAP7_75t_L g2751 ( 
.A(n_2617),
.B(n_241),
.Y(n_2751)
);

AOI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2534),
.A2(n_1763),
.B(n_1761),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2621),
.Y(n_2753)
);

INVx4_ASAP7_75t_L g2754 ( 
.A(n_2548),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2527),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2563),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_SL g2757 ( 
.A(n_2500),
.B(n_1764),
.Y(n_2757)
);

AOI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2535),
.A2(n_1766),
.B(n_1765),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2536),
.Y(n_2759)
);

AND2x4_ASAP7_75t_L g2760 ( 
.A(n_2615),
.B(n_1771),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2492),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2558),
.B(n_1774),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2545),
.B(n_2574),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2499),
.A2(n_2570),
.B(n_2509),
.Y(n_2764)
);

AOI21xp5_ASAP7_75t_L g2765 ( 
.A1(n_2594),
.A2(n_1782),
.B(n_1781),
.Y(n_2765)
);

OAI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2476),
.A2(n_1788),
.B(n_1787),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2561),
.A2(n_1793),
.B(n_1792),
.Y(n_2767)
);

AOI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2562),
.A2(n_1796),
.B(n_1795),
.Y(n_2768)
);

NOR2xp67_ASAP7_75t_L g2769 ( 
.A(n_2596),
.B(n_1797),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2477),
.A2(n_1802),
.B(n_1801),
.Y(n_2770)
);

NOR2xp67_ASAP7_75t_L g2771 ( 
.A(n_2607),
.B(n_1805),
.Y(n_2771)
);

AOI21xp5_ASAP7_75t_L g2772 ( 
.A1(n_2481),
.A2(n_1809),
.B(n_1806),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2483),
.A2(n_1813),
.B(n_1810),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2484),
.A2(n_1819),
.B(n_1816),
.Y(n_2774)
);

O2A1O1Ixp33_ASAP7_75t_L g2775 ( 
.A1(n_2567),
.A2(n_1822),
.B(n_1824),
.C(n_1820),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2578),
.Y(n_2776)
);

AOI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2538),
.A2(n_1828),
.B(n_1827),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2541),
.A2(n_1837),
.B(n_1835),
.Y(n_2778)
);

NOR2x1p5_ASAP7_75t_SL g2779 ( 
.A(n_2581),
.B(n_1850),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2584),
.B(n_1851),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2595),
.Y(n_2781)
);

AOI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2543),
.A2(n_1855),
.B(n_1854),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2654),
.B(n_2648),
.Y(n_2783)
);

BUFx6f_ASAP7_75t_L g2784 ( 
.A(n_2519),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2579),
.B(n_1859),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2582),
.B(n_1860),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2511),
.B(n_1878),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2550),
.B(n_2560),
.Y(n_2788)
);

O2A1O1Ixp33_ASAP7_75t_L g2789 ( 
.A1(n_2572),
.A2(n_1885),
.B(n_1889),
.C(n_1884),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2593),
.B(n_2599),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2528),
.A2(n_2614),
.B(n_2588),
.Y(n_2791)
);

INVxp67_ASAP7_75t_L g2792 ( 
.A(n_2616),
.Y(n_2792)
);

BUFx12f_ASAP7_75t_L g2793 ( 
.A(n_2559),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2591),
.B(n_1892),
.Y(n_2794)
);

AOI21xp5_ASAP7_75t_L g2795 ( 
.A1(n_2586),
.A2(n_1895),
.B(n_1893),
.Y(n_2795)
);

AOI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2553),
.A2(n_1897),
.B(n_1896),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2568),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2577),
.B(n_1904),
.Y(n_2798)
);

AOI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2573),
.A2(n_2575),
.B(n_2589),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2487),
.Y(n_2800)
);

AOI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2542),
.A2(n_1907),
.B(n_1906),
.Y(n_2801)
);

A2O1A1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2618),
.A2(n_1913),
.B(n_1914),
.C(n_1912),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2585),
.B(n_1918),
.Y(n_2803)
);

INVx3_ASAP7_75t_SL g2804 ( 
.A(n_2664),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2763),
.B(n_2576),
.Y(n_2805)
);

INVx4_ASAP7_75t_L g2806 ( 
.A(n_2685),
.Y(n_2806)
);

INVx3_ASAP7_75t_L g2807 ( 
.A(n_2659),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2675),
.B(n_2520),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2656),
.Y(n_2809)
);

NAND3xp33_ASAP7_75t_L g2810 ( 
.A(n_2658),
.B(n_2608),
.C(n_2486),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2764),
.A2(n_2580),
.B(n_2598),
.Y(n_2811)
);

AOI21xp5_ASAP7_75t_L g2812 ( 
.A1(n_2674),
.A2(n_2605),
.B(n_2592),
.Y(n_2812)
);

BUFx2_ASAP7_75t_L g2813 ( 
.A(n_2660),
.Y(n_2813)
);

A2O1A1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2666),
.A2(n_2590),
.B(n_2611),
.C(n_2569),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_2745),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_SL g2816 ( 
.A(n_2731),
.B(n_2610),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2687),
.B(n_2524),
.Y(n_2817)
);

HB1xp67_ASAP7_75t_SL g2818 ( 
.A(n_2685),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2668),
.B(n_2721),
.Y(n_2819)
);

BUFx2_ASAP7_75t_L g2820 ( 
.A(n_2657),
.Y(n_2820)
);

AOI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2788),
.A2(n_2791),
.B(n_2671),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2762),
.B(n_2565),
.Y(n_2822)
);

OAI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2783),
.A2(n_2600),
.B1(n_2612),
.B2(n_2606),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2786),
.B(n_2522),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2713),
.Y(n_2825)
);

AOI21xp5_ASAP7_75t_L g2826 ( 
.A1(n_2673),
.A2(n_2602),
.B(n_2571),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2676),
.A2(n_2609),
.B(n_2603),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2672),
.Y(n_2828)
);

INVxp67_ASAP7_75t_L g2829 ( 
.A(n_2692),
.Y(n_2829)
);

NAND3xp33_ASAP7_75t_SL g2830 ( 
.A(n_2780),
.B(n_2601),
.C(n_2587),
.Y(n_2830)
);

A2O1A1Ixp33_ASAP7_75t_L g2831 ( 
.A1(n_2718),
.A2(n_2546),
.B(n_2622),
.C(n_2552),
.Y(n_2831)
);

OAI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2677),
.A2(n_2497),
.B1(n_2619),
.B2(n_2635),
.Y(n_2832)
);

INVx1_ASAP7_75t_SL g2833 ( 
.A(n_2756),
.Y(n_2833)
);

NOR2x1_ASAP7_75t_L g2834 ( 
.A(n_2754),
.B(n_2649),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2733),
.B(n_2537),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2693),
.A2(n_1924),
.B(n_1923),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2682),
.Y(n_2837)
);

BUFx3_ASAP7_75t_L g2838 ( 
.A(n_2717),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2691),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2702),
.A2(n_1929),
.B(n_1927),
.Y(n_2840)
);

AOI21x1_ASAP7_75t_L g2841 ( 
.A1(n_2785),
.A2(n_246),
.B(n_245),
.Y(n_2841)
);

O2A1O1Ixp33_ASAP7_75t_L g2842 ( 
.A1(n_2679),
.A2(n_247),
.B(n_248),
.C(n_246),
.Y(n_2842)
);

OR2x6_ASAP7_75t_L g2843 ( 
.A(n_2664),
.B(n_247),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2705),
.A2(n_249),
.B(n_248),
.Y(n_2844)
);

CKINVDCx11_ASAP7_75t_R g2845 ( 
.A(n_2793),
.Y(n_2845)
);

AOI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2708),
.A2(n_251),
.B(n_250),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2711),
.B(n_2),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2714),
.B(n_2667),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2724),
.B(n_252),
.Y(n_2849)
);

AOI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2725),
.A2(n_254),
.B(n_252),
.Y(n_2850)
);

AOI21x1_ASAP7_75t_L g2851 ( 
.A1(n_2662),
.A2(n_256),
.B(n_254),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2790),
.A2(n_257),
.B1(n_258),
.B2(n_256),
.Y(n_2852)
);

INVx1_ASAP7_75t_SL g2853 ( 
.A(n_2716),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2706),
.A2(n_258),
.B1(n_259),
.B2(n_257),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2661),
.B(n_2),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2695),
.B(n_259),
.Y(n_2856)
);

BUFx12f_ASAP7_75t_L g2857 ( 
.A(n_2669),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2709),
.Y(n_2858)
);

NAND3xp33_ASAP7_75t_SL g2859 ( 
.A(n_2742),
.B(n_4),
.C(n_5),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_2716),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2732),
.A2(n_261),
.B(n_260),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2744),
.B(n_262),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2669),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2727),
.A2(n_263),
.B1(n_264),
.B2(n_262),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2728),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2799),
.A2(n_264),
.B(n_263),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2769),
.B(n_7),
.Y(n_2867)
);

OAI22x1_ASAP7_75t_L g2868 ( 
.A1(n_2736),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2868)
);

AOI22xp33_ASAP7_75t_SL g2869 ( 
.A1(n_2787),
.A2(n_267),
.B1(n_268),
.B2(n_265),
.Y(n_2869)
);

AOI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2665),
.A2(n_269),
.B(n_267),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2771),
.B(n_8),
.Y(n_2871)
);

O2A1O1Ixp33_ASAP7_75t_L g2872 ( 
.A1(n_2701),
.A2(n_270),
.B(n_271),
.C(n_269),
.Y(n_2872)
);

NOR3xp33_ASAP7_75t_L g2873 ( 
.A(n_2743),
.B(n_9),
.C(n_10),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2734),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2753),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_R g2876 ( 
.A(n_2697),
.B(n_272),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2750),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2755),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2759),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_SL g2880 ( 
.A(n_2792),
.B(n_273),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2753),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2761),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_2797),
.B(n_279),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2670),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2747),
.B(n_280),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2784),
.Y(n_2886)
);

OAI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2704),
.A2(n_12),
.B(n_13),
.Y(n_2887)
);

BUFx6f_ASAP7_75t_L g2888 ( 
.A(n_2784),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2735),
.B(n_13),
.Y(n_2889)
);

BUFx2_ASAP7_75t_SL g2890 ( 
.A(n_2800),
.Y(n_2890)
);

AO21x1_ASAP7_75t_L g2891 ( 
.A1(n_2730),
.A2(n_283),
.B(n_282),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_R g2892 ( 
.A(n_2757),
.B(n_283),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_SL g2893 ( 
.A(n_2689),
.B(n_284),
.Y(n_2893)
);

NOR3xp33_ASAP7_75t_SL g2894 ( 
.A(n_2740),
.B(n_13),
.C(n_14),
.Y(n_2894)
);

OAI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2802),
.A2(n_14),
.B(n_15),
.Y(n_2895)
);

INVx3_ASAP7_75t_SL g2896 ( 
.A(n_2760),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2696),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2698),
.A2(n_288),
.B1(n_289),
.B2(n_287),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2700),
.A2(n_292),
.B1(n_293),
.B2(n_291),
.Y(n_2899)
);

BUFx8_ASAP7_75t_L g2900 ( 
.A(n_2688),
.Y(n_2900)
);

OR2x6_ASAP7_75t_L g2901 ( 
.A(n_2699),
.B(n_294),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2746),
.Y(n_2902)
);

OR2x6_ASAP7_75t_L g2903 ( 
.A(n_2739),
.B(n_295),
.Y(n_2903)
);

INVx2_ASAP7_75t_SL g2904 ( 
.A(n_2707),
.Y(n_2904)
);

A2O1A1Ixp33_ASAP7_75t_L g2905 ( 
.A1(n_2775),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_2905)
);

AND2x4_ASAP7_75t_L g2906 ( 
.A(n_2776),
.B(n_2779),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2781),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2729),
.B(n_296),
.Y(n_2908)
);

OR2x6_ASAP7_75t_L g2909 ( 
.A(n_2751),
.B(n_297),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2712),
.Y(n_2910)
);

AO21x1_ASAP7_75t_L g2911 ( 
.A1(n_2789),
.A2(n_299),
.B(n_298),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2719),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_R g2913 ( 
.A(n_2794),
.B(n_298),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2798),
.Y(n_2914)
);

BUFx6f_ASAP7_75t_L g2915 ( 
.A(n_2749),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2694),
.A2(n_300),
.B1(n_302),
.B2(n_299),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2766),
.B(n_305),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2795),
.A2(n_307),
.B(n_306),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2748),
.B(n_308),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2663),
.B(n_308),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_R g2921 ( 
.A(n_2803),
.B(n_310),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2752),
.A2(n_312),
.B(n_311),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2678),
.B(n_20),
.Y(n_2923)
);

AOI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2758),
.A2(n_313),
.B(n_312),
.Y(n_2924)
);

CKINVDCx12_ASAP7_75t_R g2925 ( 
.A(n_2715),
.Y(n_2925)
);

HB1xp67_ASAP7_75t_L g2926 ( 
.A(n_2690),
.Y(n_2926)
);

NAND2x1p5_ASAP7_75t_L g2927 ( 
.A(n_2778),
.B(n_314),
.Y(n_2927)
);

AOI221xp5_ASAP7_75t_L g2928 ( 
.A1(n_2684),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2680),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2681),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2782),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2770),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2683),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2686),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2737),
.B(n_316),
.Y(n_2935)
);

NOR2x1_ASAP7_75t_L g2936 ( 
.A(n_2796),
.B(n_316),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2772),
.B(n_24),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2773),
.B(n_25),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2703),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2710),
.Y(n_2940)
);

INVxp67_ASAP7_75t_L g2941 ( 
.A(n_2801),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2767),
.B(n_2768),
.Y(n_2942)
);

OAI21xp33_ASAP7_75t_L g2943 ( 
.A1(n_2774),
.A2(n_25),
.B(n_26),
.Y(n_2943)
);

A2O1A1Ixp33_ASAP7_75t_SL g2944 ( 
.A1(n_2765),
.A2(n_2720),
.B(n_2723),
.C(n_2722),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2738),
.Y(n_2945)
);

NAND2x1p5_ASAP7_75t_L g2946 ( 
.A(n_2741),
.B(n_320),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2726),
.A2(n_322),
.B(n_321),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2777),
.B(n_27),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2656),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2764),
.A2(n_325),
.B(n_324),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_R g2951 ( 
.A(n_2731),
.B(n_324),
.Y(n_2951)
);

OAI21x1_ASAP7_75t_L g2952 ( 
.A1(n_2674),
.A2(n_29),
.B(n_30),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2656),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2717),
.Y(n_2954)
);

INVx3_ASAP7_75t_SL g2955 ( 
.A(n_2664),
.Y(n_2955)
);

NOR3xp33_ASAP7_75t_SL g2956 ( 
.A(n_2743),
.B(n_30),
.C(n_31),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2763),
.B(n_31),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2764),
.A2(n_328),
.B(n_326),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_2675),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2959)
);

INVx2_ASAP7_75t_SL g2960 ( 
.A(n_2717),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2763),
.B(n_32),
.Y(n_2961)
);

OAI21x1_ASAP7_75t_L g2962 ( 
.A1(n_2821),
.A2(n_33),
.B(n_34),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2809),
.Y(n_2963)
);

O2A1O1Ixp33_ASAP7_75t_SL g2964 ( 
.A1(n_2831),
.A2(n_331),
.B(n_332),
.C(n_330),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2838),
.Y(n_2965)
);

INVxp67_ASAP7_75t_SL g2966 ( 
.A(n_2820),
.Y(n_2966)
);

AO31x2_ASAP7_75t_L g2967 ( 
.A1(n_2891),
.A2(n_39),
.A3(n_36),
.B(n_38),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2808),
.B(n_2848),
.Y(n_2968)
);

OAI21x1_ASAP7_75t_L g2969 ( 
.A1(n_2952),
.A2(n_2812),
.B(n_2811),
.Y(n_2969)
);

OAI21x1_ASAP7_75t_L g2970 ( 
.A1(n_2942),
.A2(n_39),
.B(n_40),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_L g2971 ( 
.A1(n_2910),
.A2(n_40),
.B(n_41),
.Y(n_2971)
);

OAI21xp5_ASAP7_75t_L g2972 ( 
.A1(n_2810),
.A2(n_40),
.B(n_42),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2858),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2805),
.B(n_2817),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2824),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_2975)
);

INVxp67_ASAP7_75t_SL g2976 ( 
.A(n_2829),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2882),
.B(n_2954),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2949),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2835),
.B(n_333),
.Y(n_2979)
);

OAI21x1_ASAP7_75t_SL g2980 ( 
.A1(n_2895),
.A2(n_46),
.B(n_47),
.Y(n_2980)
);

AOI21xp5_ASAP7_75t_L g2981 ( 
.A1(n_2814),
.A2(n_334),
.B(n_333),
.Y(n_2981)
);

BUFx3_ASAP7_75t_L g2982 ( 
.A(n_2857),
.Y(n_2982)
);

BUFx6f_ASAP7_75t_SL g2983 ( 
.A(n_2960),
.Y(n_2983)
);

AO21x1_ASAP7_75t_L g2984 ( 
.A1(n_2889),
.A2(n_336),
.B(n_335),
.Y(n_2984)
);

BUFx12f_ASAP7_75t_L g2985 ( 
.A(n_2815),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2828),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2837),
.Y(n_2987)
);

OAI21x1_ASAP7_75t_L g2988 ( 
.A1(n_2945),
.A2(n_49),
.B(n_50),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2839),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2914),
.B(n_2957),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2961),
.B(n_50),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2819),
.B(n_50),
.Y(n_2992)
);

AND2x4_ASAP7_75t_L g2993 ( 
.A(n_2863),
.B(n_337),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2860),
.B(n_337),
.Y(n_2994)
);

AOI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2944),
.A2(n_2826),
.B(n_2827),
.Y(n_2995)
);

AOI21x1_ASAP7_75t_L g2996 ( 
.A1(n_2926),
.A2(n_51),
.B(n_52),
.Y(n_2996)
);

NAND3xp33_ASAP7_75t_L g2997 ( 
.A(n_2920),
.B(n_53),
.C(n_54),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2862),
.B(n_54),
.Y(n_2998)
);

O2A1O1Ixp5_ASAP7_75t_L g2999 ( 
.A1(n_2919),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2849),
.B(n_55),
.Y(n_3000)
);

AOI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2941),
.A2(n_340),
.B(n_339),
.Y(n_3001)
);

OAI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2816),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2950),
.A2(n_57),
.B(n_58),
.Y(n_3003)
);

BUFx6f_ASAP7_75t_L g3004 ( 
.A(n_2825),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2877),
.Y(n_3005)
);

AOI21xp5_ASAP7_75t_L g3006 ( 
.A1(n_2830),
.A2(n_342),
.B(n_341),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2856),
.B(n_60),
.Y(n_3007)
);

NOR2xp67_ASAP7_75t_L g3008 ( 
.A(n_2807),
.B(n_61),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2847),
.B(n_62),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2855),
.B(n_62),
.Y(n_3010)
);

O2A1O1Ixp33_ASAP7_75t_L g3011 ( 
.A1(n_2893),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_3011)
);

OA21x2_ASAP7_75t_L g3012 ( 
.A1(n_2887),
.A2(n_64),
.B(n_65),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2917),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_3013)
);

OAI21x1_ASAP7_75t_SL g3014 ( 
.A1(n_2911),
.A2(n_66),
.B(n_67),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2823),
.B(n_67),
.Y(n_3015)
);

AO21x1_ASAP7_75t_L g3016 ( 
.A1(n_2958),
.A2(n_345),
.B(n_344),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2934),
.A2(n_346),
.B(n_345),
.Y(n_3017)
);

AO31x2_ASAP7_75t_L g3018 ( 
.A1(n_2912),
.A2(n_71),
.A3(n_68),
.B(n_69),
.Y(n_3018)
);

AOI21xp5_ASAP7_75t_L g3019 ( 
.A1(n_2939),
.A2(n_347),
.B(n_346),
.Y(n_3019)
);

INVx5_ASAP7_75t_L g3020 ( 
.A(n_2825),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2865),
.Y(n_3021)
);

AOI21xp33_ASAP7_75t_L g3022 ( 
.A1(n_2937),
.A2(n_72),
.B(n_73),
.Y(n_3022)
);

INVx3_ASAP7_75t_L g3023 ( 
.A(n_2886),
.Y(n_3023)
);

CKINVDCx11_ASAP7_75t_R g3024 ( 
.A(n_2845),
.Y(n_3024)
);

OAI21x1_ASAP7_75t_L g3025 ( 
.A1(n_2866),
.A2(n_73),
.B(n_74),
.Y(n_3025)
);

BUFx10_ASAP7_75t_L g3026 ( 
.A(n_2886),
.Y(n_3026)
);

NAND2xp33_ASAP7_75t_R g3027 ( 
.A(n_2951),
.B(n_348),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2813),
.B(n_349),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2929),
.A2(n_352),
.B(n_350),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2874),
.Y(n_3030)
);

NAND3xp33_ASAP7_75t_L g3031 ( 
.A(n_2873),
.B(n_75),
.C(n_76),
.Y(n_3031)
);

INVx1_ASAP7_75t_SL g3032 ( 
.A(n_2818),
.Y(n_3032)
);

INVx1_ASAP7_75t_SL g3033 ( 
.A(n_2833),
.Y(n_3033)
);

OAI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2836),
.A2(n_77),
.B(n_78),
.Y(n_3034)
);

O2A1O1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2885),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2953),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2907),
.Y(n_3037)
);

AOI221xp5_ASAP7_75t_L g3038 ( 
.A1(n_2859),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.C(n_82),
.Y(n_3038)
);

OAI21xp5_ASAP7_75t_L g3039 ( 
.A1(n_2840),
.A2(n_81),
.B(n_82),
.Y(n_3039)
);

CKINVDCx5p33_ASAP7_75t_R g3040 ( 
.A(n_2890),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2878),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2884),
.Y(n_3042)
);

OAI21x1_ASAP7_75t_SL g3043 ( 
.A1(n_2851),
.A2(n_83),
.B(n_84),
.Y(n_3043)
);

OAI21x1_ASAP7_75t_L g3044 ( 
.A1(n_2930),
.A2(n_83),
.B(n_84),
.Y(n_3044)
);

HB1xp67_ASAP7_75t_L g3045 ( 
.A(n_2881),
.Y(n_3045)
);

OR2x6_ASAP7_75t_L g3046 ( 
.A(n_2888),
.B(n_2806),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_SL g3047 ( 
.A(n_2915),
.B(n_353),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2879),
.Y(n_3048)
);

CKINVDCx9p33_ASAP7_75t_R g3049 ( 
.A(n_2875),
.Y(n_3049)
);

INVxp67_ASAP7_75t_L g3050 ( 
.A(n_2888),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2933),
.A2(n_355),
.B(n_354),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2908),
.B(n_354),
.Y(n_3052)
);

NOR2x1_ASAP7_75t_L g3053 ( 
.A(n_2834),
.B(n_355),
.Y(n_3053)
);

AO32x2_ASAP7_75t_L g3054 ( 
.A1(n_2916),
.A2(n_87),
.A3(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2940),
.A2(n_357),
.B(n_356),
.Y(n_3055)
);

NOR2xp67_ASAP7_75t_L g3056 ( 
.A(n_2902),
.B(n_88),
.Y(n_3056)
);

OAI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_2956),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3057)
);

AOI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2931),
.A2(n_359),
.B(n_358),
.Y(n_3058)
);

OAI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2947),
.A2(n_89),
.B(n_91),
.Y(n_3059)
);

OR2x6_ASAP7_75t_L g3060 ( 
.A(n_2904),
.B(n_360),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_SL g3061 ( 
.A1(n_2905),
.A2(n_361),
.B(n_360),
.Y(n_3061)
);

OAI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2938),
.A2(n_96),
.B(n_97),
.Y(n_3062)
);

HB1xp67_ASAP7_75t_L g3063 ( 
.A(n_2853),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2915),
.B(n_364),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_2943),
.A2(n_2948),
.B(n_2924),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2822),
.B(n_98),
.Y(n_3066)
);

OR2x2_ASAP7_75t_L g3067 ( 
.A(n_2897),
.B(n_364),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2841),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2922),
.A2(n_366),
.B(n_365),
.Y(n_3069)
);

OAI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2870),
.A2(n_101),
.B(n_102),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2959),
.B(n_103),
.Y(n_3071)
);

OAI21x1_ASAP7_75t_L g3072 ( 
.A1(n_2918),
.A2(n_104),
.B(n_105),
.Y(n_3072)
);

AOI21xp5_ASAP7_75t_SL g3073 ( 
.A1(n_2906),
.A2(n_368),
.B(n_367),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2883),
.B(n_104),
.Y(n_3074)
);

AO31x2_ASAP7_75t_L g3075 ( 
.A1(n_2868),
.A2(n_107),
.A3(n_105),
.B(n_106),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2880),
.B(n_106),
.Y(n_3076)
);

OAI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_2832),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3077)
);

OA21x2_ASAP7_75t_L g3078 ( 
.A1(n_2867),
.A2(n_109),
.B(n_110),
.Y(n_3078)
);

AO31x2_ASAP7_75t_L g3079 ( 
.A1(n_2844),
.A2(n_2850),
.A3(n_2861),
.B(n_2846),
.Y(n_3079)
);

BUFx6f_ASAP7_75t_L g3080 ( 
.A(n_2804),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_2955),
.Y(n_3081)
);

AO31x2_ASAP7_75t_L g3082 ( 
.A1(n_2871),
.A2(n_114),
.A3(n_112),
.B(n_113),
.Y(n_3082)
);

OAI21x1_ASAP7_75t_SL g3083 ( 
.A1(n_2872),
.A2(n_112),
.B(n_114),
.Y(n_3083)
);

INVx5_ASAP7_75t_L g3084 ( 
.A(n_2843),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_SL g3085 ( 
.A1(n_2842),
.A2(n_369),
.B(n_368),
.Y(n_3085)
);

BUFx6f_ASAP7_75t_L g3086 ( 
.A(n_2896),
.Y(n_3086)
);

OAI21x1_ASAP7_75t_L g3087 ( 
.A1(n_2936),
.A2(n_115),
.B(n_116),
.Y(n_3087)
);

INVx4_ASAP7_75t_L g3088 ( 
.A(n_2843),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2894),
.B(n_2935),
.Y(n_3089)
);

OAI21x1_ASAP7_75t_L g3090 ( 
.A1(n_2969),
.A2(n_2946),
.B(n_2927),
.Y(n_3090)
);

OAI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2981),
.A2(n_2923),
.B(n_2932),
.Y(n_3091)
);

OAI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_3065),
.A2(n_2928),
.B(n_2869),
.Y(n_3092)
);

OAI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_3027),
.A2(n_2852),
.B1(n_2901),
.B2(n_2909),
.Y(n_3093)
);

OAI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2995),
.A2(n_2899),
.B(n_2898),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_SL g3095 ( 
.A1(n_2972),
.A2(n_2892),
.B1(n_2921),
.B2(n_2913),
.Y(n_3095)
);

CKINVDCx20_ASAP7_75t_R g3096 ( 
.A(n_3024),
.Y(n_3096)
);

INVxp67_ASAP7_75t_SL g3097 ( 
.A(n_2966),
.Y(n_3097)
);

OAI21x1_ASAP7_75t_L g3098 ( 
.A1(n_2962),
.A2(n_2864),
.B(n_2854),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2986),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2978),
.Y(n_3100)
);

HB1xp67_ASAP7_75t_L g3101 ( 
.A(n_3045),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2987),
.Y(n_3102)
);

OAI33xp33_ASAP7_75t_L g3103 ( 
.A1(n_3057),
.A2(n_2925),
.A3(n_2876),
.B1(n_120),
.B2(n_122),
.B3(n_118),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2974),
.B(n_2901),
.Y(n_3104)
);

AO21x2_ASAP7_75t_L g3105 ( 
.A1(n_3043),
.A2(n_2903),
.B(n_2900),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2989),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3089),
.B(n_2903),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_3005),
.Y(n_3108)
);

OAI21x1_ASAP7_75t_L g3109 ( 
.A1(n_3044),
.A2(n_118),
.B(n_119),
.Y(n_3109)
);

HB1xp67_ASAP7_75t_L g3110 ( 
.A(n_3021),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_3030),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3036),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_3048),
.Y(n_3113)
);

NAND2xp33_ASAP7_75t_L g3114 ( 
.A(n_2968),
.B(n_121),
.Y(n_3114)
);

BUFx3_ASAP7_75t_L g3115 ( 
.A(n_2977),
.Y(n_3115)
);

OAI21x1_ASAP7_75t_L g3116 ( 
.A1(n_2988),
.A2(n_121),
.B(n_123),
.Y(n_3116)
);

AOI221xp5_ASAP7_75t_L g3117 ( 
.A1(n_2998),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_3117)
);

OA21x2_ASAP7_75t_L g3118 ( 
.A1(n_2970),
.A2(n_124),
.B(n_125),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_3086),
.Y(n_3119)
);

CKINVDCx20_ASAP7_75t_R g3120 ( 
.A(n_2985),
.Y(n_3120)
);

HB1xp67_ASAP7_75t_L g3121 ( 
.A(n_3037),
.Y(n_3121)
);

OAI21x1_ASAP7_75t_L g3122 ( 
.A1(n_3003),
.A2(n_124),
.B(n_126),
.Y(n_3122)
);

OA21x2_ASAP7_75t_L g3123 ( 
.A1(n_2971),
.A2(n_127),
.B(n_128),
.Y(n_3123)
);

AOI21x1_ASAP7_75t_L g3124 ( 
.A1(n_3015),
.A2(n_127),
.B(n_128),
.Y(n_3124)
);

BUFx2_ASAP7_75t_L g3125 ( 
.A(n_3049),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_3041),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3042),
.Y(n_3127)
);

OAI21x1_ASAP7_75t_L g3128 ( 
.A1(n_3025),
.A2(n_129),
.B(n_130),
.Y(n_3128)
);

OAI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_3059),
.A2(n_131),
.B(n_132),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2990),
.B(n_370),
.Y(n_3130)
);

INVxp67_ASAP7_75t_SL g3131 ( 
.A(n_2976),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2963),
.Y(n_3132)
);

AOI221xp5_ASAP7_75t_L g3133 ( 
.A1(n_3000),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_3133)
);

INVx3_ASAP7_75t_L g3134 ( 
.A(n_3026),
.Y(n_3134)
);

BUFx12f_ASAP7_75t_L g3135 ( 
.A(n_3080),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2973),
.Y(n_3136)
);

OAI21x1_ASAP7_75t_L g3137 ( 
.A1(n_3072),
.A2(n_136),
.B(n_137),
.Y(n_3137)
);

OA21x2_ASAP7_75t_L g3138 ( 
.A1(n_3068),
.A2(n_138),
.B(n_139),
.Y(n_3138)
);

BUFx4f_ASAP7_75t_L g3139 ( 
.A(n_3080),
.Y(n_3139)
);

OA21x2_ASAP7_75t_L g3140 ( 
.A1(n_3006),
.A2(n_140),
.B(n_141),
.Y(n_3140)
);

AO32x2_ASAP7_75t_L g3141 ( 
.A1(n_2975),
.A2(n_144),
.A3(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_3141)
);

OAI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2996),
.A2(n_142),
.B(n_143),
.Y(n_3142)
);

NOR2x1_ASAP7_75t_R g3143 ( 
.A(n_3084),
.B(n_3040),
.Y(n_3143)
);

OAI21x1_ASAP7_75t_L g3144 ( 
.A1(n_3069),
.A2(n_143),
.B(n_144),
.Y(n_3144)
);

INVx1_ASAP7_75t_SL g3145 ( 
.A(n_3033),
.Y(n_3145)
);

OAI22xp33_ASAP7_75t_L g3146 ( 
.A1(n_3013),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_3146)
);

NAND2x1p5_ASAP7_75t_L g3147 ( 
.A(n_3020),
.B(n_3084),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_2965),
.Y(n_3148)
);

BUFx8_ASAP7_75t_L g3149 ( 
.A(n_2983),
.Y(n_3149)
);

NAND3xp33_ASAP7_75t_L g3150 ( 
.A(n_3034),
.B(n_145),
.C(n_146),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_3029),
.A2(n_147),
.B(n_148),
.Y(n_3151)
);

OAI21x1_ASAP7_75t_L g3152 ( 
.A1(n_3051),
.A2(n_147),
.B(n_148),
.Y(n_3152)
);

INVx4_ASAP7_75t_L g3153 ( 
.A(n_3004),
.Y(n_3153)
);

INVx4_ASAP7_75t_SL g3154 ( 
.A(n_3018),
.Y(n_3154)
);

AND2x6_ASAP7_75t_L g3155 ( 
.A(n_3053),
.B(n_372),
.Y(n_3155)
);

AOI21xp33_ASAP7_75t_L g3156 ( 
.A1(n_3039),
.A2(n_149),
.B(n_150),
.Y(n_3156)
);

CKINVDCx11_ASAP7_75t_R g3157 ( 
.A(n_3032),
.Y(n_3157)
);

CKINVDCx6p67_ASAP7_75t_R g3158 ( 
.A(n_2982),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2967),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_3067),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2964),
.A2(n_375),
.B(n_374),
.Y(n_3161)
);

OAI21x1_ASAP7_75t_L g3162 ( 
.A1(n_3055),
.A2(n_152),
.B(n_153),
.Y(n_3162)
);

BUFx2_ASAP7_75t_SL g3163 ( 
.A(n_3081),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_3070),
.A2(n_152),
.B(n_153),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3062),
.B(n_376),
.Y(n_3165)
);

OAI21x1_ASAP7_75t_L g3166 ( 
.A1(n_3087),
.A2(n_154),
.B(n_155),
.Y(n_3166)
);

OR2x6_ASAP7_75t_L g3167 ( 
.A(n_3073),
.B(n_377),
.Y(n_3167)
);

HB1xp67_ASAP7_75t_L g3168 ( 
.A(n_3063),
.Y(n_3168)
);

AOI22xp33_ASAP7_75t_L g3169 ( 
.A1(n_2997),
.A2(n_3031),
.B1(n_3038),
.B2(n_3052),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2991),
.B(n_377),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3082),
.Y(n_3171)
);

AO21x2_ASAP7_75t_L g3172 ( 
.A1(n_3014),
.A2(n_2980),
.B(n_3016),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_3088),
.B(n_379),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_3079),
.Y(n_3174)
);

INVx1_ASAP7_75t_SL g3175 ( 
.A(n_3023),
.Y(n_3175)
);

OAI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_2979),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_3022),
.A2(n_2984),
.B1(n_3071),
.B2(n_3002),
.Y(n_3177)
);

AO21x2_ASAP7_75t_L g3178 ( 
.A1(n_3083),
.A2(n_157),
.B(n_158),
.Y(n_3178)
);

OAI21x1_ASAP7_75t_L g3179 ( 
.A1(n_3090),
.A2(n_3019),
.B(n_3017),
.Y(n_3179)
);

AOI221xp5_ASAP7_75t_L g3180 ( 
.A1(n_3176),
.A2(n_3085),
.B1(n_3011),
.B2(n_3035),
.C(n_3077),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_3110),
.B(n_3007),
.Y(n_3181)
);

HB1xp67_ASAP7_75t_L g3182 ( 
.A(n_3101),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3121),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_3132),
.Y(n_3184)
);

OR2x2_ASAP7_75t_L g3185 ( 
.A(n_3126),
.B(n_3066),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_3139),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3131),
.B(n_3010),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3099),
.Y(n_3188)
);

INVx1_ASAP7_75t_SL g3189 ( 
.A(n_3145),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3102),
.Y(n_3190)
);

CKINVDCx20_ASAP7_75t_R g3191 ( 
.A(n_3096),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3136),
.Y(n_3192)
);

NAND3xp33_ASAP7_75t_L g3193 ( 
.A(n_3150),
.B(n_3001),
.C(n_3058),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3106),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_3095),
.B(n_3056),
.Y(n_3195)
);

AOI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_3091),
.A2(n_3061),
.B(n_3012),
.Y(n_3196)
);

AOI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_3092),
.A2(n_3129),
.B(n_3164),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_3111),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3097),
.B(n_3009),
.Y(n_3199)
);

OR2x6_ASAP7_75t_L g3200 ( 
.A(n_3163),
.B(n_3125),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_L g3201 ( 
.A1(n_3174),
.A2(n_2999),
.B(n_3078),
.Y(n_3201)
);

BUFx12f_ASAP7_75t_L g3202 ( 
.A(n_3157),
.Y(n_3202)
);

BUFx3_ASAP7_75t_L g3203 ( 
.A(n_3115),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_3135),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3112),
.Y(n_3205)
);

INVx3_ASAP7_75t_L g3206 ( 
.A(n_3153),
.Y(n_3206)
);

AO21x2_ASAP7_75t_L g3207 ( 
.A1(n_3159),
.A2(n_3064),
.B(n_3047),
.Y(n_3207)
);

OAI21x1_ASAP7_75t_L g3208 ( 
.A1(n_3094),
.A2(n_3074),
.B(n_3076),
.Y(n_3208)
);

OAI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3156),
.A2(n_3008),
.B(n_2992),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_3168),
.B(n_3075),
.Y(n_3210)
);

OR2x6_ASAP7_75t_L g3211 ( 
.A(n_3167),
.B(n_3046),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_3160),
.B(n_2993),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3127),
.Y(n_3213)
);

BUFx3_ASAP7_75t_L g3214 ( 
.A(n_3148),
.Y(n_3214)
);

BUFx2_ASAP7_75t_SL g3215 ( 
.A(n_3120),
.Y(n_3215)
);

BUFx4f_ASAP7_75t_SL g3216 ( 
.A(n_3149),
.Y(n_3216)
);

OA21x2_ASAP7_75t_L g3217 ( 
.A1(n_3142),
.A2(n_3028),
.B(n_3050),
.Y(n_3217)
);

AND2x4_ASAP7_75t_L g3218 ( 
.A(n_3119),
.B(n_3100),
.Y(n_3218)
);

INVx3_ASAP7_75t_L g3219 ( 
.A(n_3147),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3171),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_3161),
.A2(n_3054),
.B(n_3060),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3107),
.B(n_2994),
.Y(n_3222)
);

INVx3_ASAP7_75t_L g3223 ( 
.A(n_3134),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_3104),
.B(n_3108),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3113),
.B(n_379),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3105),
.B(n_380),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3130),
.B(n_381),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3169),
.B(n_382),
.Y(n_3228)
);

AND2x4_ASAP7_75t_L g3229 ( 
.A(n_3175),
.B(n_384),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3154),
.Y(n_3230)
);

INVx3_ASAP7_75t_L g3231 ( 
.A(n_3158),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3154),
.Y(n_3232)
);

NAND2x1p5_ASAP7_75t_L g3233 ( 
.A(n_3151),
.B(n_385),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3177),
.B(n_386),
.Y(n_3234)
);

A2O1A1Ixp33_ASAP7_75t_L g3235 ( 
.A1(n_3114),
.A2(n_389),
.B(n_390),
.C(n_386),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_3109),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3165),
.B(n_3170),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3138),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3123),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3116),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3124),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3172),
.B(n_3173),
.Y(n_3242)
);

OAI21x1_ASAP7_75t_L g3243 ( 
.A1(n_3098),
.A2(n_161),
.B(n_162),
.Y(n_3243)
);

CKINVDCx11_ASAP7_75t_R g3244 ( 
.A(n_3167),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_3118),
.Y(n_3245)
);

BUFx2_ASAP7_75t_L g3246 ( 
.A(n_3143),
.Y(n_3246)
);

NOR2x1_ASAP7_75t_SL g3247 ( 
.A(n_3178),
.B(n_393),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3122),
.Y(n_3248)
);

OR2x2_ASAP7_75t_L g3249 ( 
.A(n_3140),
.B(n_394),
.Y(n_3249)
);

OAI21x1_ASAP7_75t_L g3250 ( 
.A1(n_3128),
.A2(n_167),
.B(n_169),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3137),
.Y(n_3251)
);

INVx2_ASAP7_75t_SL g3252 ( 
.A(n_3155),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_3152),
.A2(n_169),
.B(n_170),
.Y(n_3253)
);

OAI21x1_ASAP7_75t_L g3254 ( 
.A1(n_3162),
.A2(n_169),
.B(n_170),
.Y(n_3254)
);

INVx8_ASAP7_75t_L g3255 ( 
.A(n_3093),
.Y(n_3255)
);

OAI21x1_ASAP7_75t_L g3256 ( 
.A1(n_3144),
.A2(n_171),
.B(n_172),
.Y(n_3256)
);

NOR3xp33_ASAP7_75t_L g3257 ( 
.A(n_3103),
.B(n_171),
.C(n_172),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3182),
.B(n_3166),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3190),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3194),
.Y(n_3260)
);

BUFx3_ASAP7_75t_L g3261 ( 
.A(n_3202),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3198),
.Y(n_3262)
);

BUFx3_ASAP7_75t_L g3263 ( 
.A(n_3214),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3192),
.Y(n_3264)
);

INVx2_ASAP7_75t_SL g3265 ( 
.A(n_3203),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_3181),
.B(n_3141),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3224),
.B(n_3117),
.Y(n_3267)
);

BUFx6f_ASAP7_75t_L g3268 ( 
.A(n_3204),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3205),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3183),
.B(n_3133),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3213),
.Y(n_3271)
);

OAI21x1_ASAP7_75t_L g3272 ( 
.A1(n_3179),
.A2(n_3146),
.B(n_173),
.Y(n_3272)
);

OR2x6_ASAP7_75t_L g3273 ( 
.A(n_3215),
.B(n_395),
.Y(n_3273)
);

CKINVDCx6p67_ASAP7_75t_R g3274 ( 
.A(n_3191),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3220),
.Y(n_3275)
);

INVx3_ASAP7_75t_L g3276 ( 
.A(n_3218),
.Y(n_3276)
);

AO21x2_ASAP7_75t_L g3277 ( 
.A1(n_3238),
.A2(n_173),
.B(n_174),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3184),
.Y(n_3278)
);

INVx1_ASAP7_75t_SL g3279 ( 
.A(n_3189),
.Y(n_3279)
);

BUFx2_ASAP7_75t_L g3280 ( 
.A(n_3200),
.Y(n_3280)
);

INVx4_ASAP7_75t_SL g3281 ( 
.A(n_3216),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3210),
.Y(n_3282)
);

CKINVDCx6p67_ASAP7_75t_R g3283 ( 
.A(n_3244),
.Y(n_3283)
);

INVxp67_ASAP7_75t_L g3284 ( 
.A(n_3187),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3239),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3245),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3185),
.Y(n_3287)
);

BUFx2_ASAP7_75t_L g3288 ( 
.A(n_3200),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_3222),
.B(n_396),
.Y(n_3289)
);

OR2x2_ASAP7_75t_L g3290 ( 
.A(n_3199),
.B(n_396),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3236),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3241),
.Y(n_3292)
);

INVx4_ASAP7_75t_L g3293 ( 
.A(n_3231),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3251),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3240),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_3248),
.Y(n_3296)
);

AND2x4_ASAP7_75t_L g3297 ( 
.A(n_3232),
.B(n_397),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3242),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3212),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3237),
.B(n_400),
.Y(n_3300)
);

AO21x1_ASAP7_75t_SL g3301 ( 
.A1(n_3249),
.A2(n_175),
.B(n_176),
.Y(n_3301)
);

OR2x2_ASAP7_75t_L g3302 ( 
.A(n_3217),
.B(n_401),
.Y(n_3302)
);

AO21x2_ASAP7_75t_L g3303 ( 
.A1(n_3196),
.A2(n_176),
.B(n_177),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3201),
.Y(n_3304)
);

BUFx6f_ASAP7_75t_L g3305 ( 
.A(n_3186),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3243),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3197),
.B(n_3221),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_3223),
.Y(n_3308)
);

NAND2x1p5_ASAP7_75t_L g3309 ( 
.A(n_3219),
.B(n_401),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3225),
.Y(n_3310)
);

HB1xp67_ASAP7_75t_L g3311 ( 
.A(n_3208),
.Y(n_3311)
);

AND2x4_ASAP7_75t_L g3312 ( 
.A(n_3206),
.B(n_402),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3207),
.Y(n_3313)
);

BUFx3_ASAP7_75t_L g3314 ( 
.A(n_3246),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3226),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_3252),
.Y(n_3316)
);

OA21x2_ASAP7_75t_L g3317 ( 
.A1(n_3250),
.A2(n_3253),
.B(n_3256),
.Y(n_3317)
);

INVx2_ASAP7_75t_SL g3318 ( 
.A(n_3229),
.Y(n_3318)
);

INVx3_ASAP7_75t_L g3319 ( 
.A(n_3211),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3247),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3211),
.B(n_405),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3233),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3254),
.Y(n_3323)
);

INVxp67_ASAP7_75t_SL g3324 ( 
.A(n_3193),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_L g3325 ( 
.A(n_3195),
.Y(n_3325)
);

INVx3_ASAP7_75t_L g3326 ( 
.A(n_3255),
.Y(n_3326)
);

INVx3_ASAP7_75t_L g3327 ( 
.A(n_3227),
.Y(n_3327)
);

OR2x2_ASAP7_75t_L g3328 ( 
.A(n_3234),
.B(n_406),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3228),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3209),
.B(n_407),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3257),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3235),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3180),
.B(n_408),
.Y(n_3333)
);

AO21x1_ASAP7_75t_SL g3334 ( 
.A1(n_3230),
.A2(n_178),
.B(n_179),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3188),
.Y(n_3335)
);

AO31x2_ASAP7_75t_L g3336 ( 
.A1(n_3313),
.A2(n_183),
.A3(n_181),
.B(n_182),
.Y(n_3336)
);

CKINVDCx20_ASAP7_75t_R g3337 ( 
.A(n_3274),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3285),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3331),
.A2(n_3324),
.B1(n_3333),
.B2(n_3303),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_3332),
.A2(n_410),
.B1(n_411),
.B2(n_409),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3286),
.Y(n_3341)
);

CKINVDCx5p33_ASAP7_75t_R g3342 ( 
.A(n_3283),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3298),
.B(n_185),
.Y(n_3343)
);

AOI21xp33_ASAP7_75t_L g3344 ( 
.A1(n_3329),
.A2(n_411),
.B(n_410),
.Y(n_3344)
);

AND2x4_ASAP7_75t_L g3345 ( 
.A(n_3319),
.B(n_413),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3280),
.B(n_185),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3288),
.B(n_186),
.Y(n_3347)
);

BUFx6f_ASAP7_75t_L g3348 ( 
.A(n_3268),
.Y(n_3348)
);

NAND4xp25_ASAP7_75t_L g3349 ( 
.A(n_3300),
.B(n_188),
.C(n_186),
.D(n_187),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3259),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3325),
.A2(n_417),
.B1(n_418),
.B2(n_416),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3260),
.Y(n_3352)
);

A2O1A1Ixp33_ASAP7_75t_L g3353 ( 
.A1(n_3330),
.A2(n_417),
.B(n_419),
.C(n_416),
.Y(n_3353)
);

OAI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3326),
.A2(n_194),
.B1(n_191),
.B2(n_193),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_L g3355 ( 
.A1(n_3315),
.A2(n_421),
.B1(n_422),
.B2(n_420),
.Y(n_3355)
);

INVxp67_ASAP7_75t_L g3356 ( 
.A(n_3310),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3320),
.A2(n_423),
.B1(n_424),
.B2(n_422),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_3322),
.A2(n_425),
.B1(n_426),
.B2(n_423),
.Y(n_3358)
);

NOR2x1_ASAP7_75t_SL g3359 ( 
.A(n_3334),
.B(n_191),
.Y(n_3359)
);

OR2x2_ASAP7_75t_L g3360 ( 
.A(n_3287),
.B(n_191),
.Y(n_3360)
);

OAI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3284),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_3361)
);

OR2x6_ASAP7_75t_L g3362 ( 
.A(n_3265),
.B(n_425),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3269),
.Y(n_3363)
);

AOI22xp33_ASAP7_75t_L g3364 ( 
.A1(n_3327),
.A2(n_428),
.B1(n_429),
.B2(n_427),
.Y(n_3364)
);

BUFx4f_ASAP7_75t_SL g3365 ( 
.A(n_3261),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3335),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3275),
.Y(n_3367)
);

OAI221xp5_ASAP7_75t_L g3368 ( 
.A1(n_3328),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.C(n_201),
.Y(n_3368)
);

AND2x4_ASAP7_75t_SL g3369 ( 
.A(n_3293),
.B(n_430),
.Y(n_3369)
);

AOI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_3273),
.A2(n_433),
.B1(n_434),
.B2(n_432),
.Y(n_3370)
);

OR2x2_ASAP7_75t_L g3371 ( 
.A(n_3282),
.B(n_199),
.Y(n_3371)
);

OAI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3267),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_3372)
);

HB1xp67_ASAP7_75t_L g3373 ( 
.A(n_3258),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3262),
.Y(n_3374)
);

AOI222xp33_ASAP7_75t_L g3375 ( 
.A1(n_3270),
.A2(n_207),
.B1(n_209),
.B2(n_205),
.C1(n_206),
.C2(n_208),
.Y(n_3375)
);

OAI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3302),
.A2(n_437),
.B1(n_438),
.B2(n_436),
.Y(n_3376)
);

AOI21xp33_ASAP7_75t_L g3377 ( 
.A1(n_3323),
.A2(n_441),
.B(n_439),
.Y(n_3377)
);

AOI22xp33_ASAP7_75t_L g3378 ( 
.A1(n_3277),
.A2(n_443),
.B1(n_444),
.B2(n_442),
.Y(n_3378)
);

OAI221xp5_ASAP7_75t_L g3379 ( 
.A1(n_3290),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.C(n_215),
.Y(n_3379)
);

OAI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3316),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_3308),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_3314),
.B(n_442),
.Y(n_3382)
);

INVx3_ASAP7_75t_L g3383 ( 
.A(n_3276),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3264),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3292),
.Y(n_3385)
);

AOI221xp5_ASAP7_75t_L g3386 ( 
.A1(n_3304),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.C(n_219),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3278),
.B(n_446),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3279),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_3388)
);

OA21x2_ASAP7_75t_L g3389 ( 
.A1(n_3295),
.A2(n_226),
.B(n_227),
.Y(n_3389)
);

OAI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3299),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3318),
.A2(n_448),
.B1(n_450),
.B2(n_447),
.Y(n_3391)
);

BUFx6f_ASAP7_75t_L g3392 ( 
.A(n_3305),
.Y(n_3392)
);

OAI21xp33_ASAP7_75t_L g3393 ( 
.A1(n_3311),
.A2(n_228),
.B(n_229),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3296),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3291),
.Y(n_3395)
);

OAI21xp33_ASAP7_75t_SL g3396 ( 
.A1(n_3266),
.A2(n_228),
.B(n_229),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_L g3397 ( 
.A1(n_3301),
.A2(n_450),
.B1(n_451),
.B2(n_448),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3294),
.Y(n_3398)
);

OAI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3309),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3306),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3289),
.B(n_234),
.Y(n_3401)
);

BUFx3_ASAP7_75t_L g3402 ( 
.A(n_3305),
.Y(n_3402)
);

OAI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3317),
.A2(n_452),
.B1(n_453),
.B2(n_451),
.Y(n_3403)
);

NAND4xp25_ASAP7_75t_L g3404 ( 
.A(n_3321),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_3404)
);

INVx8_ASAP7_75t_L g3405 ( 
.A(n_3312),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3272),
.Y(n_3406)
);

OAI22xp5_ASAP7_75t_L g3407 ( 
.A1(n_3297),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_3407)
);

OA21x2_ASAP7_75t_L g3408 ( 
.A1(n_3281),
.A2(n_237),
.B(n_238),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3285),
.Y(n_3409)
);

CKINVDCx5p33_ASAP7_75t_R g3410 ( 
.A(n_3274),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_3307),
.A2(n_455),
.B1(n_456),
.B2(n_454),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3298),
.B(n_239),
.Y(n_3412)
);

INVx3_ASAP7_75t_L g3413 ( 
.A(n_3263),
.Y(n_3413)
);

AND2x4_ASAP7_75t_L g3414 ( 
.A(n_3319),
.B(n_457),
.Y(n_3414)
);

AOI22xp33_ASAP7_75t_L g3415 ( 
.A1(n_3307),
.A2(n_459),
.B1(n_460),
.B2(n_457),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3285),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_L g3417 ( 
.A1(n_3307),
.A2(n_460),
.B1(n_461),
.B2(n_459),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3285),
.Y(n_3418)
);

OAI221xp5_ASAP7_75t_L g3419 ( 
.A1(n_3307),
.A2(n_466),
.B1(n_463),
.B2(n_464),
.C(n_467),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3271),
.Y(n_3420)
);

AND2x4_ASAP7_75t_L g3421 ( 
.A(n_3319),
.B(n_466),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3285),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3394),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3338),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3409),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3416),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3419),
.A2(n_473),
.B1(n_470),
.B2(n_471),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3383),
.B(n_474),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3381),
.B(n_474),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3418),
.Y(n_3430)
);

HB1xp67_ASAP7_75t_L g3431 ( 
.A(n_3406),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3339),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3422),
.Y(n_3433)
);

BUFx2_ASAP7_75t_L g3434 ( 
.A(n_3337),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3385),
.Y(n_3435)
);

AND2x4_ASAP7_75t_L g3436 ( 
.A(n_3413),
.B(n_477),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3350),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3352),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3363),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3374),
.B(n_480),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_3375),
.A2(n_483),
.B1(n_480),
.B2(n_482),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3366),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3384),
.B(n_484),
.Y(n_3443)
);

CKINVDCx16_ASAP7_75t_R g3444 ( 
.A(n_3402),
.Y(n_3444)
);

OR2x2_ASAP7_75t_L g3445 ( 
.A(n_3400),
.B(n_485),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3367),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_3392),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3420),
.B(n_487),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3341),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3395),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3398),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3343),
.B(n_488),
.Y(n_3452)
);

BUFx2_ASAP7_75t_L g3453 ( 
.A(n_3410),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3360),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_3371),
.B(n_489),
.Y(n_3455)
);

INVx1_ASAP7_75t_SL g3456 ( 
.A(n_3365),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3404),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3346),
.B(n_491),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3347),
.B(n_493),
.Y(n_3459)
);

AND2x4_ASAP7_75t_L g3460 ( 
.A(n_3412),
.B(n_494),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3389),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3349),
.A2(n_497),
.B1(n_494),
.B2(n_495),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3336),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_3348),
.B(n_498),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3387),
.Y(n_3465)
);

BUFx2_ASAP7_75t_L g3466 ( 
.A(n_3362),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3396),
.B(n_501),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3403),
.B(n_502),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3386),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3401),
.B(n_3345),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3414),
.B(n_505),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3421),
.B(n_506),
.Y(n_3472)
);

BUFx2_ASAP7_75t_L g3473 ( 
.A(n_3405),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3408),
.B(n_507),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3376),
.B(n_508),
.Y(n_3475)
);

INVx3_ASAP7_75t_L g3476 ( 
.A(n_3369),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3353),
.B(n_509),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3359),
.B(n_3382),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3393),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3379),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3377),
.B(n_510),
.Y(n_3481)
);

OR2x2_ASAP7_75t_L g3482 ( 
.A(n_3407),
.B(n_511),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3397),
.B(n_511),
.Y(n_3483)
);

INVx3_ASAP7_75t_L g3484 ( 
.A(n_3344),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3368),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3390),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3361),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3391),
.B(n_512),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3378),
.B(n_513),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3380),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3399),
.Y(n_3491)
);

INVxp33_ASAP7_75t_SL g3492 ( 
.A(n_3388),
.Y(n_3492)
);

OR2x2_ASAP7_75t_L g3493 ( 
.A(n_3372),
.B(n_514),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3411),
.B(n_515),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3354),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3355),
.B(n_519),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3370),
.B(n_521),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_L g3498 ( 
.A1(n_3415),
.A2(n_526),
.B1(n_523),
.B2(n_524),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3351),
.B(n_526),
.Y(n_3499)
);

AND2x4_ASAP7_75t_L g3500 ( 
.A(n_3417),
.B(n_527),
.Y(n_3500)
);

AND2x4_ASAP7_75t_L g3501 ( 
.A(n_3358),
.B(n_528),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3364),
.Y(n_3502)
);

INVxp67_ASAP7_75t_SL g3503 ( 
.A(n_3357),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3340),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3338),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3383),
.B(n_531),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3338),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_3373),
.B(n_533),
.Y(n_3508)
);

OR2x2_ASAP7_75t_L g3509 ( 
.A(n_3373),
.B(n_534),
.Y(n_3509)
);

INVxp67_ASAP7_75t_SL g3510 ( 
.A(n_3373),
.Y(n_3510)
);

HB1xp67_ASAP7_75t_L g3511 ( 
.A(n_3373),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3383),
.B(n_534),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3383),
.B(n_535),
.Y(n_3513)
);

BUFx12f_ASAP7_75t_L g3514 ( 
.A(n_3342),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3383),
.B(n_536),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3338),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3338),
.Y(n_3517)
);

OR2x2_ASAP7_75t_L g3518 ( 
.A(n_3373),
.B(n_538),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3356),
.B(n_539),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3394),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3444),
.B(n_540),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3424),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3425),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_3514),
.B(n_543),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_3466),
.B(n_544),
.Y(n_3525)
);

AND2x4_ASAP7_75t_L g3526 ( 
.A(n_3447),
.B(n_545),
.Y(n_3526)
);

HB1xp67_ASAP7_75t_L g3527 ( 
.A(n_3461),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3510),
.B(n_546),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3511),
.B(n_548),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3423),
.Y(n_3530)
);

HB1xp67_ASAP7_75t_L g3531 ( 
.A(n_3431),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3484),
.B(n_549),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3520),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3426),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3450),
.B(n_552),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3433),
.Y(n_3536)
);

HB1xp67_ASAP7_75t_L g3537 ( 
.A(n_3463),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3453),
.B(n_554),
.Y(n_3538)
);

AND2x4_ASAP7_75t_L g3539 ( 
.A(n_3434),
.B(n_3428),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3435),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3451),
.B(n_555),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3430),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3449),
.B(n_556),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3478),
.B(n_557),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3437),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3438),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3439),
.Y(n_3547)
);

AND2x4_ASAP7_75t_L g3548 ( 
.A(n_3506),
.B(n_558),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3442),
.Y(n_3549)
);

AND2x4_ASAP7_75t_L g3550 ( 
.A(n_3512),
.B(n_559),
.Y(n_3550)
);

AND2x4_ASAP7_75t_L g3551 ( 
.A(n_3513),
.B(n_559),
.Y(n_3551)
);

NAND2xp33_ASAP7_75t_R g3552 ( 
.A(n_3492),
.B(n_1353),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3446),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3440),
.B(n_560),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3505),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3470),
.B(n_3491),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3507),
.Y(n_3557)
);

OR2x2_ASAP7_75t_L g3558 ( 
.A(n_3508),
.B(n_561),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3516),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3517),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3445),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3443),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3448),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3486),
.B(n_562),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3429),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3509),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3515),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3490),
.B(n_562),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3518),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_3476),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3519),
.Y(n_3571)
);

AND2x2_ASAP7_75t_L g3572 ( 
.A(n_3495),
.B(n_563),
.Y(n_3572)
);

BUFx6f_ASAP7_75t_L g3573 ( 
.A(n_3436),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3487),
.B(n_564),
.Y(n_3574)
);

AND2x4_ASAP7_75t_L g3575 ( 
.A(n_3456),
.B(n_565),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3479),
.B(n_567),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3455),
.B(n_568),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3474),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3464),
.Y(n_3579)
);

INVxp67_ASAP7_75t_L g3580 ( 
.A(n_3480),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3460),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3467),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3485),
.B(n_569),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3458),
.B(n_570),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3503),
.B(n_571),
.Y(n_3585)
);

HB1xp67_ASAP7_75t_L g3586 ( 
.A(n_3502),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3459),
.B(n_571),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3471),
.B(n_572),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3472),
.B(n_573),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3452),
.B(n_573),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_3468),
.Y(n_3591)
);

HB1xp67_ASAP7_75t_L g3592 ( 
.A(n_3482),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3475),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3481),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3493),
.Y(n_3595)
);

OR2x2_ASAP7_75t_L g3596 ( 
.A(n_3477),
.B(n_575),
.Y(n_3596)
);

HB1xp67_ASAP7_75t_L g3597 ( 
.A(n_3499),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3432),
.B(n_576),
.Y(n_3598)
);

NAND2x1_ASAP7_75t_L g3599 ( 
.A(n_3497),
.B(n_578),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3427),
.B(n_577),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3483),
.B(n_577),
.Y(n_3601)
);

HB1xp67_ASAP7_75t_L g3602 ( 
.A(n_3494),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3489),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3488),
.B(n_579),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3500),
.B(n_580),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_L g3606 ( 
.A(n_3496),
.B(n_582),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3501),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3457),
.B(n_584),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_3462),
.B(n_585),
.Y(n_3609)
);

OR2x2_ASAP7_75t_L g3610 ( 
.A(n_3441),
.B(n_586),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3469),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3498),
.Y(n_3612)
);

AND2x4_ASAP7_75t_L g3613 ( 
.A(n_3504),
.B(n_586),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3465),
.B(n_587),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3424),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_3473),
.B(n_587),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3473),
.B(n_588),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3424),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3424),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3473),
.B(n_588),
.Y(n_3620)
);

OR2x2_ASAP7_75t_L g3621 ( 
.A(n_3454),
.B(n_589),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3423),
.Y(n_3622)
);

BUFx6f_ASAP7_75t_L g3623 ( 
.A(n_3514),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3473),
.B(n_592),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3473),
.B(n_594),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3473),
.B(n_595),
.Y(n_3626)
);

HB1xp67_ASAP7_75t_L g3627 ( 
.A(n_3461),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3465),
.B(n_598),
.Y(n_3628)
);

INVx4_ASAP7_75t_L g3629 ( 
.A(n_3514),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3444),
.B(n_599),
.Y(n_3630)
);

INVx1_ASAP7_75t_SL g3631 ( 
.A(n_3453),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3423),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3424),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3424),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3473),
.B(n_600),
.Y(n_3635)
);

AND2x2_ASAP7_75t_L g3636 ( 
.A(n_3473),
.B(n_601),
.Y(n_3636)
);

BUFx2_ASAP7_75t_L g3637 ( 
.A(n_3466),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3424),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3473),
.B(n_602),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3465),
.B(n_603),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_SL g3641 ( 
.A(n_3631),
.B(n_3637),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3582),
.B(n_604),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3522),
.Y(n_3643)
);

BUFx2_ASAP7_75t_L g3644 ( 
.A(n_3629),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3523),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3534),
.Y(n_3646)
);

AOI221xp5_ASAP7_75t_L g3647 ( 
.A1(n_3586),
.A2(n_607),
.B1(n_605),
.B2(n_606),
.C(n_608),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3536),
.Y(n_3648)
);

OAI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3552),
.A2(n_609),
.B1(n_606),
.B2(n_607),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3593),
.B(n_609),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3570),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3556),
.B(n_610),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_L g3653 ( 
.A(n_3623),
.B(n_612),
.Y(n_3653)
);

OAI322xp33_ASAP7_75t_L g3654 ( 
.A1(n_3585),
.A2(n_618),
.A3(n_617),
.B1(n_615),
.B2(n_613),
.C1(n_614),
.C2(n_616),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3540),
.Y(n_3655)
);

AOI221xp5_ASAP7_75t_L g3656 ( 
.A1(n_3591),
.A2(n_617),
.B1(n_613),
.B2(n_616),
.C(n_618),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3592),
.B(n_620),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3578),
.B(n_620),
.Y(n_3658)
);

AOI22xp33_ASAP7_75t_L g3659 ( 
.A1(n_3611),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3545),
.Y(n_3660)
);

HB1xp67_ASAP7_75t_L g3661 ( 
.A(n_3527),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3547),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3539),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3579),
.Y(n_3664)
);

HB1xp67_ASAP7_75t_L g3665 ( 
.A(n_3627),
.Y(n_3665)
);

BUFx3_ASAP7_75t_L g3666 ( 
.A(n_3573),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_L g3667 ( 
.A(n_3580),
.B(n_625),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3565),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3567),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3595),
.B(n_628),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3561),
.B(n_629),
.Y(n_3671)
);

AOI222xp33_ASAP7_75t_L g3672 ( 
.A1(n_3609),
.A2(n_632),
.B1(n_634),
.B2(n_630),
.C1(n_631),
.C2(n_633),
.Y(n_3672)
);

INVx3_ASAP7_75t_L g3673 ( 
.A(n_3573),
.Y(n_3673)
);

OAI21xp5_ASAP7_75t_SL g3674 ( 
.A1(n_3608),
.A2(n_637),
.B(n_636),
.Y(n_3674)
);

AOI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3602),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_3675)
);

INVx1_ASAP7_75t_SL g3676 ( 
.A(n_3521),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3555),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3597),
.B(n_639),
.Y(n_3678)
);

NAND3xp33_ASAP7_75t_SL g3679 ( 
.A(n_3630),
.B(n_641),
.C(n_642),
.Y(n_3679)
);

OAI221xp5_ASAP7_75t_L g3680 ( 
.A1(n_3596),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.C(n_647),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3557),
.Y(n_3681)
);

NOR2xp33_ASAP7_75t_L g3682 ( 
.A(n_3594),
.B(n_3571),
.Y(n_3682)
);

OAI211xp5_ASAP7_75t_L g3683 ( 
.A1(n_3600),
.A2(n_650),
.B(n_648),
.C(n_649),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_3581),
.B(n_650),
.Y(n_3684)
);

NAND4xp25_ASAP7_75t_L g3685 ( 
.A(n_3606),
.B(n_653),
.C(n_654),
.D(n_652),
.Y(n_3685)
);

AND2x4_ASAP7_75t_L g3686 ( 
.A(n_3563),
.B(n_651),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3566),
.B(n_3569),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3530),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3583),
.B(n_3576),
.Y(n_3689)
);

OR2x2_ASAP7_75t_L g3690 ( 
.A(n_3533),
.B(n_655),
.Y(n_3690)
);

OAI321xp33_ASAP7_75t_L g3691 ( 
.A1(n_3598),
.A2(n_659),
.A3(n_661),
.B1(n_657),
.B2(n_658),
.C(n_660),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3559),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3544),
.B(n_658),
.Y(n_3693)
);

HB1xp67_ASAP7_75t_L g3694 ( 
.A(n_3531),
.Y(n_3694)
);

INVx2_ASAP7_75t_SL g3695 ( 
.A(n_3616),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3562),
.B(n_660),
.Y(n_3696)
);

HB1xp67_ASAP7_75t_L g3697 ( 
.A(n_3537),
.Y(n_3697)
);

OR2x6_ASAP7_75t_L g3698 ( 
.A(n_3599),
.B(n_662),
.Y(n_3698)
);

AND2x2_ASAP7_75t_SL g3699 ( 
.A(n_3613),
.B(n_663),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3560),
.Y(n_3700)
);

AOI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3612),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3615),
.Y(n_3702)
);

AOI221xp5_ASAP7_75t_L g3703 ( 
.A1(n_3532),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.C(n_668),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3618),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3619),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3622),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3603),
.B(n_670),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3607),
.B(n_670),
.Y(n_3708)
);

HB1xp67_ASAP7_75t_L g3709 ( 
.A(n_3542),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3546),
.Y(n_3710)
);

AOI211xp5_ASAP7_75t_L g3711 ( 
.A1(n_3610),
.A2(n_674),
.B(n_671),
.C(n_673),
.Y(n_3711)
);

AO21x2_ASAP7_75t_L g3712 ( 
.A1(n_3528),
.A2(n_674),
.B(n_676),
.Y(n_3712)
);

CKINVDCx20_ASAP7_75t_R g3713 ( 
.A(n_3524),
.Y(n_3713)
);

AND2x2_ASAP7_75t_SL g3714 ( 
.A(n_3525),
.B(n_678),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_3632),
.B(n_679),
.Y(n_3715)
);

INVx1_ASAP7_75t_SL g3716 ( 
.A(n_3538),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3564),
.B(n_680),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3568),
.B(n_681),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_L g3719 ( 
.A1(n_3549),
.A2(n_683),
.B1(n_681),
.B2(n_682),
.Y(n_3719)
);

NAND3xp33_ASAP7_75t_L g3720 ( 
.A(n_3614),
.B(n_682),
.C(n_683),
.Y(n_3720)
);

HB1xp67_ASAP7_75t_L g3721 ( 
.A(n_3553),
.Y(n_3721)
);

AOI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3574),
.A2(n_686),
.B1(n_684),
.B2(n_685),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3633),
.Y(n_3723)
);

A2O1A1Ixp33_ASAP7_75t_L g3724 ( 
.A1(n_3604),
.A2(n_688),
.B(n_686),
.C(n_687),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_3529),
.B(n_690),
.Y(n_3725)
);

HB1xp67_ASAP7_75t_L g3726 ( 
.A(n_3634),
.Y(n_3726)
);

AOI211xp5_ASAP7_75t_L g3727 ( 
.A1(n_3601),
.A2(n_693),
.B(n_691),
.C(n_692),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3535),
.B(n_694),
.Y(n_3728)
);

OAI221xp5_ASAP7_75t_L g3729 ( 
.A1(n_3628),
.A2(n_699),
.B1(n_695),
.B2(n_696),
.C(n_700),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3638),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3572),
.B(n_696),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3640),
.A2(n_704),
.B1(n_701),
.B2(n_702),
.Y(n_3732)
);

AOI22xp33_ASAP7_75t_L g3733 ( 
.A1(n_3605),
.A2(n_706),
.B1(n_704),
.B2(n_705),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3590),
.B(n_706),
.Y(n_3734)
);

AND2x4_ASAP7_75t_L g3735 ( 
.A(n_3617),
.B(n_707),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3541),
.Y(n_3736)
);

AND2x4_ASAP7_75t_L g3737 ( 
.A(n_3620),
.B(n_707),
.Y(n_3737)
);

BUFx3_ASAP7_75t_L g3738 ( 
.A(n_3575),
.Y(n_3738)
);

OAI22xp33_ASAP7_75t_L g3739 ( 
.A1(n_3621),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3543),
.B(n_709),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3694),
.Y(n_3741)
);

AND2x4_ASAP7_75t_L g3742 ( 
.A(n_3666),
.B(n_3526),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3644),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3726),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3661),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3665),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3676),
.B(n_3624),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3673),
.B(n_3625),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3710),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3721),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3695),
.Y(n_3751)
);

INVx6_ASAP7_75t_L g3752 ( 
.A(n_3698),
.Y(n_3752)
);

AND2x4_ASAP7_75t_L g3753 ( 
.A(n_3651),
.B(n_3626),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3697),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3687),
.Y(n_3755)
);

INVx3_ASAP7_75t_L g3756 ( 
.A(n_3738),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3730),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3663),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3643),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3716),
.B(n_3635),
.Y(n_3760)
);

OAI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3649),
.A2(n_3554),
.B(n_3636),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3690),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3689),
.B(n_3639),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3645),
.Y(n_3764)
);

AOI21xp33_ASAP7_75t_L g3765 ( 
.A1(n_3641),
.A2(n_3577),
.B(n_3558),
.Y(n_3765)
);

INVx1_ASAP7_75t_SL g3766 ( 
.A(n_3714),
.Y(n_3766)
);

CKINVDCx16_ASAP7_75t_R g3767 ( 
.A(n_3713),
.Y(n_3767)
);

OR2x2_ASAP7_75t_L g3768 ( 
.A(n_3736),
.B(n_3584),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3664),
.B(n_3588),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3646),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3668),
.B(n_3589),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3669),
.B(n_3587),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3648),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3712),
.B(n_3548),
.Y(n_3774)
);

NOR3xp33_ASAP7_75t_L g3775 ( 
.A(n_3691),
.B(n_3551),
.C(n_3550),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3655),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3660),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3652),
.B(n_3707),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3662),
.Y(n_3779)
);

HB1xp67_ASAP7_75t_L g3780 ( 
.A(n_3709),
.Y(n_3780)
);

NOR2xp67_ASAP7_75t_L g3781 ( 
.A(n_3682),
.B(n_711),
.Y(n_3781)
);

AND2x2_ASAP7_75t_SL g3782 ( 
.A(n_3699),
.B(n_713),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3696),
.B(n_714),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3708),
.B(n_3658),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3677),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3678),
.B(n_715),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3688),
.B(n_1351),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3681),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3657),
.B(n_716),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3692),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3717),
.B(n_716),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3718),
.B(n_717),
.Y(n_3792)
);

NOR2xp67_ASAP7_75t_L g3793 ( 
.A(n_3670),
.B(n_717),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3700),
.Y(n_3794)
);

AOI22xp33_ASAP7_75t_L g3795 ( 
.A1(n_3685),
.A2(n_3679),
.B1(n_3672),
.B2(n_3729),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3702),
.Y(n_3796)
);

NAND3xp33_ASAP7_75t_L g3797 ( 
.A(n_3711),
.B(n_719),
.C(n_720),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3706),
.B(n_721),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3704),
.Y(n_3799)
);

AOI22xp5_ASAP7_75t_L g3800 ( 
.A1(n_3647),
.A2(n_3674),
.B1(n_3656),
.B2(n_3683),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3705),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3667),
.B(n_722),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3734),
.B(n_3642),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3715),
.Y(n_3804)
);

AND2x4_ASAP7_75t_L g3805 ( 
.A(n_3684),
.B(n_1363),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3671),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3731),
.B(n_724),
.Y(n_3807)
);

INVx4_ASAP7_75t_L g3808 ( 
.A(n_3735),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3725),
.B(n_725),
.Y(n_3809)
);

BUFx2_ASAP7_75t_L g3810 ( 
.A(n_3737),
.Y(n_3810)
);

NOR3xp33_ASAP7_75t_L g3811 ( 
.A(n_3654),
.B(n_725),
.C(n_726),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3650),
.B(n_727),
.Y(n_3812)
);

NAND2x1p5_ASAP7_75t_L g3813 ( 
.A(n_3686),
.B(n_728),
.Y(n_3813)
);

INVx3_ASAP7_75t_L g3814 ( 
.A(n_3808),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3767),
.B(n_3740),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3752),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3752),
.Y(n_3817)
);

AOI32xp33_ASAP7_75t_L g3818 ( 
.A1(n_3811),
.A2(n_3727),
.A3(n_3739),
.B1(n_3703),
.B2(n_3732),
.Y(n_3818)
);

CKINVDCx16_ASAP7_75t_R g3819 ( 
.A(n_3766),
.Y(n_3819)
);

INVx2_ASAP7_75t_SL g3820 ( 
.A(n_3742),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3780),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3741),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3748),
.B(n_3653),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3810),
.B(n_3722),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3747),
.B(n_3720),
.Y(n_3825)
);

OR2x2_ASAP7_75t_L g3826 ( 
.A(n_3760),
.B(n_3723),
.Y(n_3826)
);

HB1xp67_ASAP7_75t_L g3827 ( 
.A(n_3781),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3768),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3756),
.B(n_3693),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3745),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3743),
.B(n_3728),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3746),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3754),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3787),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3755),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3744),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3762),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3784),
.B(n_3724),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3778),
.B(n_3733),
.Y(n_3839)
);

OR2x2_ASAP7_75t_L g3840 ( 
.A(n_3763),
.B(n_3680),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3753),
.Y(n_3841)
);

AND2x4_ASAP7_75t_L g3842 ( 
.A(n_3751),
.B(n_3675),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3804),
.Y(n_3843)
);

OR2x2_ASAP7_75t_L g3844 ( 
.A(n_3806),
.B(n_3701),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3749),
.Y(n_3845)
);

INVx1_ASAP7_75t_SL g3846 ( 
.A(n_3782),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3769),
.B(n_3659),
.Y(n_3847)
);

INVxp67_ASAP7_75t_L g3848 ( 
.A(n_3774),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3750),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3771),
.B(n_3719),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3772),
.B(n_728),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3758),
.B(n_729),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3798),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3761),
.B(n_729),
.Y(n_3854)
);

INVxp67_ASAP7_75t_SL g3855 ( 
.A(n_3793),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3757),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3813),
.Y(n_3857)
);

OR2x2_ASAP7_75t_L g3858 ( 
.A(n_3803),
.B(n_730),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3759),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3805),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3765),
.B(n_730),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_3764),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3800),
.B(n_731),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3795),
.B(n_732),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3791),
.B(n_733),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3792),
.B(n_733),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3809),
.B(n_734),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3770),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3807),
.B(n_3789),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3786),
.B(n_735),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3783),
.B(n_736),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3773),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3775),
.B(n_737),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3776),
.B(n_738),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3777),
.B(n_3779),
.Y(n_3875)
);

OR2x2_ASAP7_75t_L g3876 ( 
.A(n_3812),
.B(n_739),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3797),
.B(n_741),
.Y(n_3877)
);

INVxp67_ASAP7_75t_L g3878 ( 
.A(n_3802),
.Y(n_3878)
);

INVxp33_ASAP7_75t_L g3879 ( 
.A(n_3785),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3788),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3790),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3794),
.B(n_742),
.Y(n_3882)
);

INVxp67_ASAP7_75t_L g3883 ( 
.A(n_3796),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3799),
.B(n_742),
.Y(n_3884)
);

AND3x2_ASAP7_75t_L g3885 ( 
.A(n_3801),
.B(n_743),
.C(n_744),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3855),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3821),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3827),
.Y(n_3888)
);

INVx1_ASAP7_75t_SL g3889 ( 
.A(n_3846),
.Y(n_3889)
);

NAND3xp33_ASAP7_75t_L g3890 ( 
.A(n_3848),
.B(n_746),
.C(n_747),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3874),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3814),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3820),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3882),
.Y(n_3894)
);

INVx1_ASAP7_75t_SL g3895 ( 
.A(n_3823),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3816),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3884),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3869),
.B(n_748),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3817),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3862),
.Y(n_3900)
);

AOI32xp33_ASAP7_75t_L g3901 ( 
.A1(n_3873),
.A2(n_751),
.A3(n_749),
.B1(n_750),
.B2(n_752),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3828),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3838),
.B(n_753),
.Y(n_3903)
);

AOI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3864),
.A2(n_756),
.B1(n_754),
.B2(n_755),
.Y(n_3904)
);

NOR3xp33_ASAP7_75t_L g3905 ( 
.A(n_3878),
.B(n_754),
.C(n_755),
.Y(n_3905)
);

OAI21xp5_ASAP7_75t_SL g3906 ( 
.A1(n_3854),
.A2(n_758),
.B(n_757),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3852),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3834),
.Y(n_3908)
);

NAND4xp25_ASAP7_75t_SL g3909 ( 
.A(n_3863),
.B(n_3824),
.C(n_3825),
.D(n_3840),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3851),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3822),
.Y(n_3911)
);

INVx1_ASAP7_75t_SL g3912 ( 
.A(n_3885),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3830),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3832),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_SL g3915 ( 
.A1(n_3847),
.A2(n_3850),
.B1(n_3839),
.B2(n_3842),
.Y(n_3915)
);

NOR2xp33_ASAP7_75t_SL g3916 ( 
.A(n_3857),
.B(n_1356),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3877),
.A2(n_759),
.B(n_760),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3833),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3837),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3860),
.B(n_761),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3829),
.B(n_3841),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3843),
.Y(n_3922)
);

OAI221xp5_ASAP7_75t_L g3923 ( 
.A1(n_3844),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.C(n_765),
.Y(n_3923)
);

AOI221xp5_ASAP7_75t_L g3924 ( 
.A1(n_3879),
.A2(n_769),
.B1(n_767),
.B2(n_768),
.C(n_770),
.Y(n_3924)
);

NOR2xp67_ASAP7_75t_SL g3925 ( 
.A(n_3858),
.B(n_772),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3831),
.B(n_1358),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3853),
.B(n_1359),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3861),
.B(n_774),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3871),
.Y(n_3929)
);

AOI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_3845),
.A2(n_777),
.B1(n_774),
.B2(n_776),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3849),
.B(n_3836),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3826),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3875),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3870),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3876),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3835),
.B(n_3865),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3866),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3867),
.Y(n_3938)
);

OAI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3883),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3859),
.Y(n_3940)
);

OAI21xp5_ASAP7_75t_L g3941 ( 
.A1(n_3856),
.A2(n_782),
.B(n_783),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3868),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3872),
.B(n_1352),
.Y(n_3943)
);

OR2x2_ASAP7_75t_L g3944 ( 
.A(n_3880),
.B(n_784),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3881),
.B(n_785),
.Y(n_3945)
);

OAI21xp5_ASAP7_75t_SL g3946 ( 
.A1(n_3818),
.A2(n_787),
.B(n_786),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3819),
.B(n_785),
.Y(n_3947)
);

AND2x2_ASAP7_75t_L g3948 ( 
.A(n_3815),
.B(n_1361),
.Y(n_3948)
);

NAND2x1_ASAP7_75t_SL g3949 ( 
.A(n_3827),
.B(n_786),
.Y(n_3949)
);

INVx1_ASAP7_75t_SL g3950 ( 
.A(n_3846),
.Y(n_3950)
);

OR2x2_ASAP7_75t_L g3951 ( 
.A(n_3819),
.B(n_789),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3815),
.Y(n_3952)
);

NOR2x1_ASAP7_75t_L g3953 ( 
.A(n_3951),
.B(n_789),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3912),
.B(n_790),
.Y(n_3954)
);

NAND3xp33_ASAP7_75t_SL g3955 ( 
.A(n_3946),
.B(n_791),
.C(n_792),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3888),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3889),
.A2(n_797),
.B1(n_793),
.B2(n_794),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3950),
.B(n_797),
.Y(n_3958)
);

OAI21xp33_ASAP7_75t_L g3959 ( 
.A1(n_3893),
.A2(n_3892),
.B(n_3895),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3921),
.B(n_798),
.Y(n_3960)
);

INVxp67_ASAP7_75t_L g3961 ( 
.A(n_3916),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3948),
.B(n_802),
.Y(n_3962)
);

AOI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3896),
.A2(n_806),
.B1(n_804),
.B2(n_805),
.Y(n_3963)
);

AOI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3899),
.A2(n_810),
.B1(n_808),
.B2(n_809),
.Y(n_3964)
);

INVxp67_ASAP7_75t_L g3965 ( 
.A(n_3925),
.Y(n_3965)
);

NAND2xp33_ASAP7_75t_L g3966 ( 
.A(n_3901),
.B(n_811),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3926),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_3906),
.B(n_812),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3936),
.Y(n_3969)
);

AOI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3910),
.A2(n_3934),
.B1(n_3937),
.B2(n_3929),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3938),
.Y(n_3971)
);

NAND3xp33_ASAP7_75t_L g3972 ( 
.A(n_3900),
.B(n_815),
.C(n_816),
.Y(n_3972)
);

OR3x1_ASAP7_75t_L g3973 ( 
.A(n_3891),
.B(n_817),
.C(n_818),
.Y(n_3973)
);

OR2x2_ASAP7_75t_L g3974 ( 
.A(n_3903),
.B(n_817),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3933),
.B(n_819),
.Y(n_3975)
);

NOR2xp33_ASAP7_75t_L g3976 ( 
.A(n_3894),
.B(n_820),
.Y(n_3976)
);

AOI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3897),
.A2(n_3905),
.B1(n_3907),
.B2(n_3887),
.Y(n_3977)
);

OAI21xp33_ASAP7_75t_SL g3978 ( 
.A1(n_3932),
.A2(n_821),
.B(n_822),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3927),
.B(n_823),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3944),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3920),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3935),
.B(n_824),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3943),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3898),
.Y(n_3984)
);

OR2x2_ASAP7_75t_L g3985 ( 
.A(n_3902),
.B(n_825),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3908),
.B(n_826),
.Y(n_3986)
);

OAI322xp33_ASAP7_75t_L g3987 ( 
.A1(n_3931),
.A2(n_3911),
.A3(n_3918),
.B1(n_3913),
.B2(n_3914),
.C1(n_3942),
.C2(n_3940),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3904),
.B(n_828),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3928),
.B(n_831),
.Y(n_3989)
);

INVxp67_ASAP7_75t_L g3990 ( 
.A(n_3923),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3945),
.Y(n_3991)
);

AOI221x1_ASAP7_75t_SL g3992 ( 
.A1(n_3919),
.A2(n_834),
.B1(n_832),
.B2(n_833),
.C(n_835),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3922),
.B(n_835),
.Y(n_3993)
);

INVxp67_ASAP7_75t_L g3994 ( 
.A(n_3890),
.Y(n_3994)
);

OAI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3930),
.A2(n_838),
.B1(n_836),
.B2(n_837),
.Y(n_3995)
);

NOR2x1_ASAP7_75t_L g3996 ( 
.A(n_3941),
.B(n_836),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3939),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3917),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3924),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3912),
.B(n_837),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3886),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3886),
.Y(n_4002)
);

OAI221xp5_ASAP7_75t_L g4003 ( 
.A1(n_3946),
.A2(n_840),
.B1(n_838),
.B2(n_839),
.C(n_841),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3952),
.B(n_839),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3912),
.B(n_842),
.Y(n_4005)
);

OAI21xp5_ASAP7_75t_SL g4006 ( 
.A1(n_3946),
.A2(n_1346),
.B(n_1345),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3886),
.Y(n_4007)
);

OAI22xp33_ASAP7_75t_SL g4008 ( 
.A1(n_3912),
.A2(n_1348),
.B1(n_1349),
.B2(n_1347),
.Y(n_4008)
);

OAI21xp33_ASAP7_75t_L g4009 ( 
.A1(n_3889),
.A2(n_843),
.B(n_844),
.Y(n_4009)
);

OAI221xp5_ASAP7_75t_L g4010 ( 
.A1(n_3946),
.A2(n_846),
.B1(n_844),
.B2(n_845),
.C(n_847),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3886),
.Y(n_4011)
);

OAI211xp5_ASAP7_75t_SL g4012 ( 
.A1(n_3889),
.A2(n_851),
.B(n_848),
.C(n_849),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3912),
.B(n_848),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3886),
.Y(n_4014)
);

HB1xp67_ASAP7_75t_L g4015 ( 
.A(n_3949),
.Y(n_4015)
);

OAI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3915),
.A2(n_856),
.B1(n_854),
.B2(n_855),
.Y(n_4016)
);

AOI221xp5_ASAP7_75t_L g4017 ( 
.A1(n_3909),
.A2(n_867),
.B1(n_874),
.B2(n_859),
.C(n_855),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3886),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3952),
.B(n_857),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3886),
.Y(n_4020)
);

NOR2xp33_ASAP7_75t_L g4021 ( 
.A(n_3889),
.B(n_860),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3912),
.B(n_861),
.Y(n_4022)
);

INVxp33_ASAP7_75t_L g4023 ( 
.A(n_3947),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3915),
.A2(n_865),
.B1(n_863),
.B2(n_864),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3912),
.B(n_866),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3886),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3952),
.B(n_866),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3912),
.B(n_868),
.Y(n_4028)
);

AOI221xp5_ASAP7_75t_L g4029 ( 
.A1(n_3909),
.A2(n_882),
.B1(n_890),
.B2(n_877),
.C(n_869),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3952),
.B(n_871),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3912),
.B(n_873),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3886),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3912),
.B(n_873),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3886),
.Y(n_4034)
);

NAND2xp33_ASAP7_75t_L g4035 ( 
.A(n_3951),
.B(n_876),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3912),
.B(n_878),
.Y(n_4036)
);

INVxp67_ASAP7_75t_L g4037 ( 
.A(n_4015),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3953),
.Y(n_4038)
);

AOI22xp33_ASAP7_75t_SL g4039 ( 
.A1(n_3999),
.A2(n_883),
.B1(n_881),
.B2(n_882),
.Y(n_4039)
);

A2O1A1Ixp33_ASAP7_75t_L g4040 ( 
.A1(n_3992),
.A2(n_884),
.B(n_881),
.C(n_883),
.Y(n_4040)
);

AOI21xp33_ASAP7_75t_L g4041 ( 
.A1(n_4023),
.A2(n_3965),
.B(n_3961),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3954),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_SL g4043 ( 
.A(n_4008),
.B(n_885),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_4000),
.Y(n_4044)
);

AOI22xp5_ASAP7_75t_L g4045 ( 
.A1(n_3959),
.A2(n_1339),
.B1(n_1340),
.B2(n_1338),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_SL g4046 ( 
.A(n_3978),
.B(n_888),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_4005),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_4013),
.Y(n_4048)
);

NOR2xp33_ASAP7_75t_L g4049 ( 
.A(n_4022),
.B(n_891),
.Y(n_4049)
);

OR2x2_ASAP7_75t_L g4050 ( 
.A(n_4025),
.B(n_893),
.Y(n_4050)
);

AOI22xp5_ASAP7_75t_L g4051 ( 
.A1(n_3955),
.A2(n_3966),
.B1(n_3997),
.B2(n_4016),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_4028),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3960),
.B(n_894),
.Y(n_4053)
);

INVx1_ASAP7_75t_SL g4054 ( 
.A(n_3973),
.Y(n_4054)
);

AOI222xp33_ASAP7_75t_L g4055 ( 
.A1(n_3990),
.A2(n_3998),
.B1(n_3994),
.B2(n_4024),
.C1(n_4029),
.C2(n_4017),
.Y(n_4055)
);

AOI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_4006),
.A2(n_1343),
.B1(n_1346),
.B2(n_1340),
.Y(n_4056)
);

AOI221xp5_ASAP7_75t_L g4057 ( 
.A1(n_3987),
.A2(n_1357),
.B1(n_1361),
.B2(n_1354),
.C(n_1350),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_4031),
.Y(n_4058)
);

AOI21xp5_ASAP7_75t_L g4059 ( 
.A1(n_4035),
.A2(n_898),
.B(n_899),
.Y(n_4059)
);

OAI322xp33_ASAP7_75t_SL g4060 ( 
.A1(n_3956),
.A2(n_905),
.A3(n_904),
.B1(n_902),
.B2(n_900),
.C1(n_901),
.C2(n_903),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_4033),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_4003),
.A2(n_908),
.B1(n_906),
.B2(n_907),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_3967),
.B(n_907),
.Y(n_4063)
);

OAI211xp5_ASAP7_75t_SL g4064 ( 
.A1(n_3977),
.A2(n_910),
.B(n_908),
.C(n_909),
.Y(n_4064)
);

XOR2xp5_ASAP7_75t_L g4065 ( 
.A(n_3970),
.B(n_909),
.Y(n_4065)
);

AOI21xp33_ASAP7_75t_L g4066 ( 
.A1(n_3980),
.A2(n_910),
.B(n_911),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_4036),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_4004),
.Y(n_4068)
);

A2O1A1Ixp33_ASAP7_75t_L g4069 ( 
.A1(n_4012),
.A2(n_914),
.B(n_911),
.C(n_913),
.Y(n_4069)
);

OR2x2_ASAP7_75t_L g4070 ( 
.A(n_3958),
.B(n_916),
.Y(n_4070)
);

NOR2xp33_ASAP7_75t_L g4071 ( 
.A(n_4009),
.B(n_917),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_4021),
.B(n_921),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_4019),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_4027),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3983),
.B(n_4030),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3975),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_3985),
.Y(n_4077)
);

AOI32xp33_ASAP7_75t_L g4078 ( 
.A1(n_3996),
.A2(n_924),
.A3(n_922),
.B1(n_923),
.B2(n_925),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3962),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3982),
.Y(n_4080)
);

NAND2x1_ASAP7_75t_SL g4081 ( 
.A(n_3986),
.B(n_924),
.Y(n_4081)
);

NOR2xp33_ASAP7_75t_L g4082 ( 
.A(n_4010),
.B(n_926),
.Y(n_4082)
);

INVx1_ASAP7_75t_SL g4083 ( 
.A(n_3974),
.Y(n_4083)
);

OAI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_3957),
.A2(n_929),
.B1(n_927),
.B2(n_928),
.Y(n_4084)
);

AOI22xp5_ASAP7_75t_L g4085 ( 
.A1(n_3969),
.A2(n_1335),
.B1(n_1337),
.B2(n_1334),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3979),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4001),
.Y(n_4087)
);

AOI211xp5_ASAP7_75t_L g4088 ( 
.A1(n_3995),
.A2(n_940),
.B(n_944),
.C(n_930),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_4002),
.Y(n_4089)
);

OAI21xp33_ASAP7_75t_L g4090 ( 
.A1(n_3984),
.A2(n_931),
.B(n_932),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4007),
.Y(n_4091)
);

AOI322xp5_ASAP7_75t_L g4092 ( 
.A1(n_3968),
.A2(n_940),
.A3(n_939),
.B1(n_936),
.B2(n_933),
.C1(n_935),
.C2(n_938),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4011),
.Y(n_4093)
);

AOI21xp33_ASAP7_75t_L g4094 ( 
.A1(n_3971),
.A2(n_935),
.B(n_936),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4014),
.Y(n_4095)
);

OAI21xp33_ASAP7_75t_SL g4096 ( 
.A1(n_4018),
.A2(n_938),
.B(n_941),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4020),
.Y(n_4097)
);

OR2x2_ASAP7_75t_L g4098 ( 
.A(n_4026),
.B(n_941),
.Y(n_4098)
);

OAI221xp5_ASAP7_75t_L g4099 ( 
.A1(n_4057),
.A2(n_4034),
.B1(n_4032),
.B2(n_3981),
.C(n_3991),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_4054),
.B(n_3976),
.Y(n_4100)
);

OAI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_4040),
.A2(n_3972),
.B(n_3988),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_4046),
.A2(n_3993),
.B(n_3989),
.Y(n_4102)
);

OAI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_4037),
.A2(n_3964),
.B(n_3963),
.Y(n_4103)
);

AOI21xp33_ASAP7_75t_SL g4104 ( 
.A1(n_4043),
.A2(n_943),
.B(n_942),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4075),
.B(n_948),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_4053),
.B(n_950),
.Y(n_4106)
);

AOI221xp5_ASAP7_75t_L g4107 ( 
.A1(n_4060),
.A2(n_954),
.B1(n_952),
.B2(n_953),
.C(n_955),
.Y(n_4107)
);

AOI311xp33_ASAP7_75t_L g4108 ( 
.A1(n_4042),
.A2(n_4044),
.A3(n_4052),
.B(n_4048),
.C(n_4047),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_SL g4109 ( 
.A1(n_4083),
.A2(n_961),
.B1(n_956),
.B2(n_959),
.Y(n_4109)
);

OAI221xp5_ASAP7_75t_L g4110 ( 
.A1(n_4065),
.A2(n_964),
.B1(n_962),
.B2(n_963),
.C(n_965),
.Y(n_4110)
);

OAI221xp5_ASAP7_75t_L g4111 ( 
.A1(n_4078),
.A2(n_966),
.B1(n_964),
.B2(n_965),
.C(n_967),
.Y(n_4111)
);

NOR4xp25_ASAP7_75t_L g4112 ( 
.A(n_4087),
.B(n_968),
.C(n_966),
.D(n_967),
.Y(n_4112)
);

NOR4xp25_ASAP7_75t_L g4113 ( 
.A(n_4089),
.B(n_971),
.C(n_969),
.D(n_970),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4063),
.Y(n_4114)
);

INVx1_ASAP7_75t_SL g4115 ( 
.A(n_4050),
.Y(n_4115)
);

A2O1A1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_4069),
.A2(n_4096),
.B(n_4082),
.C(n_4059),
.Y(n_4116)
);

NAND3xp33_ASAP7_75t_SL g4117 ( 
.A(n_4088),
.B(n_976),
.C(n_975),
.Y(n_4117)
);

AOI211xp5_ASAP7_75t_L g4118 ( 
.A1(n_4064),
.A2(n_1324),
.B(n_1325),
.C(n_1323),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_L g4119 ( 
.A(n_4090),
.B(n_977),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_4098),
.Y(n_4120)
);

OAI21xp33_ASAP7_75t_SL g4121 ( 
.A1(n_4068),
.A2(n_978),
.B(n_980),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_4039),
.B(n_981),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_4080),
.B(n_984),
.Y(n_4123)
);

OAI211xp5_ASAP7_75t_L g4124 ( 
.A1(n_4045),
.A2(n_987),
.B(n_985),
.C(n_986),
.Y(n_4124)
);

OAI21xp5_ASAP7_75t_SL g4125 ( 
.A1(n_4058),
.A2(n_986),
.B(n_987),
.Y(n_4125)
);

NAND3xp33_ASAP7_75t_L g4126 ( 
.A(n_4091),
.B(n_988),
.C(n_989),
.Y(n_4126)
);

OAI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_4056),
.A2(n_992),
.B1(n_990),
.B2(n_991),
.Y(n_4127)
);

OAI221xp5_ASAP7_75t_SL g4128 ( 
.A1(n_4061),
.A2(n_1329),
.B1(n_1330),
.B2(n_1328),
.C(n_1327),
.Y(n_4128)
);

NAND4xp25_ASAP7_75t_L g4129 ( 
.A(n_4067),
.B(n_996),
.C(n_994),
.D(n_995),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_SL g4130 ( 
.A(n_4076),
.B(n_996),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_4073),
.B(n_997),
.Y(n_4131)
);

NAND4xp25_ASAP7_75t_L g4132 ( 
.A(n_4074),
.B(n_1001),
.C(n_998),
.D(n_999),
.Y(n_4132)
);

XNOR2x1_ASAP7_75t_L g4133 ( 
.A(n_4062),
.B(n_1002),
.Y(n_4133)
);

AOI21xp33_ASAP7_75t_SL g4134 ( 
.A1(n_4077),
.A2(n_1003),
.B(n_1002),
.Y(n_4134)
);

AOI21xp5_ASAP7_75t_L g4135 ( 
.A1(n_4072),
.A2(n_1005),
.B(n_1007),
.Y(n_4135)
);

AOI221xp5_ASAP7_75t_L g4136 ( 
.A1(n_4093),
.A2(n_4095),
.B1(n_4097),
.B2(n_4084),
.C(n_4066),
.Y(n_4136)
);

AOI21xp33_ASAP7_75t_SL g4137 ( 
.A1(n_4070),
.A2(n_1011),
.B(n_1010),
.Y(n_4137)
);

NAND4xp25_ASAP7_75t_L g4138 ( 
.A(n_4079),
.B(n_1014),
.C(n_1012),
.D(n_1013),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_4094),
.A2(n_4086),
.B(n_4049),
.Y(n_4139)
);

AOI221xp5_ASAP7_75t_L g4140 ( 
.A1(n_4071),
.A2(n_1021),
.B1(n_1019),
.B2(n_1020),
.C(n_1022),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4085),
.Y(n_4141)
);

OAI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_4092),
.A2(n_1023),
.B(n_1024),
.Y(n_4142)
);

NOR3xp33_ASAP7_75t_L g4143 ( 
.A(n_4041),
.B(n_1026),
.C(n_1027),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_4054),
.B(n_1028),
.Y(n_4144)
);

NAND4xp25_ASAP7_75t_L g4145 ( 
.A(n_4055),
.B(n_1031),
.C(n_1029),
.D(n_1030),
.Y(n_4145)
);

NAND3xp33_ASAP7_75t_L g4146 ( 
.A(n_4057),
.B(n_1032),
.C(n_1033),
.Y(n_4146)
);

AOI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_4046),
.A2(n_1034),
.B(n_1035),
.Y(n_4147)
);

OAI21xp33_ASAP7_75t_SL g4148 ( 
.A1(n_4038),
.A2(n_1034),
.B(n_1035),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4081),
.Y(n_4149)
);

NOR3xp33_ASAP7_75t_L g4150 ( 
.A(n_4041),
.B(n_1036),
.C(n_1037),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4054),
.B(n_1037),
.Y(n_4151)
);

NOR3xp33_ASAP7_75t_L g4152 ( 
.A(n_4041),
.B(n_1040),
.C(n_1041),
.Y(n_4152)
);

OAI21xp5_ASAP7_75t_SL g4153 ( 
.A1(n_4051),
.A2(n_1046),
.B(n_1047),
.Y(n_4153)
);

NAND3xp33_ASAP7_75t_SL g4154 ( 
.A(n_4054),
.B(n_1052),
.C(n_1051),
.Y(n_4154)
);

NOR2xp33_ASAP7_75t_L g4155 ( 
.A(n_4054),
.B(n_1050),
.Y(n_4155)
);

XOR2x2_ASAP7_75t_L g4156 ( 
.A(n_4081),
.B(n_1051),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_SL g4157 ( 
.A(n_4038),
.B(n_1052),
.Y(n_4157)
);

NAND4xp25_ASAP7_75t_L g4158 ( 
.A(n_4055),
.B(n_1059),
.C(n_1057),
.D(n_1058),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_4155),
.A2(n_1061),
.B1(n_1059),
.B2(n_1060),
.Y(n_4159)
);

AOI322xp5_ASAP7_75t_L g4160 ( 
.A1(n_4107),
.A2(n_1069),
.A3(n_1068),
.B1(n_1066),
.B2(n_1064),
.C1(n_1065),
.C2(n_1067),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4156),
.Y(n_4161)
);

OAI322xp33_ASAP7_75t_SL g4162 ( 
.A1(n_4100),
.A2(n_1081),
.A3(n_1080),
.B1(n_1078),
.B2(n_1075),
.C1(n_1077),
.C2(n_1079),
.Y(n_4162)
);

AOI221xp5_ASAP7_75t_L g4163 ( 
.A1(n_4145),
.A2(n_1084),
.B1(n_1086),
.B2(n_1083),
.C(n_1085),
.Y(n_4163)
);

AOI221xp5_ASAP7_75t_L g4164 ( 
.A1(n_4158),
.A2(n_1091),
.B1(n_1093),
.B2(n_1090),
.C(n_1092),
.Y(n_4164)
);

AOI221xp5_ASAP7_75t_L g4165 ( 
.A1(n_4142),
.A2(n_1096),
.B1(n_1098),
.B2(n_1095),
.C(n_1097),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_4149),
.B(n_1094),
.Y(n_4166)
);

AOI321xp33_ASAP7_75t_L g4167 ( 
.A1(n_4108),
.A2(n_1098),
.A3(n_1100),
.B1(n_1096),
.B2(n_1097),
.C(n_1099),
.Y(n_4167)
);

AOI322xp5_ASAP7_75t_L g4168 ( 
.A1(n_4117),
.A2(n_4141),
.A3(n_4154),
.B1(n_4136),
.B2(n_4150),
.C1(n_4143),
.C2(n_4152),
.Y(n_4168)
);

OAI221xp5_ASAP7_75t_L g4169 ( 
.A1(n_4153),
.A2(n_1104),
.B1(n_1102),
.B2(n_1103),
.C(n_1105),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_4105),
.B(n_1104),
.Y(n_4170)
);

OAI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_4146),
.A2(n_1110),
.B1(n_1106),
.B2(n_1109),
.Y(n_4171)
);

AOI31xp33_ASAP7_75t_L g4172 ( 
.A1(n_4104),
.A2(n_1115),
.A3(n_1116),
.B(n_1114),
.Y(n_4172)
);

OAI221xp5_ASAP7_75t_L g4173 ( 
.A1(n_4101),
.A2(n_4103),
.B1(n_4116),
.B2(n_4099),
.C(n_4148),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4144),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4112),
.B(n_1112),
.Y(n_4175)
);

BUFx2_ASAP7_75t_L g4176 ( 
.A(n_4121),
.Y(n_4176)
);

AOI221xp5_ASAP7_75t_L g4177 ( 
.A1(n_4113),
.A2(n_1119),
.B1(n_1121),
.B2(n_1118),
.C(n_1120),
.Y(n_4177)
);

OR2x2_ASAP7_75t_L g4178 ( 
.A(n_4151),
.B(n_1122),
.Y(n_4178)
);

NAND4xp25_ASAP7_75t_L g4179 ( 
.A(n_4102),
.B(n_4139),
.C(n_4114),
.D(n_4115),
.Y(n_4179)
);

NOR2x1p5_ASAP7_75t_L g4180 ( 
.A(n_4122),
.B(n_4120),
.Y(n_4180)
);

BUFx3_ASAP7_75t_L g4181 ( 
.A(n_4106),
.Y(n_4181)
);

OAI22xp5_ASAP7_75t_L g4182 ( 
.A1(n_4111),
.A2(n_4118),
.B1(n_4110),
.B2(n_4109),
.Y(n_4182)
);

AOI31xp33_ASAP7_75t_L g4183 ( 
.A1(n_4147),
.A2(n_1125),
.A3(n_1127),
.B(n_1124),
.Y(n_4183)
);

AOI211xp5_ASAP7_75t_SL g4184 ( 
.A1(n_4124),
.A2(n_1134),
.B(n_1131),
.C(n_1133),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_SL g4185 ( 
.A(n_4167),
.B(n_4137),
.Y(n_4185)
);

OAI21xp33_ASAP7_75t_L g4186 ( 
.A1(n_4168),
.A2(n_4133),
.B(n_4131),
.Y(n_4186)
);

OAI21xp33_ASAP7_75t_L g4187 ( 
.A1(n_4179),
.A2(n_4123),
.B(n_4119),
.Y(n_4187)
);

AOI21x1_ASAP7_75t_L g4188 ( 
.A1(n_4176),
.A2(n_4157),
.B(n_4130),
.Y(n_4188)
);

O2A1O1Ixp33_ASAP7_75t_L g4189 ( 
.A1(n_4175),
.A2(n_4134),
.B(n_4128),
.C(n_4125),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_SL g4190 ( 
.A1(n_4173),
.A2(n_4127),
.B1(n_4126),
.B2(n_4135),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_4178),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4184),
.B(n_4160),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4170),
.Y(n_4193)
);

NOR2x1p5_ASAP7_75t_L g4194 ( 
.A(n_4161),
.B(n_4132),
.Y(n_4194)
);

AOI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_4182),
.A2(n_4140),
.B1(n_4129),
.B2(n_4138),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4172),
.Y(n_4196)
);

AOI322xp5_ASAP7_75t_L g4197 ( 
.A1(n_4165),
.A2(n_1139),
.A3(n_1138),
.B1(n_1136),
.B2(n_1134),
.C1(n_1135),
.C2(n_1137),
.Y(n_4197)
);

AOI22xp5_ASAP7_75t_L g4198 ( 
.A1(n_4180),
.A2(n_1142),
.B1(n_1140),
.B2(n_1141),
.Y(n_4198)
);

NOR3xp33_ASAP7_75t_L g4199 ( 
.A(n_4171),
.B(n_1148),
.C(n_1149),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4183),
.Y(n_4200)
);

AOI221xp5_ASAP7_75t_L g4201 ( 
.A1(n_4162),
.A2(n_1153),
.B1(n_1151),
.B2(n_1152),
.C(n_1154),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_4181),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4166),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4159),
.Y(n_4204)
);

OAI22xp5_ASAP7_75t_L g4205 ( 
.A1(n_4169),
.A2(n_1159),
.B1(n_1157),
.B2(n_1158),
.Y(n_4205)
);

OAI211xp5_ASAP7_75t_SL g4206 ( 
.A1(n_4174),
.A2(n_1162),
.B(n_1160),
.C(n_1161),
.Y(n_4206)
);

NAND4xp25_ASAP7_75t_SL g4207 ( 
.A(n_4201),
.B(n_4177),
.C(n_4163),
.D(n_4164),
.Y(n_4207)
);

OAI21xp33_ASAP7_75t_SL g4208 ( 
.A1(n_4185),
.A2(n_4192),
.B(n_4194),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4188),
.Y(n_4209)
);

OAI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_4195),
.A2(n_4190),
.B1(n_4196),
.B2(n_4198),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_4189),
.A2(n_1164),
.B(n_1165),
.Y(n_4211)
);

OAI21xp33_ASAP7_75t_SL g4212 ( 
.A1(n_4200),
.A2(n_1166),
.B(n_1167),
.Y(n_4212)
);

NOR3xp33_ASAP7_75t_L g4213 ( 
.A(n_4186),
.B(n_1168),
.C(n_1169),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4202),
.B(n_4203),
.Y(n_4214)
);

AOI221xp5_ASAP7_75t_L g4215 ( 
.A1(n_4187),
.A2(n_1175),
.B1(n_1172),
.B2(n_1173),
.C(n_1176),
.Y(n_4215)
);

AOI21xp33_ASAP7_75t_L g4216 ( 
.A1(n_4204),
.A2(n_1173),
.B(n_1175),
.Y(n_4216)
);

AND2x4_ASAP7_75t_L g4217 ( 
.A(n_4191),
.B(n_1177),
.Y(n_4217)
);

OAI21xp33_ASAP7_75t_L g4218 ( 
.A1(n_4193),
.A2(n_4199),
.B(n_4197),
.Y(n_4218)
);

NOR2x1_ASAP7_75t_L g4219 ( 
.A(n_4209),
.B(n_4206),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_L g4220 ( 
.A(n_4212),
.B(n_4205),
.Y(n_4220)
);

HB1xp67_ASAP7_75t_L g4221 ( 
.A(n_4217),
.Y(n_4221)
);

AOI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4207),
.A2(n_1180),
.B1(n_1178),
.B2(n_1179),
.Y(n_4222)
);

AOI22xp5_ASAP7_75t_L g4223 ( 
.A1(n_4208),
.A2(n_1183),
.B1(n_1181),
.B2(n_1182),
.Y(n_4223)
);

BUFx6f_ASAP7_75t_L g4224 ( 
.A(n_4214),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4213),
.B(n_1183),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4221),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4224),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4222),
.Y(n_4228)
);

XNOR2xp5_ASAP7_75t_L g4229 ( 
.A(n_4223),
.B(n_4210),
.Y(n_4229)
);

NAND4xp75_ASAP7_75t_L g4230 ( 
.A(n_4219),
.B(n_4211),
.C(n_4215),
.D(n_4216),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4220),
.Y(n_4231)
);

AND2x2_ASAP7_75t_L g4232 ( 
.A(n_4225),
.B(n_4218),
.Y(n_4232)
);

NOR3xp33_ASAP7_75t_L g4233 ( 
.A(n_4226),
.B(n_1184),
.C(n_1185),
.Y(n_4233)
);

XNOR2xp5_ASAP7_75t_L g4234 ( 
.A(n_4229),
.B(n_1185),
.Y(n_4234)
);

AOI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_4231),
.A2(n_1190),
.B1(n_1188),
.B2(n_1189),
.Y(n_4235)
);

OAI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4227),
.A2(n_1193),
.B1(n_1191),
.B2(n_1192),
.Y(n_4236)
);

NAND5xp2_ASAP7_75t_L g4237 ( 
.A(n_4228),
.B(n_1197),
.C(n_1195),
.D(n_1196),
.E(n_1198),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4234),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_4237),
.B(n_4230),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_4238),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_4239),
.B(n_4233),
.Y(n_4241)
);

CKINVDCx5p33_ASAP7_75t_R g4242 ( 
.A(n_4240),
.Y(n_4242)
);

XNOR2x1_ASAP7_75t_L g4243 ( 
.A(n_4242),
.B(n_4232),
.Y(n_4243)
);

OAI22xp5_ASAP7_75t_L g4244 ( 
.A1(n_4243),
.A2(n_4241),
.B1(n_4235),
.B2(n_4236),
.Y(n_4244)
);

XNOR2x1_ASAP7_75t_L g4245 ( 
.A(n_4244),
.B(n_1196),
.Y(n_4245)
);

OR2x2_ASAP7_75t_L g4246 ( 
.A(n_4245),
.B(n_1197),
.Y(n_4246)
);

XNOR2xp5_ASAP7_75t_L g4247 ( 
.A(n_4246),
.B(n_1199),
.Y(n_4247)
);

AOI222xp33_ASAP7_75t_L g4248 ( 
.A1(n_4247),
.A2(n_1203),
.B1(n_1205),
.B2(n_1200),
.C1(n_1202),
.C2(n_1204),
.Y(n_4248)
);

OA21x2_ASAP7_75t_L g4249 ( 
.A1(n_4248),
.A2(n_1206),
.B(n_1208),
.Y(n_4249)
);

AOI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_4249),
.A2(n_1209),
.B(n_1210),
.Y(n_4250)
);

AOI211xp5_ASAP7_75t_L g4251 ( 
.A1(n_4250),
.A2(n_1319),
.B(n_1211),
.C(n_1210),
.Y(n_4251)
);


endmodule