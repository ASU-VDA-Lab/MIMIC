module real_jpeg_155_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_1),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_1),
.A2(n_24),
.B1(n_31),
.B2(n_43),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_21),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_62),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_3),
.B(n_36),
.C(n_54),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_24),
.B1(n_29),
.B2(n_31),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_3),
.B(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_58),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_24),
.B1(n_31),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_36),
.B1(n_44),
.B2(n_51),
.Y(n_99)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_36),
.B1(n_44),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_9),
.A2(n_24),
.B1(n_31),
.B2(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_9),
.A2(n_36),
.B1(n_44),
.B2(n_65),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_21),
.B1(n_22),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_24),
.B1(n_31),
.B2(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_10),
.A2(n_36),
.B1(n_44),
.B2(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_12),
.A2(n_36),
.B1(n_44),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_90),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_81),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_81),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_59),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_48),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_33),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.A3(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_32),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_21),
.A2(n_22),
.B1(n_74),
.B2(n_76),
.Y(n_73)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_31),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

AO22x2_ASAP7_75t_SL g62 ( 
.A1(n_24),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_107),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_29),
.A2(n_35),
.B1(n_39),
.B2(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B1(n_41),
.B2(n_45),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_34),
.A2(n_38),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_35),
.A2(n_39),
.B1(n_46),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_35),
.A2(n_39),
.B1(n_42),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_35),
.A2(n_39),
.B1(n_119),
.B2(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_36),
.B(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_56),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_58),
.B1(n_89),
.B2(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_52),
.A2(n_58),
.B1(n_96),
.B2(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_69),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_64),
.B1(n_66),
.B2(n_84),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_77),
.B2(n_80),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_74),
.Y(n_76)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.C(n_86),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_86),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_102),
.B(n_132),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_100),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_97),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_113),
.B(n_131),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_125),
.B(n_130),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_120),
.B(n_124),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_122),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_129),
.Y(n_130)
);


endmodule