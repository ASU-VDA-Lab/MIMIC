module fake_netlist_5_228_n_811 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_811);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_811;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_753;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_804;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_95),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_170),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_82),
.B(n_140),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_84),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_9),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_52),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_29),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_50),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_35),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_92),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_12),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_11),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_98),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_57),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_22),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_32),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_128),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_141),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_73),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_33),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_66),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_1),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_94),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_100),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_126),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_37),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_142),
.B(n_7),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_40),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_80),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_67),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_106),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_111),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_18),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_77),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_169),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_0),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_215),
.B(n_0),
.Y(n_244)
);

AOI22x1_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

BUFx8_ASAP7_75t_SL g249 ( 
.A(n_234),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_19),
.Y(n_250)
);

BUFx8_ASAP7_75t_SL g251 ( 
.A(n_198),
.Y(n_251)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_20),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_198),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_181),
.B(n_2),
.Y(n_254)
);

OAI22x1_ASAP7_75t_L g255 ( 
.A1(n_182),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx11_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_6),
.Y(n_260)
);

OAI22x1_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_209),
.B1(n_200),
.B2(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_196),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_196),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_173),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

OAI22x1_ASAP7_75t_SL g272 ( 
.A1(n_175),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_188),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

OA21x2_ASAP7_75t_L g275 ( 
.A1(n_193),
.A2(n_201),
.B(n_195),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_179),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_204),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_180),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_194),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_183),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_222),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_184),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_214),
.B(n_8),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_178),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_189),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_266),
.B(n_192),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_253),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_276),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_291),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_251),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_291),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_248),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_287),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_251),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_R g306 ( 
.A(n_264),
.B(n_197),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_256),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

AND3x2_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_232),
.C(n_228),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_258),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_249),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_177),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_289),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_249),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_263),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_257),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_R g329 ( 
.A(n_290),
.B(n_203),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_246),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_R g332 ( 
.A(n_267),
.B(n_206),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_283),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_246),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_243),
.B(n_269),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_283),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_286),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_282),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_262),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_282),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_259),
.C(n_269),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_333),
.B(n_263),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_292),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_322),
.B(n_263),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_280),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_298),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_275),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_254),
.B1(n_244),
.B2(n_288),
.Y(n_356)
);

AO221x1_ASAP7_75t_L g357 ( 
.A1(n_342),
.A2(n_255),
.B1(n_241),
.B2(n_233),
.C(n_240),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_263),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_299),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_340),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_288),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_315),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_332),
.B(n_243),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_339),
.B(n_260),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_303),
.B(n_317),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_280),
.Y(n_372)
);

NAND2xp33_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_250),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_250),
.Y(n_374)
);

NOR3xp33_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_259),
.C(n_265),
.Y(n_375)
);

AO221x1_ASAP7_75t_L g376 ( 
.A1(n_321),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.C(n_277),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_280),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_311),
.B(n_278),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_311),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_250),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_250),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_274),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_278),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_274),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_314),
.B(n_207),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_281),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_293),
.B(n_277),
.Y(n_393)
);

AO221x1_ASAP7_75t_L g394 ( 
.A1(n_328),
.A2(n_285),
.B1(n_284),
.B2(n_281),
.C(n_272),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_300),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_296),
.B(n_281),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_309),
.B(n_284),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_304),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_320),
.B(n_208),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_210),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_306),
.A2(n_261),
.B1(n_212),
.B2(n_229),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_294),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_333),
.B(n_217),
.Y(n_405)
);

NOR3xp33_ASAP7_75t_L g406 ( 
.A(n_295),
.B(n_252),
.C(n_218),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_391),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_345),
.B(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_355),
.B(n_284),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_355),
.A2(n_357),
.B1(n_373),
.B2(n_356),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_363),
.A2(n_245),
.B1(n_219),
.B2(n_237),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_374),
.A2(n_285),
.B1(n_242),
.B2(n_235),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_396),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_366),
.B(n_285),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

OR2x4_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_10),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_225),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_226),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

NAND2x1p5_ASAP7_75t_L g426 ( 
.A(n_371),
.B(n_23),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_348),
.B(n_230),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_10),
.Y(n_428)
);

BUFx12f_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_11),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_359),
.B(n_403),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_351),
.B(n_393),
.Y(n_435)
);

NOR2x1p5_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_13),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_24),
.Y(n_437)
);

AO21x1_ASAP7_75t_L g438 ( 
.A1(n_385),
.A2(n_14),
.B(n_15),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_380),
.Y(n_440)
);

BUFx8_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_388),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_388),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_367),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_384),
.A2(n_97),
.B(n_171),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_376),
.A2(n_406),
.B1(n_344),
.B2(n_375),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_25),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_362),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_372),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_379),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_26),
.Y(n_456)
);

NAND2x1p5_ASAP7_75t_L g457 ( 
.A(n_347),
.B(n_27),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_28),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

BUFx8_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_15),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_377),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_402),
.A2(n_16),
.B1(n_17),
.B2(n_30),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_379),
.B(n_31),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_397),
.A2(n_16),
.B1(n_17),
.B2(n_34),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_431),
.A2(n_395),
.B(n_38),
.C(n_39),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_415),
.B(n_36),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_SL g471 ( 
.A(n_415),
.B(n_41),
.C(n_43),
.Y(n_471)
);

O2A1O1Ixp5_ASAP7_75t_L g472 ( 
.A1(n_433),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_424),
.A2(n_410),
.B(n_416),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_47),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_432),
.B(n_48),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_418),
.A2(n_49),
.B(n_51),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_54),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_55),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_56),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_59),
.Y(n_482)
);

NOR3xp33_ASAP7_75t_SL g483 ( 
.A(n_413),
.B(n_60),
.C(n_61),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_444),
.B(n_62),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_429),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_65),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_453),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_412),
.A2(n_68),
.B(n_69),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_70),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_409),
.A2(n_71),
.B(n_72),
.C(n_74),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_407),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_454),
.A2(n_79),
.B(n_83),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_435),
.B(n_85),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_428),
.A2(n_89),
.B(n_90),
.C(n_93),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_408),
.B(n_99),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_465),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_423),
.A2(n_466),
.B1(n_414),
.B2(n_451),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_427),
.B(n_101),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_419),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_462),
.A2(n_108),
.B(n_109),
.C(n_110),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_423),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_115),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_450),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_437),
.A2(n_116),
.B(n_117),
.C(n_119),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_460),
.B(n_120),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_425),
.A2(n_124),
.B(n_127),
.C(n_131),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_465),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_439),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_460),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_450),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_455),
.B(n_139),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_491),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_487),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_518),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_491),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_474),
.A2(n_459),
.B(n_456),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_514),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_473),
.B(n_407),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_480),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_501),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_440),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_504),
.A2(n_438),
.B1(n_436),
.B2(n_426),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_503),
.Y(n_534)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_481),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_458),
.Y(n_537)
);

NOR2x1_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_467),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

AO21x2_ASAP7_75t_L g540 ( 
.A1(n_489),
.A2(n_452),
.B(n_459),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_478),
.B(n_463),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_482),
.Y(n_543)
);

OA21x2_ASAP7_75t_L g544 ( 
.A1(n_497),
.A2(n_452),
.B(n_447),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_488),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_506),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_516),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_510),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_519),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_457),
.Y(n_551)
);

BUFx8_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_519),
.Y(n_553)
);

AOI22x1_ASAP7_75t_L g554 ( 
.A1(n_477),
.A2(n_468),
.B1(n_413),
.B2(n_461),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_502),
.A2(n_468),
.B(n_144),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_486),
.A2(n_143),
.B(n_145),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_509),
.Y(n_560)
);

OA21x2_ASAP7_75t_L g561 ( 
.A1(n_472),
.A2(n_148),
.B(n_149),
.Y(n_561)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_490),
.Y(n_562)
);

AOI22x1_ASAP7_75t_L g563 ( 
.A1(n_496),
.A2(n_461),
.B1(n_151),
.B2(n_152),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_469),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_499),
.A2(n_150),
.B(n_153),
.Y(n_565)
);

BUFx2_ASAP7_75t_SL g566 ( 
.A(n_512),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

INVx3_ASAP7_75t_SL g568 ( 
.A(n_534),
.Y(n_568)
);

INVx8_ASAP7_75t_L g569 ( 
.A(n_562),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_483),
.C(n_505),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_522),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_536),
.Y(n_572)
);

CKINVDCx11_ASAP7_75t_R g573 ( 
.A(n_534),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_536),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_530),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_547),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_560),
.B(n_476),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_547),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_527),
.B(n_470),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_539),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_545),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_548),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_537),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_530),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_551),
.A2(n_517),
.B1(n_508),
.B2(n_441),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_527),
.B(n_511),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_539),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_531),
.Y(n_590)
);

CKINVDCx11_ASAP7_75t_R g591 ( 
.A(n_529),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_554),
.A2(n_495),
.B1(n_507),
.B2(n_498),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_535),
.Y(n_593)
);

AO21x1_ASAP7_75t_SL g594 ( 
.A1(n_533),
.A2(n_493),
.B(n_513),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_541),
.B(n_441),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_535),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_527),
.B(n_154),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_532),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_523),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_556),
.B(n_160),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

CKINVDCx6p67_ASAP7_75t_R g602 ( 
.A(n_529),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_552),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_564),
.A2(n_172),
.B(n_163),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_564),
.A2(n_161),
.B1(n_165),
.B2(n_168),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_576),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_568),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_572),
.B(n_559),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_562),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_526),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_577),
.B(n_543),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_573),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_573),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_SL g617 ( 
.A(n_570),
.B(n_586),
.C(n_595),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_R g618 ( 
.A(n_571),
.B(n_551),
.Y(n_618)
);

AO31x2_ASAP7_75t_L g619 ( 
.A1(n_600),
.A2(n_559),
.A3(n_540),
.B(n_525),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_602),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_569),
.B(n_562),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_578),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_591),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_R g624 ( 
.A(n_607),
.B(n_561),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_575),
.Y(n_625)
);

AO21x2_ASAP7_75t_L g626 ( 
.A1(n_592),
.A2(n_525),
.B(n_540),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_591),
.Y(n_627)
);

NOR3xp33_ASAP7_75t_SL g628 ( 
.A(n_598),
.B(n_521),
.C(n_524),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_590),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_542),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_575),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_582),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_568),
.Y(n_633)
);

OAI21xp33_ASAP7_75t_L g634 ( 
.A1(n_608),
.A2(n_538),
.B(n_563),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_574),
.B(n_553),
.Y(n_635)
);

CKINVDCx11_ASAP7_75t_R g636 ( 
.A(n_583),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_585),
.B(n_566),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_603),
.B(n_553),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_569),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_585),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_581),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_567),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_603),
.B(n_549),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_604),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_608),
.A2(n_558),
.B1(n_566),
.B2(n_562),
.Y(n_646)
);

AND2x2_ASAP7_75t_SL g647 ( 
.A(n_587),
.B(n_561),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_604),
.B(n_549),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_SL g649 ( 
.A(n_598),
.B(n_558),
.C(n_528),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_582),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_599),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_528),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_528),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_605),
.B(n_555),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_609),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_612),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_632),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_612),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_629),
.B(n_584),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_639),
.B(n_582),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_622),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_648),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_617),
.B(n_582),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_642),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_635),
.B(n_555),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_645),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_653),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_653),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_647),
.B(n_557),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_625),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_631),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_611),
.B(n_589),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_618),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_632),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_614),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_654),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_626),
.B(n_557),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_654),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_654),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_641),
.B(n_557),
.Y(n_680)
);

AND2x6_ASAP7_75t_SL g681 ( 
.A(n_652),
.B(n_605),
.Y(n_681)
);

AND2x4_ASAP7_75t_SL g682 ( 
.A(n_650),
.B(n_589),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_651),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_638),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_611),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_619),
.B(n_565),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_SL g688 ( 
.A1(n_646),
.A2(n_592),
.B(n_565),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_634),
.A2(n_563),
.B1(n_594),
.B2(n_540),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_626),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_667),
.B(n_610),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_668),
.B(n_630),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_673),
.B(n_610),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_684),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_655),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_655),
.Y(n_696)
);

AOI221xp5_ASAP7_75t_SL g697 ( 
.A1(n_663),
.A2(n_646),
.B1(n_634),
.B2(n_637),
.C(n_633),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_689),
.B(n_628),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_662),
.B(n_613),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_675),
.B(n_619),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_686),
.B(n_619),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_664),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_664),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_661),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_688),
.B(n_612),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_660),
.B(n_613),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_681),
.B(n_636),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_678),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_659),
.B(n_615),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_666),
.B(n_616),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_670),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_656),
.B(n_627),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_670),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_685),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_680),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_700),
.B(n_678),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_694),
.B(n_676),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_708),
.B(n_676),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_695),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_695),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_692),
.B(n_679),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_693),
.B(n_679),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_694),
.B(n_669),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_706),
.B(n_679),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_702),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_701),
.B(n_669),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_715),
.B(n_676),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_714),
.B(n_685),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_696),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_699),
.B(n_665),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_696),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_711),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_708),
.B(n_665),
.Y(n_733)
);

OAI222xp33_ASAP7_75t_L g734 ( 
.A1(n_726),
.A2(n_698),
.B1(n_705),
.B2(n_691),
.C1(n_709),
.C2(n_710),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_726),
.B(n_723),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_725),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_732),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_723),
.B(n_704),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_732),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_719),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_719),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_L g742 ( 
.A1(n_716),
.A2(n_698),
.B(n_688),
.Y(n_742)
);

AOI211x1_ASAP7_75t_L g743 ( 
.A1(n_734),
.A2(n_722),
.B(n_721),
.C(n_728),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_742),
.A2(n_705),
.B1(n_649),
.B2(n_712),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_734),
.A2(n_707),
.B(n_697),
.C(n_735),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_738),
.A2(n_705),
.B1(n_658),
.B2(n_656),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_736),
.A2(n_707),
.B1(n_656),
.B2(n_658),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_745),
.B(n_730),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_744),
.A2(n_623),
.B(n_620),
.C(n_718),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_746),
.A2(n_747),
.B(n_728),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_743),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_SL g753 ( 
.A(n_744),
.B(n_658),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_751),
.B(n_739),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_SL g755 ( 
.A(n_750),
.B(n_658),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_752),
.Y(n_756)
);

OAI21xp33_ASAP7_75t_L g757 ( 
.A1(n_748),
.A2(n_717),
.B(n_733),
.Y(n_757)
);

AOI211x1_ASAP7_75t_L g758 ( 
.A1(n_756),
.A2(n_753),
.B(n_749),
.C(n_737),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_755),
.A2(n_718),
.B1(n_658),
.B2(n_724),
.Y(n_759)
);

AOI211x1_ASAP7_75t_SL g760 ( 
.A1(n_758),
.A2(n_754),
.B(n_757),
.C(n_720),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_759),
.B(n_741),
.Y(n_761)
);

AOI211xp5_ASAP7_75t_L g762 ( 
.A1(n_758),
.A2(n_526),
.B(n_677),
.C(n_672),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_761),
.B(n_740),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_760),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

OA22x2_ASAP7_75t_L g766 ( 
.A1(n_761),
.A2(n_657),
.B1(n_729),
.B2(n_731),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_761),
.Y(n_767)
);

NOR2x1_ASAP7_75t_L g768 ( 
.A(n_761),
.B(n_621),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_767),
.B(n_640),
.Y(n_769)
);

NAND4xp75_ASAP7_75t_L g770 ( 
.A(n_764),
.B(n_657),
.C(n_552),
.D(n_713),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_765),
.A2(n_677),
.B(n_720),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_768),
.Y(n_772)
);

NOR3x1_ASAP7_75t_L g773 ( 
.A(n_766),
.B(n_727),
.C(n_690),
.Y(n_773)
);

AOI221xp5_ASAP7_75t_L g774 ( 
.A1(n_763),
.A2(n_690),
.B1(n_703),
.B2(n_687),
.C(n_711),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_768),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_772),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_775),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_770),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_769),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_771),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_774),
.A2(n_674),
.B(n_640),
.C(n_682),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_773),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_776),
.Y(n_783)
);

XOR2xp5_ASAP7_75t_L g784 ( 
.A(n_779),
.B(n_632),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_777),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_778),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_780),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_782),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_781),
.Y(n_789)
);

OAI22xp33_ASAP7_75t_L g790 ( 
.A1(n_782),
.A2(n_621),
.B1(n_674),
.B2(n_624),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_778),
.A2(n_621),
.B1(n_682),
.B2(n_589),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_783),
.B(n_589),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_786),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_785),
.B(n_715),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_787),
.A2(n_788),
.B1(n_789),
.B2(n_790),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_784),
.A2(n_596),
.B1(n_593),
.B2(n_687),
.Y(n_796)
);

OAI31xp33_ASAP7_75t_L g797 ( 
.A1(n_791),
.A2(n_580),
.A3(n_567),
.B(n_643),
.Y(n_797)
);

AO22x2_ASAP7_75t_L g798 ( 
.A1(n_787),
.A2(n_596),
.B1(n_593),
.B2(n_588),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_786),
.B(n_683),
.Y(n_799)
);

OAI31xp33_ASAP7_75t_L g800 ( 
.A1(n_787),
.A2(n_580),
.A3(n_643),
.B(n_680),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_793),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_792),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_798),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_799),
.Y(n_804)
);

OAI22x1_ASAP7_75t_L g805 ( 
.A1(n_796),
.A2(n_588),
.B1(n_606),
.B2(n_671),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_801),
.A2(n_795),
.B1(n_794),
.B2(n_798),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_804),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_806),
.B(n_803),
.C(n_802),
.Y(n_808)
);

AOI222xp33_ASAP7_75t_L g809 ( 
.A1(n_808),
.A2(n_807),
.B1(n_805),
.B2(n_797),
.C1(n_800),
.C2(n_535),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_809),
.B(n_683),
.Y(n_810)
);

OAI211xp5_ASAP7_75t_L g811 ( 
.A1(n_810),
.A2(n_535),
.B(n_544),
.C(n_671),
.Y(n_811)
);


endmodule