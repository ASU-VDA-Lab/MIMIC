module fake_jpeg_17891_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_1),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_20),
.Y(n_25)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_4),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_12),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_27),
.B(n_31),
.Y(n_34)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_6),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.C(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_36),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);


endmodule