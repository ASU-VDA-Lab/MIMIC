module fake_jpeg_6138_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_19),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_19),
.B1(n_30),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_49),
.A2(n_53),
.B1(n_82),
.B2(n_4),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_76),
.B1(n_84),
.B2(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_62),
.Y(n_114)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_65),
.A2(n_78),
.B1(n_9),
.B2(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_69),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_39),
.A2(n_18),
.B1(n_16),
.B2(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_2),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_14),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_79),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_111),
.B1(n_87),
.B2(n_70),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_55),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_82),
.B1(n_53),
.B2(n_50),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_9),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_115),
.B(n_120),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_117),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_92),
.B1(n_93),
.B2(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_54),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_52),
.B1(n_56),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_129),
.B1(n_134),
.B2(n_140),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_61),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_62),
.B(n_74),
.C(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_135),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_56),
.B1(n_52),
.B2(n_71),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_81),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_103),
.B(n_11),
.C(n_13),
.D(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_85),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_81),
.B1(n_77),
.B2(n_51),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_85),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_87),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_99),
.Y(n_163)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_97),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_88),
.Y(n_154)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_117),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_103),
.A3(n_104),
.B1(n_95),
.B2(n_102),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_152),
.B1(n_163),
.B2(n_154),
.C(n_164),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_92),
.B(n_11),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_134),
.B(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_128),
.B1(n_124),
.B2(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_100),
.B1(n_99),
.B2(n_13),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_134),
.B(n_133),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_142),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_119),
.B1(n_134),
.B2(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_181),
.B(n_152),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_180),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_123),
.B(n_142),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_139),
.B(n_129),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_122),
.C(n_137),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_176),
.C(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_11),
.C(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_173),
.C(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_165),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_143),
.B1(n_145),
.B2(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_189),
.B(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_157),
.C(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_176),
.C(n_182),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_196),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_182),
.C(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_194),
.C(n_195),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_196),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_209),
.Y(n_212)
);


endmodule